module fake_netlist_5_1556_n_5157 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_5157);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_5157;

wire n_924;
wire n_977;
wire n_2253;
wire n_2756;
wire n_2417;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_2091;
wire n_1517;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_882;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_4255;
wire n_1796;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_2100;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_1385;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_870;
wire n_1711;
wire n_1891;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_1194;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_4391;
wire n_949;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1994;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_757;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_4918;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_978;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_4294;
wire n_1732;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_962;
wire n_723;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_974;
wire n_727;
wire n_4967;
wire n_957;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_815;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_4452;
wire n_4348;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_885;
wire n_5063;
wire n_2125;
wire n_3771;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_802;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_3178;
wire n_873;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_972;
wire n_3040;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_943;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_789;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_1109;
wire n_2605;
wire n_1310;
wire n_4747;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_4538;
wire n_766;
wire n_1117;
wire n_2754;
wire n_1742;
wire n_2489;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_3691;
wire n_3628;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_886;
wire n_1221;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_2476;
wire n_704;
wire n_4399;
wire n_2781;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_816;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1012;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_781;
wire n_3521;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_1018;
wire n_2247;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_5088;
wire n_2302;
wire n_951;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_902;
wire n_4991;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_3060;
wire n_4276;
wire n_3013;
wire n_1984;
wire n_2408;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_1097;
wire n_1036;
wire n_798;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_3985;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_858;
wire n_2985;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_892;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_4353;
wire n_2042;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_822;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_705;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_906;
wire n_919;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_1132;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_2878;
wire n_874;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_921;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_967;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_2637;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_984;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_1176;
wire n_1149;
wire n_1020;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_849;
wire n_1786;
wire n_4997;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_969;
wire n_1401;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_1702;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_2649;
wire n_1187;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_1174;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_1059;
wire n_1133;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_985;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3973;
wire n_3670;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_1178;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_1625;
wire n_2130;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1238;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_2260;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_3289;
wire n_1973;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_1087;
wire n_3472;
wire n_2874;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_844;
wire n_3497;
wire n_1601;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2505;
wire n_2427;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_1130;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_4881;
wire n_5089;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_4636;
wire n_4584;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_927;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_915;
wire n_864;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_947;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_1230;
wire n_4144;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_4483;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_955;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_897;
wire n_1428;
wire n_1216;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_1248;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_857;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_2808;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_914;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_946;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_1090;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_1639;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_1017;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_743;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_765;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3927;
wire n_3698;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_4891;
wire n_1023;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_1060;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_4608;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_1504;
wire n_3956;
wire n_3572;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_842;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_894;
wire n_3253;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_830;
wire n_3085;
wire n_1655;
wire n_749;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_1653;
wire n_1506;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_2608;
wire n_2657;
wire n_770;
wire n_2852;
wire n_2392;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_4679;
wire n_4115;
wire n_726;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1777;
wire n_1335;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_707;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_895;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_732;
wire n_4743;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_916;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_823;
wire n_725;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_719;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_1063;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_3852;
wire n_812;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_905;
wire n_5077;
wire n_782;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_4723;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_787;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_1028;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_3512;
wire n_4939;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_720;
wire n_2500;
wire n_1918;
wire n_863;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_2004;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_4474;
wire n_1089;
wire n_1004;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_1528;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_1545;
wire n_2374;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_1799;
wire n_2396;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_4197;
wire n_4829;
wire n_976;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_4944;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_1547;
wire n_777;
wire n_1755;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_923;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_1202;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_1072;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_706;
wire n_746;
wire n_784;
wire n_3978;
wire n_4809;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_913;
wire n_3833;
wire n_865;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_3471;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_724;
wire n_2084;
wire n_1781;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5108;
wire n_4692;
wire n_959;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_750;
wire n_742;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_5054;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_1209;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_4541;
wire n_3824;
wire n_3388;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_764;
wire n_1424;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_1432;
wire n_3875;
wire n_4003;
wire n_2402;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3382;
wire n_3574;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_896;
wire n_3316;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_4682;
wire n_3708;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_1188;
wire n_3957;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_1110;
wire n_3123;
wire n_5056;
wire n_1088;
wire n_3393;
wire n_866;
wire n_4887;
wire n_4617;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_1375;
wire n_3727;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_4987;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_899;
wire n_2722;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_710;
wire n_3090;
wire n_1168;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_791;
wire n_1533;
wire n_5036;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_3757;
wire n_3381;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_1170;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_825;
wire n_2819;
wire n_737;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_792;
wire n_3140;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_1225;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_3302;
wire n_1223;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_1086;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_852;
wire n_4602;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1975;
wire n_1321;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_2135;
wire n_3493;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_1076;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_730;
wire n_795;
wire n_4345;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_712;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_2839;
wire n_1588;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

INVx1_ASAP7_75t_L g703 ( 
.A(n_244),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_680),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_578),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_590),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_199),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_131),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_518),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_600),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_279),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_173),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_632),
.Y(n_713)
);

CKINVDCx16_ASAP7_75t_R g714 ( 
.A(n_696),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_217),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_478),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_144),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_247),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_363),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_658),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_585),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_233),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_507),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_582),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_300),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_695),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_653),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_372),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_207),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_240),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_601),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_691),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_113),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_248),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_654),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_3),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_369),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_559),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_489),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_397),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_277),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_165),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_343),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_8),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_414),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_120),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_598),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_383),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_193),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_419),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_323),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_129),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_57),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_40),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_400),
.Y(n_755)
);

BUFx2_ASAP7_75t_SL g756 ( 
.A(n_153),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_113),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_539),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_93),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_86),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_416),
.Y(n_761)
);

CKINVDCx14_ASAP7_75t_R g762 ( 
.A(n_264),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_642),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_120),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_654),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_451),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_285),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_68),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_506),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_373),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_343),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_572),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_110),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_685),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_334),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_433),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_328),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_453),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_687),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_468),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_657),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_10),
.Y(n_783)
);

BUFx10_ASAP7_75t_L g784 ( 
.A(n_667),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_660),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_580),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_699),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_146),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_137),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_481),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_594),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_550),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_566),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_311),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_402),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_183),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_674),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_259),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_98),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_134),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_229),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_257),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_346),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_527),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_168),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_633),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_319),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_525),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_203),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_317),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_650),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_361),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_664),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_544),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_135),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_463),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_73),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_491),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_532),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_374),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_552),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_386),
.Y(n_822)
);

BUFx10_ASAP7_75t_L g823 ( 
.A(n_570),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_563),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_65),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_12),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_326),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_338),
.Y(n_828)
);

BUFx10_ASAP7_75t_L g829 ( 
.A(n_240),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_496),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_436),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_177),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_642),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_262),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_309),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_275),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_595),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_59),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_515),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_214),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_42),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_439),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_386),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_179),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_658),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_662),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_437),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_641),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_357),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_663),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_569),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_651),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_648),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_9),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_182),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_149),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_473),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_68),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_652),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_57),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_347),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_490),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_530),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_246),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_126),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_233),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_362),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_539),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_634),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_656),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_318),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_514),
.Y(n_872)
);

BUFx8_ASAP7_75t_SL g873 ( 
.A(n_69),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_264),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_481),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_290),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_519),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_443),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_477),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_498),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_45),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_460),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_302),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_582),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_4),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_333),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_374),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_627),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_148),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_202),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_202),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_419),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_583),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_502),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_541),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_359),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_631),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_597),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_625),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_101),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_18),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_442),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_691),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_411),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_536),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_524),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_332),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_211),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_254),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_488),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_84),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_640),
.Y(n_912)
);

BUFx5_ASAP7_75t_L g913 ( 
.A(n_5),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_1),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_242),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_585),
.Y(n_916)
);

CKINVDCx14_ASAP7_75t_R g917 ( 
.A(n_661),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_663),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_548),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_268),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_307),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_108),
.Y(n_922)
);

BUFx8_ASAP7_75t_SL g923 ( 
.A(n_455),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_617),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_572),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_166),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_340),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_415),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_697),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_617),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_524),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_175),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_476),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_99),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_73),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_655),
.Y(n_936)
);

CKINVDCx16_ASAP7_75t_R g937 ( 
.A(n_509),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_609),
.Y(n_938)
);

BUFx10_ASAP7_75t_L g939 ( 
.A(n_571),
.Y(n_939)
);

INVxp33_ASAP7_75t_L g940 ( 
.A(n_491),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_579),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_659),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_335),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_85),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_430),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_674),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_589),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_413),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_186),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_220),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_409),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_681),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_440),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_621),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_625),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_80),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_218),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_597),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_643),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_359),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_402),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_592),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_117),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_4),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_559),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_60),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_82),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_485),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_241),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_309),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_127),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_519),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_131),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_229),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_278),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_280),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_358),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_440),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_377),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_373),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_64),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_344),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_141),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_666),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_311),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_665),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_257),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_363),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_564),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_37),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_689),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_185),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_339),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_69),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_615),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_353),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_574),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_599),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_549),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_99),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_379),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_700),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_101),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_210),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_205),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_589),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_635),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_444),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_484),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_586),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_669),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_648),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_608),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_659),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_253),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_667),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_356),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_504),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_449),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_547),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_7),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_245),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_603),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_457),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_310),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_668),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_261),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_88),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_317),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_414),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_600),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_449),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_16),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_666),
.Y(n_1034)
);

BUFx2_ASAP7_75t_SL g1035 ( 
.A(n_673),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_672),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_573),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_81),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_913),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_913),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_741),
.Y(n_1041)
);

BUFx8_ASAP7_75t_SL g1042 ( 
.A(n_914),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_873),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_913),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_923),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_913),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_913),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_913),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_913),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_899),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_899),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_899),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_740),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_751),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_762),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_736),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_730),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_917),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_714),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_730),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_734),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_761),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_739),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_734),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_941),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_941),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_955),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_740),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_740),
.Y(n_1069)
);

INVx4_ASAP7_75t_R g1070 ( 
.A(n_709),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_769),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_740),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_740),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_914),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_757),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_916),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_758),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_757),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_758),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_758),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_961),
.Y(n_1081)
);

INVxp33_ASAP7_75t_SL g1082 ( 
.A(n_770),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_981),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_758),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_937),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_758),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_781),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_781),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_847),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_744),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_949),
.Y(n_1091)
);

INVxp33_ASAP7_75t_SL g1092 ( 
.A(n_744),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1001),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_710),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_781),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_781),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_781),
.Y(n_1097)
);

BUFx5_ASAP7_75t_L g1098 ( 
.A(n_703),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_822),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_822),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_885),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_822),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_822),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_822),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_855),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_855),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_855),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_783),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_855),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_855),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_940),
.B(n_0),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_936),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_826),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1037),
.B(n_0),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_936),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_854),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_964),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_713),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_885),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_767),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_936),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_936),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_936),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_715),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_705),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_708),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_717),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_711),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_763),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_712),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_720),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_784),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_764),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_721),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_727),
.Y(n_1135)
);

INVxp33_ASAP7_75t_SL g1136 ( 
.A(n_1021),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_728),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_784),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_732),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_784),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_1021),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_765),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_766),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_743),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_767),
.Y(n_1145)
);

CKINVDCx16_ASAP7_75t_R g1146 ( 
.A(n_793),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_793),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_745),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_746),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_747),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_748),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_768),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_750),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_793),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_753),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_773),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_774),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_796),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_823),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_817),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_754),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_778),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_779),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_980),
.B(n_0),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_823),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_759),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_782),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_760),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_785),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_771),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_823),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_775),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_786),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_788),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_772),
.Y(n_1175)
);

INVxp33_ASAP7_75t_SL g1176 ( 
.A(n_704),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_792),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_776),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_777),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_716),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_780),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_798),
.Y(n_1182)
);

CKINVDCx14_ASAP7_75t_R g1183 ( 
.A(n_829),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_799),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_800),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_716),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_704),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_787),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_795),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_829),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_997),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_706),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_797),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_718),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_801),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_802),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_804),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_803),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_808),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_810),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_812),
.Y(n_1201)
);

CKINVDCx14_ASAP7_75t_R g1202 ( 
.A(n_829),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_818),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_772),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_718),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_825),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_791),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_827),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_805),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_833),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_837),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_806),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_789),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_807),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_809),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_811),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_839),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_789),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_843),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_814),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_849),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_819),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_853),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_848),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_857),
.Y(n_1225)
);

BUFx5_ASAP7_75t_L g1226 ( 
.A(n_858),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_848),
.Y(n_1227)
);

INVxp33_ASAP7_75t_SL g1228 ( 
.A(n_706),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_848),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_859),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_886),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_862),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_865),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_820),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_790),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_866),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_790),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_868),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_870),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_821),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_877),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_824),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_878),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1024),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_879),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_895),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_886),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_900),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_907),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_723),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_830),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_908),
.Y(n_1252)
);

BUFx2_ASAP7_75t_SL g1253 ( 
.A(n_886),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_831),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_888),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_911),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_912),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_794),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_927),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_928),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_794),
.Y(n_1261)
);

INVxp33_ASAP7_75t_L g1262 ( 
.A(n_816),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_888),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_931),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_935),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_834),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_938),
.Y(n_1267)
);

CKINVDCx14_ASAP7_75t_R g1268 ( 
.A(n_888),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_835),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_709),
.B(n_2),
.Y(n_1270)
);

XNOR2xp5_ASAP7_75t_SL g1271 ( 
.A(n_723),
.B(n_724),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_942),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_944),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_719),
.B(n_1),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_947),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_898),
.Y(n_1276)
);

NOR2xp67_ASAP7_75t_L g1277 ( 
.A(n_719),
.B(n_1),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_898),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_950),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_957),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_898),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_836),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_958),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_959),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_963),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_791),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_971),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_840),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_979),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_815),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_841),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_985),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_986),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_987),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_988),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_989),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_993),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_934),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_844),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_996),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_845),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_816),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_998),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_755),
.B(n_2),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_724),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1005),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_846),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1011),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1012),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1020),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1023),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_842),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1025),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_934),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1026),
.Y(n_1315)
);

INVxp33_ASAP7_75t_L g1316 ( 
.A(n_842),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1027),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_934),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1028),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_755),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1030),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1032),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_863),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_881),
.B(n_707),
.Y(n_1324)
);

BUFx2_ASAP7_75t_SL g1325 ( 
.A(n_939),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_881),
.B(n_2),
.Y(n_1326)
);

BUFx8_ASAP7_75t_SL g1327 ( 
.A(n_815),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_828),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_828),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_850),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_863),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_920),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_920),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_965),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_965),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1007),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1007),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1029),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1029),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_939),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_851),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_852),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_939),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_756),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1035),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_856),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_860),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_722),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_861),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_864),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_867),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_869),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_874),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_875),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_876),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_882),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_891),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_892),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_893),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_894),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_832),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_896),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_897),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_901),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_832),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_903),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_904),
.Y(n_1367)
);

CKINVDCx16_ASAP7_75t_R g1368 ( 
.A(n_838),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_905),
.Y(n_1369)
);

CKINVDCx16_ASAP7_75t_R g1370 ( 
.A(n_838),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_906),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_909),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_910),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_880),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_915),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_918),
.Y(n_1376)
);

BUFx5_ASAP7_75t_L g1377 ( 
.A(n_919),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_921),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_922),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_924),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_752),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_926),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_929),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_930),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_932),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_933),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_943),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_880),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_945),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_L g1390 ( 
.A(n_946),
.B(n_3),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_951),
.B(n_3),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_952),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_953),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_954),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_962),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_966),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_967),
.Y(n_1397)
);

INVxp33_ASAP7_75t_L g1398 ( 
.A(n_925),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_968),
.Y(n_1399)
);

CKINVDCx16_ASAP7_75t_R g1400 ( 
.A(n_925),
.Y(n_1400)
);

BUFx2_ASAP7_75t_SL g1401 ( 
.A(n_956),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_956),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1069),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1118),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1053),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1123),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1077),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1059),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1079),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1084),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1124),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1127),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1086),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1087),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1129),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1133),
.B(n_969),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1075),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1169),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_1173),
.B(n_4),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1174),
.B(n_5),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1053),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1177),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1182),
.B(n_970),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1088),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1184),
.B(n_972),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1059),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1095),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1071),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1185),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1096),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1253),
.Y(n_1431)
);

INVxp33_ASAP7_75t_L g1432 ( 
.A(n_1090),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1048),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1075),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1195),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1078),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1196),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1078),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1097),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1120),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1099),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1197),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1100),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1209),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1212),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1048),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1214),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1348),
.B(n_973),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1068),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1123),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1103),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1215),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1216),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1104),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1071),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1220),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_L g1457 ( 
.A(n_1222),
.B(n_1362),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1105),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1325),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1076),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1106),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1107),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1367),
.B(n_974),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1369),
.B(n_975),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1109),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1375),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1110),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1382),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1381),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1076),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1112),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1392),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1120),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1121),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1122),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1072),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1396),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1072),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1399),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1045),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1108),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1068),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1039),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1113),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1187),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1044),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1145),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1046),
.Y(n_1488)
);

INVxp33_ASAP7_75t_L g1489 ( 
.A(n_1101),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1145),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1047),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1377),
.B(n_976),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1116),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1052),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1117),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1327),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1052),
.Y(n_1497)
);

CKINVDCx16_ASAP7_75t_R g1498 ( 
.A(n_1183),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1261),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1327),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1085),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1094),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1323),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1175),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1094),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1050),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1175),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1051),
.Y(n_1508)
);

CKINVDCx14_ASAP7_75t_R g1509 ( 
.A(n_1183),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1073),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1073),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1204),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1080),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1055),
.B(n_977),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1142),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1080),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1204),
.Y(n_1517)
);

XNOR2xp5_ASAP7_75t_L g1518 ( 
.A(n_1398),
.B(n_1019),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1102),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1102),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1115),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1115),
.Y(n_1522)
);

CKINVDCx16_ASAP7_75t_R g1523 ( 
.A(n_1202),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1123),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1142),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1125),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1143),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1377),
.B(n_978),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1258),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1126),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1377),
.B(n_982),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1143),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1207),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1128),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1152),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1130),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1207),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1131),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1134),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1135),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1085),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1137),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1139),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1360),
.Y(n_1545)
);

CKINVDCx16_ASAP7_75t_R g1546 ( 
.A(n_1202),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1058),
.B(n_983),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1040),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1144),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_SL g1550 ( 
.A(n_1141),
.Y(n_1550)
);

CKINVDCx16_ASAP7_75t_R g1551 ( 
.A(n_1268),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1152),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1286),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1156),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1286),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_SL g1556 ( 
.A(n_1141),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1290),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1148),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1156),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_SL g1560 ( 
.A(n_1141),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1057),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1157),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1149),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1290),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1150),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1151),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1258),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1328),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1328),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1329),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1153),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1157),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1155),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1161),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1162),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1162),
.B(n_984),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1163),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1166),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1163),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1168),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1329),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1167),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1361),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1377),
.B(n_1346),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1167),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1234),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1234),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1170),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_R g1589 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1172),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1250),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1178),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1361),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1365),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_R g1595 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1251),
.Y(n_1596)
);

BUFx10_ASAP7_75t_L g1597 ( 
.A(n_1091),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1040),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1179),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1251),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1181),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1254),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1254),
.B(n_991),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1266),
.B(n_992),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1365),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1374),
.Y(n_1606)
);

NOR2xp67_ASAP7_75t_L g1607 ( 
.A(n_1266),
.B(n_5),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1374),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1188),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1305),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1360),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1189),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1402),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1402),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1193),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1119),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1198),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1269),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1368),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1199),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1269),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1200),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1282),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1201),
.Y(n_1624)
);

CKINVDCx20_ASAP7_75t_R g1625 ( 
.A(n_1042),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1378),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1042),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1378),
.B(n_994),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1203),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1377),
.B(n_1350),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1282),
.Y(n_1631)
);

CKINVDCx16_ASAP7_75t_R g1632 ( 
.A(n_1268),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1206),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1192),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1370),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1388),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1208),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1210),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_R g1639 ( 
.A(n_1288),
.B(n_725),
.Y(n_1639)
);

CKINVDCx16_ASAP7_75t_R g1640 ( 
.A(n_1400),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1288),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1211),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1091),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1049),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1217),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1291),
.B(n_995),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1291),
.B(n_6),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1299),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1074),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1258),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1219),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1299),
.Y(n_1652)
);

NOR2xp67_ASAP7_75t_L g1653 ( 
.A(n_1301),
.B(n_6),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1221),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_1132),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1074),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1223),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1301),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1307),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1225),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1230),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1307),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1043),
.Y(n_1663)
);

INVxp33_ASAP7_75t_SL g1664 ( 
.A(n_1093),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1330),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1049),
.Y(n_1666)
);

INVxp33_ASAP7_75t_L g1667 ( 
.A(n_1324),
.Y(n_1667)
);

INVxp33_ASAP7_75t_SL g1668 ( 
.A(n_1093),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1330),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1389),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1159),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1171),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1232),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1341),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1341),
.B(n_1342),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1233),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1342),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1401),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_1043),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1236),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_1138),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1347),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1238),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1239),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1241),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1243),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1146),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1245),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1258),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1347),
.B(n_999),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1246),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1248),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1249),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1255),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1252),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1256),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1355),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1257),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1355),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1389),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1259),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1349),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1061),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1263),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1190),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1260),
.Y(n_1706)
);

INVxp67_ASAP7_75t_SL g1707 ( 
.A(n_1394),
.Y(n_1707)
);

CKINVDCx16_ASAP7_75t_R g1708 ( 
.A(n_1140),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1483),
.B(n_1486),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1492),
.B(n_1377),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1650),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1526),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1530),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1619),
.A2(n_1009),
.B1(n_1019),
.B2(n_990),
.Y(n_1714)
);

AND2x6_ASAP7_75t_L g1715 ( 
.A(n_1584),
.B(n_1394),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1650),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1529),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1671),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1529),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1469),
.B(n_1092),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1529),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1650),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1667),
.A2(n_1316),
.B1(n_1262),
.B2(n_1270),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1535),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1537),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1488),
.B(n_1377),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1639),
.A2(n_1082),
.B1(n_1136),
.B2(n_1092),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1539),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1667),
.A2(n_1114),
.B1(n_1082),
.B2(n_1009),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1672),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1649),
.Y(n_1731)
);

INVx5_ASAP7_75t_L g1732 ( 
.A(n_1529),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1540),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1567),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1576),
.A2(n_1136),
.B1(n_1228),
.B2(n_1176),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1476),
.B(n_1060),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1603),
.A2(n_1176),
.B1(n_1228),
.B2(n_1063),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1567),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1567),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1541),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1543),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1544),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1491),
.B(n_1098),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1567),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1478),
.B(n_1060),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1448),
.B(n_1062),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1549),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1558),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1689),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1563),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1565),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1566),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1571),
.Y(n_1754)
);

OA21x2_ASAP7_75t_L g1755 ( 
.A1(n_1630),
.A2(n_1397),
.B(n_1352),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1604),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1573),
.Y(n_1757)
);

AOI22x1_ASAP7_75t_SL g1758 ( 
.A1(n_1625),
.A2(n_1031),
.B1(n_1033),
.B2(n_990),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1689),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1548),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1574),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1578),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1548),
.B(n_1098),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1406),
.B(n_1450),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1509),
.B(n_1054),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1509),
.B(n_1397),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1646),
.A2(n_1351),
.B1(n_1354),
.B2(n_1353),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1580),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1406),
.B(n_1064),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1588),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1450),
.Y(n_1771)
);

CKINVDCx11_ASAP7_75t_R g1772 ( 
.A(n_1625),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1524),
.B(n_1065),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1607),
.A2(n_1033),
.B1(n_1031),
.B2(n_1041),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1561),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1590),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1690),
.A2(n_1675),
.B1(n_1423),
.B2(n_1425),
.Y(n_1777)
);

AND2x6_ASAP7_75t_L g1778 ( 
.A(n_1628),
.B(n_1356),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1561),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1703),
.B(n_1066),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1528),
.B(n_1098),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1598),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_SL g1783 ( 
.A(n_1647),
.B(n_813),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1703),
.Y(n_1784)
);

OA21x2_ASAP7_75t_L g1785 ( 
.A1(n_1531),
.A2(n_1358),
.B(n_1357),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1592),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1498),
.B(n_1229),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1598),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1599),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1644),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1601),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1635),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1644),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1523),
.B(n_1318),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1609),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1666),
.B(n_1433),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1612),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1499),
.B(n_1359),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1615),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1482),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1404),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1514),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1482),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1666),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1482),
.Y(n_1805)
);

BUFx8_ASAP7_75t_L g1806 ( 
.A(n_1550),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1403),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1411),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1407),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1409),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1410),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_L g1812 ( 
.A(n_1503),
.B(n_1098),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1546),
.B(n_1551),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_SL g1814 ( 
.A(n_1653),
.B(n_872),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1413),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1617),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1414),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1632),
.B(n_1363),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1424),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1616),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1427),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1547),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1432),
.B(n_1364),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1430),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1432),
.B(n_1489),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1620),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1439),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1441),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1443),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1416),
.B(n_1387),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1419),
.B(n_902),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1451),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1622),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1454),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1420),
.B(n_1098),
.Y(n_1835)
);

INVx5_ASAP7_75t_L g1836 ( 
.A(n_1405),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1458),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1412),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1461),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1545),
.B(n_1366),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1489),
.B(n_1431),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1624),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1611),
.B(n_1626),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1462),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1459),
.B(n_1371),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1629),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1670),
.B(n_1372),
.Y(n_1847)
);

INVx3_ASAP7_75t_L g1848 ( 
.A(n_1405),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1465),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1633),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1700),
.B(n_1707),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1421),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1637),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1467),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1446),
.B(n_1098),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1471),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1474),
.Y(n_1857)
);

BUFx8_ASAP7_75t_L g1858 ( 
.A(n_1550),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1463),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1475),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1421),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1449),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1636),
.A2(n_1518),
.B1(n_1398),
.B2(n_1640),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1681),
.A2(n_726),
.B1(n_729),
.B2(n_725),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1449),
.Y(n_1865)
);

NAND2xp33_ASAP7_75t_SL g1866 ( 
.A(n_1550),
.B(n_726),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1638),
.Y(n_1867)
);

AND2x6_ASAP7_75t_L g1868 ( 
.A(n_1464),
.B(n_1373),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1510),
.B(n_1098),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1485),
.B(n_1376),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1642),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1591),
.A2(n_1081),
.B1(n_1083),
.B2(n_1067),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1610),
.A2(n_1634),
.B1(n_1457),
.B2(n_1534),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1645),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1506),
.Y(n_1875)
);

INVx6_ASAP7_75t_L g1876 ( 
.A(n_1708),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1511),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1508),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1651),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1654),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1657),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1589),
.B(n_1595),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1513),
.B(n_1226),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1415),
.B(n_1226),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1660),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1516),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_L g1887 ( 
.A(n_1661),
.B(n_1380),
.C(n_1379),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1673),
.B(n_1383),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1519),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1676),
.B(n_1384),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1680),
.B(n_1385),
.Y(n_1891)
);

INVx4_ASAP7_75t_L g1892 ( 
.A(n_1418),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1683),
.B(n_1393),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1684),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1520),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1685),
.B(n_1395),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1686),
.B(n_1344),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1688),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1678),
.B(n_1262),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1691),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1692),
.B(n_1345),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1521),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1693),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1695),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1696),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1522),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1494),
.B(n_1226),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1698),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1497),
.B(n_1226),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1701),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1556),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1706),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1408),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1597),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1422),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1597),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1426),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1597),
.Y(n_1918)
);

BUFx8_ASAP7_75t_L g1919 ( 
.A(n_1556),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1429),
.B(n_1226),
.Y(n_1920)
);

OA21x2_ASAP7_75t_L g1921 ( 
.A1(n_1435),
.A2(n_1186),
.B(n_1180),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1437),
.B(n_1226),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1442),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1444),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1445),
.B(n_1226),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1447),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1452),
.B(n_1312),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1428),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1455),
.B(n_1056),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1453),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1460),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1502),
.A2(n_1111),
.B1(n_1160),
.B2(n_1158),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1505),
.A2(n_1244),
.B1(n_1191),
.B2(n_1274),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1456),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1470),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1466),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_SL g1937 ( 
.A1(n_1681),
.A2(n_731),
.B1(n_733),
.B2(n_729),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1468),
.B(n_1312),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1472),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1477),
.Y(n_1940)
);

INVx5_ASAP7_75t_L g1941 ( 
.A(n_1655),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1501),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1542),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1479),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1481),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1687),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1484),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1493),
.B(n_1312),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1643),
.Y(n_1949)
);

BUFx8_ASAP7_75t_L g1950 ( 
.A(n_1556),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1515),
.A2(n_1304),
.B1(n_1326),
.B2(n_1277),
.Y(n_1951)
);

OAI22x1_ASAP7_75t_SL g1952 ( 
.A1(n_1649),
.A2(n_733),
.B1(n_735),
.B2(n_731),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1495),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1525),
.B(n_1312),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1527),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1532),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1536),
.B(n_1331),
.Y(n_1957)
);

OAI21x1_ASAP7_75t_L g1958 ( 
.A1(n_1560),
.A2(n_1186),
.B(n_1180),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1552),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1554),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1559),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1704),
.B(n_1140),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1702),
.B(n_1349),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1562),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1572),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1575),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1577),
.B(n_1316),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1579),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1687),
.A2(n_737),
.B1(n_738),
.B2(n_735),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1582),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1664),
.A2(n_1668),
.B1(n_1586),
.B2(n_1587),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1585),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1596),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1600),
.Y(n_1974)
);

CKINVDCx11_ASAP7_75t_R g1975 ( 
.A(n_1627),
.Y(n_1975)
);

INVx5_ASAP7_75t_L g1976 ( 
.A(n_1560),
.Y(n_1976)
);

BUFx8_ASAP7_75t_L g1977 ( 
.A(n_1560),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1602),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1618),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1621),
.B(n_1154),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1623),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1631),
.B(n_1331),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1641),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1648),
.B(n_1331),
.Y(n_1984)
);

NOR2x1_ASAP7_75t_L g1985 ( 
.A(n_1694),
.B(n_1154),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1652),
.B(n_1227),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1658),
.B(n_1264),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1659),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1662),
.B(n_1227),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1665),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1669),
.A2(n_1340),
.B1(n_1165),
.B2(n_1224),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1674),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1677),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1682),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1697),
.B(n_1231),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1699),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1480),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1923),
.Y(n_1998)
);

NAND2xp33_ASAP7_75t_R g1999 ( 
.A(n_1718),
.B(n_1496),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1712),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1930),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1731),
.Y(n_2002)
);

BUFx3_ASAP7_75t_L g2003 ( 
.A(n_1775),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1930),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1713),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1731),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1930),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1775),
.Y(n_2008)
);

CKINVDCx20_ASAP7_75t_R g2009 ( 
.A(n_1863),
.Y(n_2009)
);

CKINVDCx20_ASAP7_75t_R g2010 ( 
.A(n_1714),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1946),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1930),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1760),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1934),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1724),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1934),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1934),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1730),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1782),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1934),
.Y(n_2020)
);

BUFx2_ASAP7_75t_L g2021 ( 
.A(n_1730),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1944),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1944),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1944),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_R g2025 ( 
.A(n_1911),
.B(n_1500),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1944),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1772),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_R g2028 ( 
.A(n_1911),
.B(n_1627),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1772),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_R g2030 ( 
.A(n_1866),
.B(n_1608),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1975),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1975),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1725),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1801),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1801),
.Y(n_2035)
);

CKINVDCx16_ASAP7_75t_R g2036 ( 
.A(n_1813),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1792),
.Y(n_2037)
);

AOI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1835),
.A2(n_1164),
.B(n_1390),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1728),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1808),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1808),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1733),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1775),
.Y(n_2043)
);

CKINVDCx16_ASAP7_75t_R g2044 ( 
.A(n_1765),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1838),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1756),
.B(n_1349),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1838),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_1743),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_R g2049 ( 
.A(n_1866),
.B(n_1613),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1756),
.B(n_1386),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1788),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1892),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1790),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1775),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1892),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1793),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1865),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1924),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1848),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_R g2060 ( 
.A(n_1997),
.B(n_1614),
.Y(n_2060)
);

NOR2xp67_ASAP7_75t_L g2061 ( 
.A(n_1976),
.B(n_1147),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1740),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1924),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1947),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1848),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1779),
.Y(n_2066)
);

NOR2xp67_ASAP7_75t_L g2067 ( 
.A(n_1976),
.B(n_1298),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1947),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1955),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1955),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1955),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1955),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1741),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1966),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_R g2075 ( 
.A(n_1997),
.B(n_1663),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1966),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1742),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_1966),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1966),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1899),
.B(n_1340),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1748),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1749),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1973),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1879),
.B(n_1265),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1973),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_1743),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1825),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1973),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1747),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1751),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1843),
.A2(n_1694),
.B1(n_1704),
.B2(n_1391),
.Y(n_2091)
);

CKINVDCx20_ASAP7_75t_R g2092 ( 
.A(n_1968),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1752),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1973),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1753),
.Y(n_2095)
);

INVxp33_ASAP7_75t_L g2096 ( 
.A(n_1967),
.Y(n_2096)
);

CKINVDCx20_ASAP7_75t_R g2097 ( 
.A(n_1968),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_R g2098 ( 
.A(n_1956),
.B(n_1663),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1994),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_1784),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1852),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1843),
.A2(n_1272),
.B1(n_1273),
.B2(n_1267),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1754),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1994),
.Y(n_2104)
);

HB1xp67_ASAP7_75t_L g2105 ( 
.A(n_1784),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1757),
.Y(n_2106)
);

BUFx4f_ASAP7_75t_L g2107 ( 
.A(n_1914),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1994),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1994),
.Y(n_2109)
);

CKINVDCx20_ASAP7_75t_R g2110 ( 
.A(n_1876),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_1996),
.Y(n_2111)
);

BUFx10_ASAP7_75t_L g2112 ( 
.A(n_1967),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_1996),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1761),
.Y(n_2114)
);

NOR2xp67_ASAP7_75t_L g2115 ( 
.A(n_1976),
.B(n_1314),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1762),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1768),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1996),
.Y(n_2118)
);

AO21x2_ASAP7_75t_L g2119 ( 
.A1(n_1710),
.A2(n_1333),
.B(n_1332),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1830),
.A2(n_1279),
.B1(n_1280),
.B2(n_1275),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1996),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1770),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1852),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1806),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1806),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1776),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_R g2127 ( 
.A(n_1956),
.B(n_1679),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_R g2128 ( 
.A(n_1974),
.B(n_1679),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_1858),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1858),
.Y(n_2130)
);

CKINVDCx20_ASAP7_75t_R g2131 ( 
.A(n_1876),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1786),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_1919),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1919),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_1841),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1950),
.Y(n_2136)
);

INVx8_ASAP7_75t_L g2137 ( 
.A(n_1778),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1789),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1791),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1861),
.Y(n_2140)
);

HB1xp67_ASAP7_75t_L g2141 ( 
.A(n_1954),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1954),
.Y(n_2142)
);

CKINVDCx20_ASAP7_75t_R g2143 ( 
.A(n_1876),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1950),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1977),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1977),
.Y(n_2146)
);

BUFx10_ASAP7_75t_L g2147 ( 
.A(n_1989),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1941),
.Y(n_2148)
);

CKINVDCx20_ASAP7_75t_R g2149 ( 
.A(n_1971),
.Y(n_2149)
);

OA21x2_ASAP7_75t_L g2150 ( 
.A1(n_1744),
.A2(n_1855),
.B(n_1726),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_1779),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1941),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1941),
.Y(n_2153)
);

BUFx3_ASAP7_75t_L g2154 ( 
.A(n_1779),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1941),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1914),
.Y(n_2156)
);

BUFx2_ASAP7_75t_L g2157 ( 
.A(n_1820),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1795),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_1859),
.B(n_1386),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1914),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1914),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1916),
.Y(n_2162)
);

AND2x6_ASAP7_75t_L g2163 ( 
.A(n_1920),
.B(n_1343),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1916),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1797),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1799),
.Y(n_2166)
);

NAND2xp33_ASAP7_75t_R g2167 ( 
.A(n_1787),
.B(n_737),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1916),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1916),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1816),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1861),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1759),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_R g2173 ( 
.A(n_1974),
.B(n_1553),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1750),
.Y(n_2174)
);

CKINVDCx6p67_ASAP7_75t_R g2175 ( 
.A(n_1976),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_1957),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_1918),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_1720),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1918),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1826),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1833),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1918),
.Y(n_2182)
);

CKINVDCx20_ASAP7_75t_R g2183 ( 
.A(n_1727),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1918),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1915),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1842),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1750),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1926),
.Y(n_2188)
);

CKINVDCx20_ASAP7_75t_R g2189 ( 
.A(n_1794),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1846),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1936),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1939),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1940),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1945),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1953),
.Y(n_2195)
);

INVx5_ASAP7_75t_L g2196 ( 
.A(n_1804),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1983),
.Y(n_2197)
);

NOR2xp67_ASAP7_75t_L g2198 ( 
.A(n_1993),
.B(n_1231),
.Y(n_2198)
);

BUFx2_ASAP7_75t_L g2199 ( 
.A(n_1820),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_1983),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1800),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1850),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1777),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_1804),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_1767),
.B(n_1002),
.C(n_1000),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1859),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1800),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1882),
.Y(n_2208)
);

CKINVDCx20_ASAP7_75t_R g2209 ( 
.A(n_1864),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1882),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1823),
.B(n_1247),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1853),
.Y(n_2212)
);

INVxp67_ASAP7_75t_SL g2213 ( 
.A(n_1804),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1867),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1957),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1960),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_1970),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_R g2218 ( 
.A(n_1959),
.B(n_1564),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1972),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1979),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1990),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1989),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1995),
.Y(n_2223)
);

CKINVDCx20_ASAP7_75t_R g2224 ( 
.A(n_1937),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_R g2225 ( 
.A(n_1961),
.B(n_1564),
.Y(n_2225)
);

BUFx3_ASAP7_75t_L g2226 ( 
.A(n_1779),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1871),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1995),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1720),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1874),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1880),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1881),
.Y(n_2232)
);

INVx3_ASAP7_75t_L g2233 ( 
.A(n_1804),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_1802),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_1894),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1885),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1803),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1802),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1822),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1803),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1898),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1870),
.B(n_1247),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1851),
.B(n_1920),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1900),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1805),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1822),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_1982),
.B(n_1386),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1805),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1905),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1908),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_1982),
.B(n_1089),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_R g2252 ( 
.A(n_1964),
.B(n_1570),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1965),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1978),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1912),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_1981),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1894),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1912),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1886),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1988),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1886),
.Y(n_2261)
);

CKINVDCx20_ASAP7_75t_R g2262 ( 
.A(n_1969),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1902),
.Y(n_2263)
);

CKINVDCx20_ASAP7_75t_R g2264 ( 
.A(n_1758),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1992),
.Y(n_2265)
);

CKINVDCx20_ASAP7_75t_R g2266 ( 
.A(n_1873),
.Y(n_2266)
);

INVx8_ASAP7_75t_L g2267 ( 
.A(n_1778),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1796),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1796),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_R g2270 ( 
.A(n_1913),
.B(n_1570),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_1927),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1780),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1927),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_1938),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1780),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1938),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1879),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_1948),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1875),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1948),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_1735),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_1980),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1986),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1984),
.Y(n_2284)
);

CKINVDCx20_ASAP7_75t_R g2285 ( 
.A(n_1737),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_1984),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_1830),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1902),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_1830),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1830),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_R g2291 ( 
.A(n_1917),
.B(n_1581),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1830),
.Y(n_2292)
);

BUFx2_ASAP7_75t_L g2293 ( 
.A(n_1987),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_1868),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1875),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1868),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1878),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1868),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_1987),
.B(n_1276),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_1862),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1878),
.Y(n_2301)
);

CKINVDCx20_ASAP7_75t_R g2302 ( 
.A(n_1963),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1862),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_1888),
.B(n_1283),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1868),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_1868),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_1932),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1862),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1932),
.Y(n_2309)
);

CKINVDCx20_ASAP7_75t_R g2310 ( 
.A(n_1729),
.Y(n_2310)
);

NOR2xp67_ASAP7_75t_L g2311 ( 
.A(n_1771),
.B(n_1276),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_R g2312 ( 
.A(n_1928),
.B(n_1593),
.Y(n_2312)
);

CKINVDCx20_ASAP7_75t_R g2313 ( 
.A(n_1729),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_R g2314 ( 
.A(n_1931),
.B(n_1593),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_R g2315 ( 
.A(n_1935),
.B(n_1594),
.Y(n_2315)
);

CKINVDCx20_ASAP7_75t_R g2316 ( 
.A(n_1774),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_1933),
.Y(n_2317)
);

NOR2xp67_ASAP7_75t_L g2318 ( 
.A(n_1771),
.B(n_1278),
.Y(n_2318)
);

INVx4_ASAP7_75t_SL g2319 ( 
.A(n_2163),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2268),
.B(n_1922),
.Y(n_2320)
);

INVx4_ASAP7_75t_L g2321 ( 
.A(n_2156),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2269),
.B(n_1922),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_2054),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2243),
.A2(n_1884),
.B(n_1925),
.Y(n_2324)
);

INVx4_ASAP7_75t_L g2325 ( 
.A(n_2160),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2141),
.B(n_1925),
.Y(n_2326)
);

INVx2_ASAP7_75t_SL g2327 ( 
.A(n_2018),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2013),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2203),
.A2(n_1723),
.B1(n_1847),
.B2(n_1840),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2013),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2019),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_SL g2332 ( 
.A(n_2107),
.B(n_1783),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2110),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2142),
.B(n_1715),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2019),
.Y(n_2335)
);

INVx4_ASAP7_75t_L g2336 ( 
.A(n_2161),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2176),
.B(n_1715),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_SL g2338 ( 
.A(n_2271),
.B(n_1840),
.Y(n_2338)
);

INVx1_ASAP7_75t_SL g2339 ( 
.A(n_2021),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_2178),
.B(n_1783),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2051),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2215),
.B(n_1715),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2089),
.B(n_1942),
.Y(n_2343)
);

AOI22xp33_ASAP7_75t_L g2344 ( 
.A1(n_2163),
.A2(n_1785),
.B1(n_1715),
.B2(n_1778),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2277),
.B(n_1764),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1998),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2273),
.B(n_1715),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2274),
.B(n_1778),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2051),
.Y(n_2349)
);

CKINVDCx6p67_ASAP7_75t_R g2350 ( 
.A(n_2002),
.Y(n_2350)
);

INVx4_ASAP7_75t_SL g2351 ( 
.A(n_2163),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2053),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2272),
.B(n_2275),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2053),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2056),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2110),
.Y(n_2356)
);

NAND2xp33_ASAP7_75t_L g2357 ( 
.A(n_2287),
.B(n_1778),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2276),
.B(n_1855),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2056),
.Y(n_2359)
);

INVx2_ASAP7_75t_SL g2360 ( 
.A(n_2157),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_SL g2361 ( 
.A(n_2112),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2278),
.B(n_1847),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2084),
.B(n_1764),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2057),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2131),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2131),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2057),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2259),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2001),
.Y(n_2369)
);

OR2x6_ASAP7_75t_L g2370 ( 
.A(n_2293),
.B(n_1962),
.Y(n_2370)
);

BUFx3_ASAP7_75t_L g2371 ( 
.A(n_2143),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2280),
.B(n_2229),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2259),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2163),
.B(n_1785),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2284),
.B(n_1831),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2172),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2087),
.B(n_1943),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2172),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2004),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2163),
.B(n_1755),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_SL g2381 ( 
.A(n_2107),
.B(n_1814),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2163),
.B(n_1755),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2199),
.B(n_1949),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2080),
.B(n_1929),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2286),
.B(n_1831),
.Y(n_2385)
);

AOI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_2289),
.A2(n_1884),
.B1(n_1812),
.B2(n_1798),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_2211),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2162),
.B(n_1814),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2164),
.B(n_1894),
.Y(n_2389)
);

OR2x6_ASAP7_75t_L g2390 ( 
.A(n_2086),
.B(n_1985),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2261),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2150),
.B(n_1921),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2096),
.B(n_2206),
.Y(n_2393)
);

AND2x6_ASAP7_75t_L g2394 ( 
.A(n_2120),
.B(n_2299),
.Y(n_2394)
);

OAI22xp33_ASAP7_75t_L g2395 ( 
.A1(n_2307),
.A2(n_2309),
.B1(n_2313),
.B2(n_2310),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2150),
.B(n_1921),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2168),
.B(n_1894),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2261),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2048),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2169),
.B(n_1903),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2048),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2177),
.B(n_1903),
.Y(n_2402)
);

INVx3_ASAP7_75t_L g2403 ( 
.A(n_2054),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2201),
.Y(n_2404)
);

INVx5_ASAP7_75t_L g2405 ( 
.A(n_2137),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2179),
.B(n_1903),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2084),
.B(n_1888),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2135),
.B(n_1933),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_2007),
.Y(n_2409)
);

BUFx10_ASAP7_75t_L g2410 ( 
.A(n_2046),
.Y(n_2410)
);

XNOR2xp5_ASAP7_75t_L g2411 ( 
.A(n_2037),
.B(n_1473),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2242),
.B(n_1929),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2150),
.B(n_1726),
.Y(n_2413)
);

AOI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_2310),
.A2(n_1798),
.B1(n_1812),
.B2(n_1891),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2096),
.B(n_1766),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2201),
.Y(n_2416)
);

INVx4_ASAP7_75t_L g2417 ( 
.A(n_2182),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2234),
.B(n_1963),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_2313),
.A2(n_1891),
.B1(n_1893),
.B2(n_1901),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2263),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2054),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2238),
.B(n_1723),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2263),
.Y(n_2423)
);

INVx4_ASAP7_75t_SL g2424 ( 
.A(n_2235),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_SL g2425 ( 
.A(n_2184),
.B(n_1903),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2288),
.B(n_2255),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2288),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2207),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2054),
.Y(n_2429)
);

INVx5_ASAP7_75t_L g2430 ( 
.A(n_2137),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_SL g2431 ( 
.A(n_2012),
.B(n_1904),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_2066),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2258),
.B(n_1709),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_2014),
.B(n_1904),
.Y(n_2434)
);

AND3x2_ASAP7_75t_L g2435 ( 
.A(n_2159),
.B(n_1818),
.C(n_1845),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2207),
.Y(n_2436)
);

AOI22xp33_ASAP7_75t_L g2437 ( 
.A1(n_2000),
.A2(n_1893),
.B1(n_1901),
.B2(n_1709),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2237),
.Y(n_2438)
);

AND2x6_ASAP7_75t_L g2439 ( 
.A(n_2279),
.B(n_1773),
.Y(n_2439)
);

INVx4_ASAP7_75t_L g2440 ( 
.A(n_2066),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_2066),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2005),
.A2(n_1910),
.B1(n_1904),
.B2(n_1896),
.Y(n_2442)
);

INVx4_ASAP7_75t_SL g2443 ( 
.A(n_2235),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2237),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2240),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_2066),
.Y(n_2446)
);

NAND2xp33_ASAP7_75t_L g2447 ( 
.A(n_2290),
.B(n_1904),
.Y(n_2447)
);

OAI22xp33_ASAP7_75t_SL g2448 ( 
.A1(n_2208),
.A2(n_1774),
.B1(n_1951),
.B2(n_1991),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2295),
.B(n_1896),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2297),
.B(n_2301),
.Y(n_2450)
);

AOI22xp33_ASAP7_75t_L g2451 ( 
.A1(n_2015),
.A2(n_1910),
.B1(n_1890),
.B2(n_1835),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2240),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2016),
.B(n_1910),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2044),
.B(n_1872),
.Y(n_2454)
);

INVx2_ASAP7_75t_SL g2455 ( 
.A(n_2304),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2239),
.B(n_1951),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2247),
.B(n_1890),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2245),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2245),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2248),
.Y(n_2460)
);

INVx1_ASAP7_75t_SL g2461 ( 
.A(n_2069),
.Y(n_2461)
);

AND2x6_ASAP7_75t_L g2462 ( 
.A(n_2248),
.B(n_1773),
.Y(n_2462)
);

OR2x2_ASAP7_75t_SL g2463 ( 
.A(n_2036),
.B(n_1656),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2059),
.Y(n_2464)
);

INVx3_ASAP7_75t_L g2465 ( 
.A(n_2235),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2246),
.B(n_1656),
.Y(n_2466)
);

OR2x2_ASAP7_75t_L g2467 ( 
.A(n_2100),
.B(n_1872),
.Y(n_2467)
);

INVx3_ASAP7_75t_L g2468 ( 
.A(n_2235),
.Y(n_2468)
);

OR2x6_ASAP7_75t_L g2469 ( 
.A(n_2137),
.B(n_2267),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2033),
.Y(n_2470)
);

AOI22xp33_ASAP7_75t_L g2471 ( 
.A1(n_2039),
.A2(n_2042),
.B1(n_2073),
.B2(n_2062),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2077),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2081),
.Y(n_2473)
);

NAND2xp33_ASAP7_75t_L g2474 ( 
.A(n_2292),
.B(n_1910),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2059),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2294),
.B(n_2296),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2065),
.Y(n_2477)
);

BUFx6f_ASAP7_75t_L g2478 ( 
.A(n_2003),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2003),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_2143),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2082),
.Y(n_2481)
);

AOI22xp33_ASAP7_75t_L g2482 ( 
.A1(n_2316),
.A2(n_948),
.B1(n_960),
.B2(n_1897),
.Y(n_2482)
);

OR2x6_ASAP7_75t_L g2483 ( 
.A(n_2137),
.B(n_1769),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2017),
.B(n_1769),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2298),
.B(n_1744),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2008),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2065),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2090),
.A2(n_1821),
.B1(n_1834),
.B2(n_1810),
.Y(n_2488)
);

CKINVDCx20_ASAP7_75t_R g2489 ( 
.A(n_2002),
.Y(n_2489)
);

OAI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2317),
.A2(n_1887),
.B1(n_1897),
.B2(n_742),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2084),
.B(n_2304),
.Y(n_2491)
);

BUFx3_ASAP7_75t_L g2492 ( 
.A(n_2037),
.Y(n_2492)
);

AND2x6_ASAP7_75t_L g2493 ( 
.A(n_2093),
.B(n_1736),
.Y(n_2493)
);

INVxp67_ASAP7_75t_SL g2494 ( 
.A(n_2257),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2305),
.B(n_1781),
.Y(n_2495)
);

OAI22xp33_ASAP7_75t_SL g2496 ( 
.A1(n_2210),
.A2(n_742),
.B1(n_749),
.B2(n_738),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2306),
.B(n_1781),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2008),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2095),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2103),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2106),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2105),
.B(n_1736),
.Y(n_2502)
);

OR2x6_ASAP7_75t_L g2503 ( 
.A(n_2267),
.B(n_1746),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2257),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2070),
.Y(n_2505)
);

BUFx2_ASAP7_75t_L g2506 ( 
.A(n_2011),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2114),
.Y(n_2507)
);

BUFx3_ASAP7_75t_L g2508 ( 
.A(n_2020),
.Y(n_2508)
);

BUFx4f_ASAP7_75t_L g2509 ( 
.A(n_2175),
.Y(n_2509)
);

INVx5_ASAP7_75t_L g2510 ( 
.A(n_2267),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2101),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2116),
.Y(n_2512)
);

INVx6_ASAP7_75t_L g2513 ( 
.A(n_2043),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2304),
.B(n_1746),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2257),
.Y(n_2515)
);

INVx6_ASAP7_75t_L g2516 ( 
.A(n_2043),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2117),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_L g2518 ( 
.A(n_2267),
.B(n_2257),
.Y(n_2518)
);

BUFx3_ASAP7_75t_L g2519 ( 
.A(n_2022),
.Y(n_2519)
);

INVx4_ASAP7_75t_SL g2520 ( 
.A(n_2151),
.Y(n_2520)
);

AND2x6_ASAP7_75t_L g2521 ( 
.A(n_2122),
.B(n_2126),
.Y(n_2521)
);

INVx4_ASAP7_75t_L g2522 ( 
.A(n_2023),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2251),
.B(n_1089),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2132),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2024),
.B(n_1857),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2138),
.B(n_1907),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2071),
.Y(n_2527)
);

NAND2xp33_ASAP7_75t_R g2528 ( 
.A(n_2270),
.B(n_2291),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_2151),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2101),
.Y(n_2530)
);

BUFx8_ASAP7_75t_SL g2531 ( 
.A(n_2006),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_L g2532 ( 
.A1(n_2139),
.A2(n_1821),
.B1(n_1834),
.B2(n_1810),
.Y(n_2532)
);

NAND3xp33_ASAP7_75t_L g2533 ( 
.A(n_2050),
.B(n_1809),
.C(n_1807),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2072),
.Y(n_2534)
);

BUFx6f_ASAP7_75t_L g2535 ( 
.A(n_2154),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2123),
.Y(n_2536)
);

AND3x1_ASAP7_75t_L g2537 ( 
.A(n_2091),
.B(n_1952),
.C(n_1271),
.Y(n_2537)
);

OAI22xp33_ASAP7_75t_SL g2538 ( 
.A1(n_2222),
.A2(n_871),
.B1(n_883),
.B2(n_749),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2026),
.B(n_2185),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2074),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2223),
.B(n_1417),
.Y(n_2541)
);

AND2x2_ASAP7_75t_SL g2542 ( 
.A(n_2010),
.B(n_1417),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2188),
.B(n_2191),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2076),
.B(n_1089),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2192),
.B(n_1810),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2158),
.Y(n_2546)
);

INVx4_ASAP7_75t_SL g2547 ( 
.A(n_2154),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2165),
.B(n_1907),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2166),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2170),
.B(n_1909),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2180),
.A2(n_1710),
.B1(n_1821),
.B2(n_1810),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2193),
.B(n_1821),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2181),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2226),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2228),
.B(n_1278),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2194),
.B(n_1834),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2186),
.B(n_1909),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_2078),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2190),
.Y(n_2559)
);

INVx2_ASAP7_75t_SL g2560 ( 
.A(n_2079),
.Y(n_2560)
);

BUFx3_ASAP7_75t_L g2561 ( 
.A(n_2083),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2226),
.Y(n_2562)
);

AND3x2_ASAP7_75t_L g2563 ( 
.A(n_2202),
.B(n_1285),
.C(n_1284),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2195),
.B(n_1839),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2123),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2085),
.B(n_1281),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2212),
.B(n_1763),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2214),
.B(n_1763),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2227),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2140),
.Y(n_2570)
);

AO22x2_ASAP7_75t_L g2571 ( 
.A1(n_2316),
.A2(n_1281),
.B1(n_1289),
.B2(n_1287),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2230),
.Y(n_2572)
);

INVx2_ASAP7_75t_SL g2573 ( 
.A(n_2088),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2231),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2232),
.B(n_1811),
.Y(n_2575)
);

INVx4_ASAP7_75t_L g2576 ( 
.A(n_2094),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2099),
.B(n_1320),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2236),
.B(n_2241),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2244),
.B(n_2249),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2104),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2112),
.B(n_1434),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2011),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2250),
.B(n_1877),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2140),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2171),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2108),
.B(n_2109),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2111),
.B(n_1320),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2171),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2119),
.A2(n_1839),
.B1(n_1849),
.B2(n_1834),
.Y(n_2589)
);

AOI22xp33_ASAP7_75t_L g2590 ( 
.A1(n_2119),
.A2(n_883),
.B1(n_884),
.B2(n_871),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2300),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2300),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2174),
.Y(n_2593)
);

BUFx6f_ASAP7_75t_L g2594 ( 
.A(n_2113),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2303),
.B(n_1889),
.Y(n_2595)
);

BUFx4f_ASAP7_75t_L g2596 ( 
.A(n_2303),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2311),
.B(n_1815),
.Y(n_2597)
);

INVx6_ASAP7_75t_L g2598 ( 
.A(n_2112),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2216),
.A2(n_1849),
.B1(n_1857),
.B2(n_1839),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2118),
.B(n_1320),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2308),
.B(n_1895),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2205),
.A2(n_1849),
.B1(n_1857),
.B2(n_1839),
.Y(n_2602)
);

INVxp33_ASAP7_75t_L g2603 ( 
.A(n_2312),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2121),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2282),
.B(n_1434),
.Y(n_2605)
);

INVx3_ASAP7_75t_L g2606 ( 
.A(n_2308),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2283),
.B(n_1817),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2174),
.Y(n_2608)
);

INVx4_ASAP7_75t_SL g2609 ( 
.A(n_2148),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2187),
.A2(n_1857),
.B1(n_1849),
.B2(n_1824),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_2281),
.B(n_1819),
.Y(n_2611)
);

AND2x6_ASAP7_75t_L g2612 ( 
.A(n_2204),
.B(n_1734),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2187),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2204),
.B(n_1906),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2217),
.B(n_1827),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2102),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2147),
.B(n_2219),
.Y(n_2617)
);

OAI22xp33_ASAP7_75t_L g2618 ( 
.A1(n_2285),
.A2(n_2265),
.B1(n_2254),
.B2(n_2256),
.Y(n_2618)
);

INVxp67_ASAP7_75t_L g2619 ( 
.A(n_2167),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2204),
.Y(n_2620)
);

NAND2xp33_ASAP7_75t_L g2621 ( 
.A(n_2034),
.B(n_1738),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2233),
.Y(n_2622)
);

INVxp67_ASAP7_75t_SL g2623 ( 
.A(n_2233),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_SL g2624 ( 
.A(n_2035),
.B(n_884),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2233),
.Y(n_2625)
);

INVx4_ASAP7_75t_L g2626 ( 
.A(n_2058),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2038),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2196),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2220),
.B(n_1828),
.Y(n_2629)
);

NOR2xp33_ASAP7_75t_SL g2630 ( 
.A(n_2040),
.B(n_887),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2183),
.A2(n_1832),
.B1(n_1837),
.B2(n_1829),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2213),
.Y(n_2632)
);

NAND2xp33_ASAP7_75t_SL g2633 ( 
.A(n_2041),
.B(n_1436),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_2147),
.B(n_1436),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2221),
.A2(n_1854),
.B1(n_1856),
.B2(n_1844),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_L g2636 ( 
.A(n_2147),
.B(n_2253),
.Y(n_2636)
);

INVx4_ASAP7_75t_L g2637 ( 
.A(n_2063),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2196),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2045),
.B(n_1860),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2260),
.B(n_1958),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2197),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2318),
.B(n_1869),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_2047),
.B(n_1717),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2196),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2052),
.B(n_2055),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2006),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2196),
.Y(n_2647)
);

INVx4_ASAP7_75t_L g2648 ( 
.A(n_2064),
.Y(n_2648)
);

BUFx2_ASAP7_75t_L g2649 ( 
.A(n_2189),
.Y(n_2649)
);

OAI21xp33_ASAP7_75t_SL g2650 ( 
.A1(n_2198),
.A2(n_1883),
.B(n_1869),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2196),
.B(n_1883),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2068),
.B(n_1862),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_L g2653 ( 
.A(n_2200),
.B(n_1438),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2061),
.B(n_1438),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2152),
.Y(n_2655)
);

INVx4_ASAP7_75t_SL g2656 ( 
.A(n_2153),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2155),
.Y(n_2657)
);

OR2x2_ASAP7_75t_L g2658 ( 
.A(n_2067),
.B(n_1292),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2115),
.B(n_1711),
.Y(n_2659)
);

BUFx10_ASAP7_75t_L g2660 ( 
.A(n_2027),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2189),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2266),
.B(n_1716),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2092),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2183),
.A2(n_1722),
.B1(n_1745),
.B2(n_1739),
.Y(n_2664)
);

INVxp67_ASAP7_75t_SL g2665 ( 
.A(n_2092),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2097),
.Y(n_2666)
);

HB1xp67_ASAP7_75t_L g2667 ( 
.A(n_2314),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2097),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2302),
.Y(n_2669)
);

INVx4_ASAP7_75t_L g2670 ( 
.A(n_2124),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2060),
.B(n_1739),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2315),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2149),
.Y(n_2673)
);

INVx4_ASAP7_75t_L g2674 ( 
.A(n_2125),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2218),
.B(n_1717),
.Y(n_2675)
);

INVx5_ASAP7_75t_L g2676 ( 
.A(n_1999),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2457),
.B(n_2173),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2457),
.B(n_2075),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2328),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2384),
.B(n_2098),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2676),
.B(n_2127),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2358),
.B(n_2326),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2358),
.B(n_2128),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2676),
.B(n_2225),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2326),
.B(n_2252),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2354),
.Y(n_2686)
);

OR2x2_ASAP7_75t_L g2687 ( 
.A(n_2661),
.B(n_2372),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2320),
.B(n_2149),
.Y(n_2688)
);

INVx3_ASAP7_75t_L g2689 ( 
.A(n_2620),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_L g2690 ( 
.A(n_2372),
.B(n_2340),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_SL g2691 ( 
.A(n_2346),
.B(n_2029),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2415),
.B(n_2030),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2320),
.B(n_1717),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2322),
.B(n_1717),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2676),
.B(n_2049),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2322),
.B(n_1719),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2470),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2433),
.B(n_1719),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2355),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2376),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2676),
.B(n_2009),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2472),
.Y(n_2702)
);

NOR2xp67_ASAP7_75t_L g2703 ( 
.A(n_2522),
.B(n_2129),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2393),
.B(n_2009),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2378),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2433),
.B(n_2449),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2332),
.B(n_2025),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2449),
.B(n_2526),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2526),
.B(n_1719),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2548),
.B(n_1719),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2548),
.B(n_1721),
.Y(n_2711)
);

INVx4_ASAP7_75t_L g2712 ( 
.A(n_2594),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_2332),
.B(n_2028),
.Y(n_2713)
);

INVxp67_ASAP7_75t_L g2714 ( 
.A(n_2383),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_2412),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2381),
.B(n_1440),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2550),
.B(n_1721),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2381),
.B(n_2414),
.Y(n_2718)
);

AOI22xp5_ASAP7_75t_SL g2719 ( 
.A1(n_2418),
.A2(n_2010),
.B1(n_1473),
.B2(n_1487),
.Y(n_2719)
);

INVxp33_ASAP7_75t_L g2720 ( 
.A(n_2605),
.Y(n_2720)
);

NOR2x1p5_ASAP7_75t_L g2721 ( 
.A(n_2508),
.B(n_2031),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2329),
.B(n_1440),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2422),
.B(n_2209),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2464),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2475),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2473),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2550),
.B(n_1721),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2619),
.B(n_2395),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2432),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2481),
.Y(n_2730)
);

BUFx3_ASAP7_75t_L g2731 ( 
.A(n_2594),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2557),
.B(n_1721),
.Y(n_2732)
);

NAND2x1_ASAP7_75t_L g2733 ( 
.A(n_2469),
.B(n_1070),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2557),
.B(n_1331),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2567),
.B(n_1003),
.Y(n_2735)
);

NOR2x1p5_ASAP7_75t_L g2736 ( 
.A(n_2519),
.B(n_2032),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2586),
.B(n_1487),
.Y(n_2737)
);

NOR2x1p5_ASAP7_75t_L g2738 ( 
.A(n_2540),
.B(n_2130),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2477),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2567),
.B(n_2568),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2487),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2568),
.B(n_1004),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2578),
.B(n_2579),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2578),
.B(n_1006),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2511),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2579),
.B(n_1038),
.Y(n_2746)
);

OR2x2_ASAP7_75t_L g2747 ( 
.A(n_2339),
.B(n_1490),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2395),
.B(n_2619),
.Y(n_2748)
);

NAND2xp33_ASAP7_75t_L g2749 ( 
.A(n_2521),
.B(n_2133),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2329),
.B(n_2209),
.Y(n_2750)
);

NOR2xp67_ASAP7_75t_L g2751 ( 
.A(n_2522),
.B(n_2134),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2499),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2500),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2491),
.B(n_1594),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2523),
.B(n_1583),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2501),
.B(n_2507),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2512),
.B(n_887),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2530),
.Y(n_2758)
);

INVx2_ASAP7_75t_SL g2759 ( 
.A(n_2327),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2339),
.B(n_1490),
.Y(n_2760)
);

NOR3xp33_ASAP7_75t_L g2761 ( 
.A(n_2618),
.B(n_2144),
.C(n_2136),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_SL g2762 ( 
.A(n_2491),
.B(n_1504),
.Y(n_2762)
);

OAI221xp5_ASAP7_75t_L g2763 ( 
.A1(n_2482),
.A2(n_1008),
.B1(n_1010),
.B2(n_890),
.C(n_889),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_SL g2764 ( 
.A(n_2369),
.B(n_2379),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2517),
.B(n_889),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2524),
.B(n_890),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2461),
.B(n_1504),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2546),
.B(n_2549),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2338),
.A2(n_1512),
.B1(n_1517),
.B2(n_1507),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2536),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2565),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2570),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2553),
.B(n_1008),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_SL g2774 ( 
.A(n_2594),
.B(n_1507),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2584),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2588),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2608),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2613),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2559),
.Y(n_2779)
);

NAND3xp33_ASAP7_75t_L g2780 ( 
.A(n_2482),
.B(n_1517),
.C(n_1512),
.Y(n_2780)
);

INVxp67_ASAP7_75t_L g2781 ( 
.A(n_2343),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2569),
.B(n_2572),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2408),
.B(n_2224),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_2620),
.Y(n_2784)
);

NAND3xp33_ASAP7_75t_L g2785 ( 
.A(n_2466),
.B(n_1538),
.C(n_1533),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2574),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2467),
.B(n_2224),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2432),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2652),
.B(n_1010),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2618),
.B(n_1555),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2652),
.B(n_1013),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2407),
.B(n_1555),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2407),
.B(n_1557),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2616),
.B(n_1013),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2471),
.B(n_1014),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2387),
.B(n_1014),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2386),
.B(n_1015),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2485),
.B(n_1015),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_2461),
.B(n_1581),
.Y(n_2799)
);

NAND3xp33_ASAP7_75t_L g2800 ( 
.A(n_2541),
.B(n_1583),
.C(n_1569),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2419),
.B(n_2611),
.Y(n_2801)
);

NOR3xp33_ASAP7_75t_L g2802 ( 
.A(n_2456),
.B(n_2146),
.C(n_2145),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2485),
.B(n_1016),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2330),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_SL g2805 ( 
.A(n_2409),
.B(n_1605),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2331),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2335),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2341),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2362),
.A2(n_1538),
.B1(n_1553),
.B2(n_1533),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2375),
.B(n_2262),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2349),
.Y(n_2811)
);

BUFx5_ASAP7_75t_L g2812 ( 
.A(n_2521),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2385),
.B(n_2262),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2437),
.B(n_1016),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2442),
.B(n_1017),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2352),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2583),
.B(n_1017),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2583),
.B(n_1018),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_2558),
.B(n_1557),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2450),
.B(n_1018),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2450),
.B(n_1022),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2451),
.B(n_1022),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2359),
.Y(n_2823)
);

NOR3xp33_ASAP7_75t_L g2824 ( 
.A(n_2581),
.B(n_1294),
.C(n_1293),
.Y(n_2824)
);

NOR2xp67_ASAP7_75t_L g2825 ( 
.A(n_2576),
.B(n_1295),
.Y(n_2825)
);

OAI22xp33_ASAP7_75t_L g2826 ( 
.A1(n_2490),
.A2(n_1036),
.B1(n_1034),
.B2(n_1568),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2514),
.B(n_1568),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2413),
.B(n_1034),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2364),
.Y(n_2829)
);

INVxp67_ASAP7_75t_SL g2830 ( 
.A(n_2494),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_SL g2831 ( 
.A(n_2514),
.B(n_1569),
.Y(n_2831)
);

NAND2xp33_ASAP7_75t_L g2832 ( 
.A(n_2521),
.B(n_1036),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2413),
.B(n_1194),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_SL g2834 ( 
.A(n_2561),
.Y(n_2834)
);

INVx1_ASAP7_75t_SL g2835 ( 
.A(n_2360),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2607),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2454),
.B(n_1605),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2566),
.B(n_1606),
.Y(n_2838)
);

INVxp67_ASAP7_75t_L g2839 ( 
.A(n_2377),
.Y(n_2839)
);

NOR2xp67_ASAP7_75t_L g2840 ( 
.A(n_2576),
.B(n_1296),
.Y(n_2840)
);

BUFx5_ASAP7_75t_L g2841 ( 
.A(n_2521),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_L g2842 ( 
.A(n_2662),
.B(n_1606),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2577),
.B(n_1297),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2367),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2662),
.B(n_2264),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2347),
.B(n_1194),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2587),
.B(n_1300),
.Y(n_2847)
);

O2A1O1Ixp33_ASAP7_75t_L g2848 ( 
.A1(n_2347),
.A2(n_1306),
.B(n_1308),
.C(n_1303),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2448),
.B(n_2264),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2363),
.B(n_1309),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2600),
.B(n_1310),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2348),
.B(n_1205),
.Y(n_2852)
);

NOR2xp33_ASAP7_75t_L g2853 ( 
.A(n_2388),
.B(n_6),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2348),
.B(n_1205),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2426),
.B(n_1213),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2426),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2404),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2494),
.B(n_1213),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2416),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2575),
.B(n_1218),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2363),
.B(n_1311),
.Y(n_2861)
);

AOI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2394),
.A2(n_1315),
.B1(n_1317),
.B2(n_1313),
.Y(n_2862)
);

INVxp67_ASAP7_75t_SL g2863 ( 
.A(n_2432),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2575),
.B(n_1218),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2438),
.Y(n_2865)
);

HB1xp67_ASAP7_75t_L g2866 ( 
.A(n_2505),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2599),
.B(n_1235),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2617),
.B(n_1235),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2455),
.B(n_1319),
.Y(n_2869)
);

NAND2xp33_ASAP7_75t_L g2870 ( 
.A(n_2521),
.B(n_1732),
.Y(n_2870)
);

INVxp67_ASAP7_75t_L g2871 ( 
.A(n_2505),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2334),
.B(n_1237),
.Y(n_2872)
);

INVxp67_ASAP7_75t_L g2873 ( 
.A(n_2527),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2334),
.B(n_1237),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2337),
.B(n_2342),
.Y(n_2875)
);

INVxp67_ASAP7_75t_L g2876 ( 
.A(n_2527),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2444),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2368),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2373),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2636),
.B(n_7),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2458),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2459),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2337),
.B(n_1302),
.Y(n_2883)
);

OAI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2495),
.A2(n_1836),
.B1(n_1321),
.B2(n_1322),
.Y(n_2884)
);

NOR2xp67_ASAP7_75t_L g2885 ( 
.A(n_2604),
.B(n_1334),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2391),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2342),
.B(n_1302),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2632),
.B(n_1335),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2597),
.B(n_1336),
.Y(n_2889)
);

INVxp67_ASAP7_75t_L g2890 ( 
.A(n_2502),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2398),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2597),
.B(n_1337),
.Y(n_2892)
);

INVx2_ASAP7_75t_SL g2893 ( 
.A(n_2580),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2543),
.B(n_2669),
.Y(n_2894)
);

NOR2xp67_ASAP7_75t_L g2895 ( 
.A(n_2604),
.B(n_1338),
.Y(n_2895)
);

INVxp67_ASAP7_75t_SL g2896 ( 
.A(n_2623),
.Y(n_2896)
);

BUFx6f_ASAP7_75t_L g2897 ( 
.A(n_2478),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2420),
.Y(n_2898)
);

OAI22xp33_ASAP7_75t_L g2899 ( 
.A1(n_2490),
.A2(n_1339),
.B1(n_9),
.B2(n_7),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2423),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2603),
.B(n_8),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2590),
.B(n_1836),
.Y(n_2902)
);

INVxp67_ASAP7_75t_L g2903 ( 
.A(n_2649),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2427),
.Y(n_2904)
);

INVx5_ASAP7_75t_L g2905 ( 
.A(n_2469),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2585),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2590),
.B(n_1836),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2529),
.B(n_2554),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2529),
.B(n_1836),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2593),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2554),
.B(n_8),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2428),
.Y(n_2912)
);

NAND3xp33_ASAP7_75t_L g2913 ( 
.A(n_2631),
.B(n_1732),
.C(n_9),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_2673),
.B(n_16),
.Y(n_2914)
);

INVx8_ASAP7_75t_L g2915 ( 
.A(n_2483),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_SL g2916 ( 
.A(n_2534),
.B(n_1732),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2623),
.B(n_10),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2560),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2545),
.B(n_10),
.Y(n_2919)
);

INVxp67_ASAP7_75t_SL g2920 ( 
.A(n_2478),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2436),
.Y(n_2921)
);

BUFx3_ASAP7_75t_L g2922 ( 
.A(n_2333),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2445),
.Y(n_2923)
);

NAND2x1_ASAP7_75t_L g2924 ( 
.A(n_2469),
.B(n_1732),
.Y(n_2924)
);

INVx2_ASAP7_75t_SL g2925 ( 
.A(n_2573),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2452),
.Y(n_2926)
);

O2A1O1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_2324),
.A2(n_2495),
.B(n_2497),
.C(n_2374),
.Y(n_2927)
);

NOR2xp33_ASAP7_75t_L g2928 ( 
.A(n_2539),
.B(n_11),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2555),
.B(n_11),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2321),
.B(n_17),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2460),
.Y(n_2931)
);

NAND2xp33_ASAP7_75t_L g2932 ( 
.A(n_2493),
.B(n_2405),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2595),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2321),
.B(n_17),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2591),
.Y(n_2935)
);

INVx3_ASAP7_75t_L g2936 ( 
.A(n_2620),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2591),
.Y(n_2937)
);

NAND2xp33_ASAP7_75t_L g2938 ( 
.A(n_2493),
.B(n_2405),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2552),
.B(n_11),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2592),
.Y(n_2940)
);

NAND3xp33_ASAP7_75t_L g2941 ( 
.A(n_2624),
.B(n_12),
.C(n_13),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2556),
.B(n_12),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2564),
.B(n_13),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2592),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2595),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2642),
.B(n_13),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2642),
.B(n_14),
.Y(n_2947)
);

NAND2xp33_ASAP7_75t_L g2948 ( 
.A(n_2493),
.B(n_2405),
.Y(n_2948)
);

BUFx6f_ASAP7_75t_L g2949 ( 
.A(n_2478),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2497),
.B(n_2394),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2410),
.B(n_2624),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2394),
.B(n_14),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2325),
.B(n_18),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2394),
.B(n_14),
.Y(n_2954)
);

NOR2xp33_ASAP7_75t_L g2955 ( 
.A(n_2410),
.B(n_15),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2394),
.B(n_15),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2544),
.B(n_693),
.Y(n_2957)
);

NOR2xp67_ASAP7_75t_L g2958 ( 
.A(n_2325),
.B(n_15),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2431),
.B(n_2434),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2453),
.B(n_19),
.Y(n_2960)
);

NOR2x1p5_ASAP7_75t_L g2961 ( 
.A(n_2336),
.B(n_20),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2630),
.B(n_2634),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2525),
.B(n_19),
.Y(n_2963)
);

INVx3_ASAP7_75t_L g2964 ( 
.A(n_2440),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2606),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2601),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2353),
.B(n_20),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2630),
.B(n_696),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_SL g2969 ( 
.A(n_2336),
.B(n_21),
.Y(n_2969)
);

INVx4_ASAP7_75t_L g2970 ( 
.A(n_2479),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2731),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2682),
.B(n_2435),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2697),
.Y(n_2973)
);

INVxp67_ASAP7_75t_L g2974 ( 
.A(n_2866),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2702),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2726),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2730),
.Y(n_2977)
);

AO22x2_ASAP7_75t_L g2978 ( 
.A1(n_2718),
.A2(n_2665),
.B1(n_2666),
.B2(n_2663),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2752),
.Y(n_2979)
);

AO22x2_ASAP7_75t_L g2980 ( 
.A1(n_2780),
.A2(n_2665),
.B1(n_2668),
.B2(n_2351),
.Y(n_2980)
);

AO22x2_ASAP7_75t_L g2981 ( 
.A1(n_2722),
.A2(n_2351),
.B1(n_2319),
.B2(n_2374),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2753),
.Y(n_2982)
);

AO22x2_ASAP7_75t_L g2983 ( 
.A1(n_2952),
.A2(n_2351),
.B1(n_2319),
.B2(n_2571),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2779),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2786),
.Y(n_2985)
);

CKINVDCx5p33_ASAP7_75t_R g2986 ( 
.A(n_2834),
.Y(n_2986)
);

INVx2_ASAP7_75t_SL g2987 ( 
.A(n_2712),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2712),
.Y(n_2988)
);

AO22x2_ASAP7_75t_L g2989 ( 
.A1(n_2954),
.A2(n_2956),
.B1(n_2913),
.B2(n_2941),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2756),
.Y(n_2990)
);

NAND2x1p5_ASAP7_75t_L g2991 ( 
.A(n_2835),
.B(n_2417),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2768),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2782),
.Y(n_2993)
);

INVxp67_ASAP7_75t_L g2994 ( 
.A(n_2866),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2811),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2816),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2823),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2690),
.B(n_2435),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2844),
.Y(n_2999)
);

OAI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2740),
.A2(n_2476),
.B1(n_2532),
.B2(n_2488),
.Y(n_3000)
);

BUFx2_ASAP7_75t_L g3001 ( 
.A(n_2903),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2688),
.B(n_2542),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2878),
.Y(n_3003)
);

AO22x2_ASAP7_75t_L g3004 ( 
.A1(n_2801),
.A2(n_2319),
.B1(n_2571),
.B2(n_2640),
.Y(n_3004)
);

BUFx8_ASAP7_75t_L g3005 ( 
.A(n_2834),
.Y(n_3005)
);

INVxp67_ASAP7_75t_L g3006 ( 
.A(n_2687),
.Y(n_3006)
);

HB1xp67_ASAP7_75t_L g3007 ( 
.A(n_2836),
.Y(n_3007)
);

CKINVDCx16_ASAP7_75t_R g3008 ( 
.A(n_2764),
.Y(n_3008)
);

NOR2xp67_ASAP7_75t_L g3009 ( 
.A(n_2893),
.B(n_2626),
.Y(n_3009)
);

NAND2x1p5_ASAP7_75t_L g3010 ( 
.A(n_2970),
.B(n_2417),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2690),
.B(n_2641),
.Y(n_3011)
);

OAI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2743),
.A2(n_2476),
.B1(n_2596),
.B2(n_2551),
.Y(n_3012)
);

AO22x2_ASAP7_75t_L g3013 ( 
.A1(n_2950),
.A2(n_2790),
.B1(n_2800),
.B2(n_2785),
.Y(n_3013)
);

AO22x2_ASAP7_75t_L g3014 ( 
.A1(n_2716),
.A2(n_2571),
.B1(n_2382),
.B2(n_2380),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2879),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2804),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2886),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2891),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2898),
.Y(n_3019)
);

AND2x2_ASAP7_75t_SL g3020 ( 
.A(n_2750),
.B(n_2537),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2706),
.B(n_2353),
.Y(n_3021)
);

AO22x2_ASAP7_75t_L g3022 ( 
.A1(n_2701),
.A2(n_2382),
.B1(n_2380),
.B2(n_2533),
.Y(n_3022)
);

AOI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2842),
.A2(n_2653),
.B1(n_2633),
.B2(n_2528),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2904),
.Y(n_3024)
);

OA22x2_ASAP7_75t_L g3025 ( 
.A1(n_2769),
.A2(n_2411),
.B1(n_2390),
.B2(n_2401),
.Y(n_3025)
);

INVx2_ASAP7_75t_SL g3026 ( 
.A(n_2759),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2906),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2910),
.Y(n_3028)
);

BUFx8_ASAP7_75t_L g3029 ( 
.A(n_2767),
.Y(n_3029)
);

AND2x4_ASAP7_75t_L g3030 ( 
.A(n_2922),
.B(n_2918),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2806),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2912),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2708),
.B(n_2345),
.Y(n_3033)
);

AO22x2_ASAP7_75t_L g3034 ( 
.A1(n_2797),
.A2(n_2672),
.B1(n_2654),
.B2(n_2675),
.Y(n_3034)
);

OAI221xp5_ASAP7_75t_L g3035 ( 
.A1(n_2750),
.A2(n_2635),
.B1(n_2615),
.B2(n_2629),
.C(n_2667),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2807),
.Y(n_3036)
);

AO22x2_ASAP7_75t_L g3037 ( 
.A1(n_2677),
.A2(n_2675),
.B1(n_2627),
.B2(n_2397),
.Y(n_3037)
);

AO22x2_ASAP7_75t_L g3038 ( 
.A1(n_2678),
.A2(n_2400),
.B1(n_2402),
.B2(n_2389),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2808),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2923),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2926),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2842),
.A2(n_2645),
.B1(n_2667),
.B2(n_2484),
.Y(n_3042)
);

OAI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_2896),
.A2(n_2596),
.B1(n_2344),
.B2(n_2516),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2931),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2856),
.B(n_2345),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2829),
.Y(n_3046)
);

HB1xp67_ASAP7_75t_L g3047 ( 
.A(n_2871),
.Y(n_3047)
);

AO22x2_ASAP7_75t_L g3048 ( 
.A1(n_2685),
.A2(n_2425),
.B1(n_2406),
.B2(n_2626),
.Y(n_3048)
);

NAND2x1p5_ASAP7_75t_L g3049 ( 
.A(n_2970),
.B(n_2479),
.Y(n_3049)
);

AOI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_2837),
.A2(n_2370),
.B1(n_2390),
.B2(n_2637),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2860),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_2925),
.B(n_2356),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2864),
.Y(n_3053)
);

NAND2x1p5_ASAP7_75t_L g3054 ( 
.A(n_2905),
.B(n_2479),
.Y(n_3054)
);

OR2x2_ASAP7_75t_L g3055 ( 
.A(n_2747),
.B(n_2399),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2900),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2921),
.Y(n_3057)
);

AO22x2_ASAP7_75t_L g3058 ( 
.A1(n_2896),
.A2(n_2637),
.B1(n_2648),
.B2(n_2392),
.Y(n_3058)
);

BUFx8_ASAP7_75t_L g3059 ( 
.A(n_2737),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2683),
.B(n_2783),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2735),
.B(n_2658),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2679),
.Y(n_3062)
);

AO22x2_ASAP7_75t_L g3063 ( 
.A1(n_2830),
.A2(n_2648),
.B1(n_2392),
.B2(n_2396),
.Y(n_3063)
);

AO22x2_ASAP7_75t_L g3064 ( 
.A1(n_2830),
.A2(n_2396),
.B1(n_2671),
.B2(n_2656),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2686),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2699),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2700),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2705),
.Y(n_3068)
);

INVxp67_ASAP7_75t_L g3069 ( 
.A(n_2760),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2742),
.B(n_2671),
.Y(n_3070)
);

OR2x6_ASAP7_75t_L g3071 ( 
.A(n_2915),
.B(n_2506),
.Y(n_3071)
);

OR2x2_ASAP7_75t_SL g3072 ( 
.A(n_2914),
.B(n_2598),
.Y(n_3072)
);

AOI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_2837),
.A2(n_2370),
.B1(n_2390),
.B2(n_2639),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2783),
.B(n_2370),
.Y(n_3074)
);

NAND2x1p5_ASAP7_75t_L g3075 ( 
.A(n_2905),
.B(n_2486),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2787),
.B(n_2655),
.Y(n_3076)
);

INVx4_ASAP7_75t_L g3077 ( 
.A(n_2897),
.Y(n_3077)
);

AO22x2_ASAP7_75t_L g3078 ( 
.A1(n_2930),
.A2(n_2656),
.B1(n_2609),
.B2(n_2643),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2724),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2798),
.B(n_2664),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2725),
.Y(n_3081)
);

AO22x2_ASAP7_75t_L g3082 ( 
.A1(n_2934),
.A2(n_2656),
.B1(n_2609),
.B2(n_2646),
.Y(n_3082)
);

AND2x4_ASAP7_75t_L g3083 ( 
.A(n_2738),
.B(n_2365),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2739),
.Y(n_3084)
);

INVxp67_ASAP7_75t_L g3085 ( 
.A(n_2894),
.Y(n_3085)
);

AO22x2_ASAP7_75t_L g3086 ( 
.A1(n_2953),
.A2(n_2609),
.B1(n_2657),
.B2(n_2371),
.Y(n_3086)
);

BUFx4f_ASAP7_75t_L g3087 ( 
.A(n_2897),
.Y(n_3087)
);

CKINVDCx20_ASAP7_75t_R g3088 ( 
.A(n_2809),
.Y(n_3088)
);

AND2x4_ASAP7_75t_L g3089 ( 
.A(n_2715),
.B(n_2366),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2741),
.Y(n_3090)
);

AO22x2_ASAP7_75t_L g3091 ( 
.A1(n_2969),
.A2(n_2480),
.B1(n_2492),
.B2(n_2463),
.Y(n_3091)
);

NAND2x1p5_ASAP7_75t_L g3092 ( 
.A(n_2905),
.B(n_2486),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2723),
.B(n_2582),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2745),
.Y(n_3094)
);

NAND2x1p5_ASAP7_75t_L g3095 ( 
.A(n_2905),
.B(n_2486),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2758),
.Y(n_3096)
);

AO22x2_ASAP7_75t_L g3097 ( 
.A1(n_2713),
.A2(n_2622),
.B1(n_2625),
.B2(n_2496),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2723),
.B(n_2489),
.Y(n_3098)
);

AO22x2_ASAP7_75t_L g3099 ( 
.A1(n_2899),
.A2(n_2674),
.B1(n_2670),
.B2(n_2538),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2770),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2771),
.Y(n_3101)
);

AO22x2_ASAP7_75t_L g3102 ( 
.A1(n_2899),
.A2(n_2674),
.B1(n_2670),
.B2(n_2547),
.Y(n_3102)
);

AO22x2_ASAP7_75t_L g3103 ( 
.A1(n_2799),
.A2(n_2547),
.B1(n_2520),
.B2(n_2606),
.Y(n_3103)
);

BUFx8_ASAP7_75t_L g3104 ( 
.A(n_2838),
.Y(n_3104)
);

AND2x4_ASAP7_75t_L g3105 ( 
.A(n_2715),
.B(n_2483),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2890),
.B(n_2483),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2772),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2775),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2776),
.Y(n_3109)
);

NAND2x1p5_ASAP7_75t_L g3110 ( 
.A(n_2897),
.B(n_2498),
.Y(n_3110)
);

OAI221xp5_ASAP7_75t_L g3111 ( 
.A1(n_2880),
.A2(n_2962),
.B1(n_2968),
.B2(n_2849),
.C(n_2928),
.Y(n_3111)
);

OAI22xp5_ASAP7_75t_SL g3112 ( 
.A1(n_2704),
.A2(n_2598),
.B1(n_2503),
.B2(n_2531),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2777),
.Y(n_3113)
);

HB1xp67_ASAP7_75t_L g3114 ( 
.A(n_2871),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2778),
.Y(n_3115)
);

AO22x2_ASAP7_75t_L g3116 ( 
.A1(n_2754),
.A2(n_2547),
.B1(n_2520),
.B2(n_2601),
.Y(n_3116)
);

AO22x2_ASAP7_75t_L g3117 ( 
.A1(n_2762),
.A2(n_2520),
.B1(n_2443),
.B2(n_2424),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2857),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2949),
.Y(n_3119)
);

NAND2x1p5_ASAP7_75t_L g3120 ( 
.A(n_2949),
.B(n_2498),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2890),
.B(n_2503),
.Y(n_3121)
);

BUFx3_ASAP7_75t_L g3122 ( 
.A(n_2949),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2803),
.B(n_2598),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2859),
.Y(n_3124)
);

BUFx3_ASAP7_75t_L g3125 ( 
.A(n_2894),
.Y(n_3125)
);

INVx1_ASAP7_75t_SL g3126 ( 
.A(n_2720),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2744),
.B(n_2498),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2865),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2877),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2746),
.B(n_2535),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2748),
.B(n_2350),
.Y(n_3131)
);

AND2x4_ASAP7_75t_L g3132 ( 
.A(n_2721),
.B(n_2736),
.Y(n_3132)
);

HB1xp67_ASAP7_75t_L g3133 ( 
.A(n_2873),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2881),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2933),
.B(n_2535),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2882),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2888),
.Y(n_3137)
);

HB1xp67_ASAP7_75t_L g3138 ( 
.A(n_2873),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2917),
.Y(n_3139)
);

BUFx2_ASAP7_75t_L g3140 ( 
.A(n_2903),
.Y(n_3140)
);

AO22x2_ASAP7_75t_L g3141 ( 
.A1(n_2919),
.A2(n_2443),
.B1(n_2424),
.B2(n_2614),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2787),
.B(n_2535),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2889),
.Y(n_3143)
);

INVx2_ASAP7_75t_SL g3144 ( 
.A(n_2774),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2892),
.Y(n_3145)
);

OR2x2_ASAP7_75t_SL g3146 ( 
.A(n_2814),
.B(n_2361),
.Y(n_3146)
);

OAI221xp5_ASAP7_75t_L g3147 ( 
.A1(n_2880),
.A2(n_2602),
.B1(n_2650),
.B2(n_2509),
.C(n_2621),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2935),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2937),
.Y(n_3149)
);

HB1xp67_ASAP7_75t_L g3150 ( 
.A(n_2876),
.Y(n_3150)
);

INVxp67_ASAP7_75t_L g3151 ( 
.A(n_2714),
.Y(n_3151)
);

BUFx2_ASAP7_75t_L g3152 ( 
.A(n_2876),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2940),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2944),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2704),
.B(n_2361),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2945),
.B(n_2562),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2748),
.B(n_2660),
.Y(n_3157)
);

BUFx8_ASAP7_75t_L g3158 ( 
.A(n_2680),
.Y(n_3158)
);

INVxp67_ASAP7_75t_L g3159 ( 
.A(n_2714),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2965),
.Y(n_3160)
);

INVx8_ASAP7_75t_L g3161 ( 
.A(n_2915),
.Y(n_3161)
);

INVx3_ASAP7_75t_L g3162 ( 
.A(n_2689),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2843),
.B(n_2660),
.Y(n_3163)
);

AO22x2_ASAP7_75t_L g3164 ( 
.A1(n_2939),
.A2(n_2443),
.B1(n_2424),
.B2(n_2614),
.Y(n_3164)
);

AND2x6_ASAP7_75t_L g3165 ( 
.A(n_2862),
.B(n_2562),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2966),
.B(n_2817),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2858),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2911),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2855),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_2703),
.B(n_2503),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2946),
.Y(n_3171)
);

AND2x2_ASAP7_75t_SL g3172 ( 
.A(n_2962),
.B(n_2509),
.Y(n_3172)
);

OR2x6_ASAP7_75t_L g3173 ( 
.A(n_2915),
.B(n_2513),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2947),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2818),
.B(n_2562),
.Y(n_3175)
);

OAI221xp5_ASAP7_75t_L g3176 ( 
.A1(n_2968),
.A2(n_2610),
.B1(n_2589),
.B2(n_2659),
.C(n_2474),
.Y(n_3176)
);

OAI221xp5_ASAP7_75t_L g3177 ( 
.A1(n_2849),
.A2(n_2659),
.B1(n_2447),
.B2(n_2357),
.C(n_2651),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2872),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_2847),
.B(n_2563),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2851),
.B(n_2563),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2942),
.Y(n_3181)
);

AO22x2_ASAP7_75t_L g3182 ( 
.A1(n_2943),
.A2(n_2468),
.B1(n_2504),
.B2(n_2465),
.Y(n_3182)
);

INVxp33_ASAP7_75t_SL g3183 ( 
.A(n_2691),
.Y(n_3183)
);

AO22x2_ASAP7_75t_L g3184 ( 
.A1(n_2792),
.A2(n_2468),
.B1(n_2504),
.B2(n_2465),
.Y(n_3184)
);

CKINVDCx20_ASAP7_75t_R g3185 ( 
.A(n_2805),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2728),
.B(n_2513),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2789),
.B(n_2493),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_2810),
.B(n_2513),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2846),
.Y(n_3189)
);

HB1xp67_ASAP7_75t_L g3190 ( 
.A(n_2781),
.Y(n_3190)
);

AO22x2_ASAP7_75t_L g3191 ( 
.A1(n_2793),
.A2(n_2963),
.B1(n_2960),
.B2(n_2831),
.Y(n_3191)
);

AO22x2_ASAP7_75t_L g3192 ( 
.A1(n_2827),
.A2(n_2515),
.B1(n_2403),
.B2(n_2421),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2791),
.B(n_2493),
.Y(n_3193)
);

AO22x2_ASAP7_75t_L g3194 ( 
.A1(n_2755),
.A2(n_2515),
.B1(n_2403),
.B2(n_2421),
.Y(n_3194)
);

AO22x2_ASAP7_75t_L g3195 ( 
.A1(n_2707),
.A2(n_2429),
.B1(n_2446),
.B2(n_2323),
.Y(n_3195)
);

CKINVDCx10_ASAP7_75t_R g3196 ( 
.A(n_3008),
.Y(n_3196)
);

OAI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_3111),
.A2(n_2927),
.B(n_2875),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_3060),
.B(n_2781),
.Y(n_3198)
);

INVx2_ASAP7_75t_SL g3199 ( 
.A(n_3030),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_3085),
.A2(n_2813),
.B1(n_2810),
.B2(n_2951),
.Y(n_3200)
);

AOI22xp33_ASAP7_75t_L g3201 ( 
.A1(n_3013),
.A2(n_2813),
.B1(n_2853),
.B2(n_2928),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3166),
.B(n_2839),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_3125),
.A2(n_2951),
.B1(n_2839),
.B2(n_2845),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_3043),
.A2(n_2870),
.B(n_2932),
.Y(n_3204)
);

CKINVDCx10_ASAP7_75t_R g3205 ( 
.A(n_3071),
.Y(n_3205)
);

AOI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_3012),
.A2(n_2948),
.B(n_2938),
.Y(n_3206)
);

NOR2x1p5_ASAP7_75t_SL g3207 ( 
.A(n_3178),
.B(n_2812),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_3011),
.B(n_2692),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3147),
.A2(n_2518),
.B(n_2927),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2973),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2975),
.Y(n_3211)
);

BUFx6f_ASAP7_75t_L g3212 ( 
.A(n_3087),
.Y(n_3212)
);

NAND3xp33_ASAP7_75t_L g3213 ( 
.A(n_3070),
.B(n_2853),
.C(n_2901),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_3042),
.B(n_2684),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3137),
.B(n_2820),
.Y(n_3215)
);

A2O1A1Ixp33_ASAP7_75t_L g3216 ( 
.A1(n_3061),
.A2(n_2848),
.B(n_2929),
.C(n_2955),
.Y(n_3216)
);

AO21x1_ASAP7_75t_L g3217 ( 
.A1(n_2998),
.A2(n_2848),
.B(n_2828),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3002),
.B(n_2957),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3186),
.B(n_2929),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3021),
.B(n_2821),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_3093),
.B(n_2819),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3171),
.B(n_3174),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2990),
.B(n_2992),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_3188),
.B(n_2901),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2993),
.B(n_2794),
.Y(n_3225)
);

AOI21x1_ASAP7_75t_L g3226 ( 
.A1(n_3064),
.A2(n_2833),
.B(n_2874),
.Y(n_3226)
);

OR2x2_ASAP7_75t_L g3227 ( 
.A(n_3055),
.B(n_2868),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3176),
.A2(n_2694),
.B(n_2693),
.Y(n_3228)
);

CKINVDCx20_ASAP7_75t_R g3229 ( 
.A(n_3005),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_3177),
.A2(n_2696),
.B(n_2709),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2976),
.Y(n_3231)
);

INVxp67_ASAP7_75t_L g3232 ( 
.A(n_3152),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_3183),
.B(n_2845),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3139),
.B(n_2826),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_3035),
.B(n_2719),
.Y(n_3235)
);

OAI22xp5_ASAP7_75t_L g3236 ( 
.A1(n_3023),
.A2(n_2681),
.B1(n_2695),
.B2(n_2959),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_3187),
.A2(n_2711),
.B(n_2710),
.Y(n_3237)
);

OAI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3080),
.A2(n_2822),
.B(n_2852),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3193),
.A2(n_2727),
.B(n_2717),
.Y(n_3239)
);

BUFx6f_ASAP7_75t_L g3240 ( 
.A(n_3161),
.Y(n_3240)
);

NAND2x1p5_ASAP7_75t_L g3241 ( 
.A(n_3142),
.B(n_2964),
.Y(n_3241)
);

NAND3xp33_ASAP7_75t_L g3242 ( 
.A(n_2972),
.B(n_2955),
.C(n_2824),
.Y(n_3242)
);

OAI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_3000),
.A2(n_2854),
.B(n_2883),
.Y(n_3243)
);

A2O1A1Ixp33_ASAP7_75t_L g3244 ( 
.A1(n_3168),
.A2(n_2832),
.B(n_2967),
.C(n_2795),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_3189),
.A2(n_2732),
.B(n_2734),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3033),
.B(n_2826),
.Y(n_3246)
);

AOI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_3169),
.A2(n_2698),
.B(n_2430),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3167),
.A2(n_2430),
.B(n_2405),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3006),
.B(n_2824),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3143),
.B(n_2757),
.Y(n_3250)
);

A2O1A1Ixp33_ASAP7_75t_L g3251 ( 
.A1(n_3181),
.A2(n_2815),
.B(n_2840),
.C(n_2825),
.Y(n_3251)
);

XOR2x2_ASAP7_75t_R g3252 ( 
.A(n_3102),
.B(n_2961),
.Y(n_3252)
);

OAI21xp33_ASAP7_75t_L g3253 ( 
.A1(n_3145),
.A2(n_2763),
.B(n_2765),
.Y(n_3253)
);

NOR2xp67_ASAP7_75t_L g3254 ( 
.A(n_3026),
.B(n_2751),
.Y(n_3254)
);

BUFx2_ASAP7_75t_L g3255 ( 
.A(n_3007),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3016),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_3157),
.B(n_2796),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_3126),
.B(n_2850),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3063),
.A2(n_2510),
.B(n_2430),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3063),
.A2(n_2510),
.B(n_2430),
.Y(n_3260)
);

CKINVDCx10_ASAP7_75t_R g3261 ( 
.A(n_3071),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_3064),
.A2(n_2510),
.B(n_2651),
.Y(n_3262)
);

BUFx4f_ASAP7_75t_L g3263 ( 
.A(n_3132),
.Y(n_3263)
);

OAI22xp5_ASAP7_75t_L g3264 ( 
.A1(n_3088),
.A2(n_2773),
.B1(n_2766),
.B2(n_2920),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_L g3265 ( 
.A1(n_3013),
.A2(n_2802),
.B1(n_2761),
.B2(n_2958),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2977),
.Y(n_3266)
);

NOR2xp67_ASAP7_75t_L g3267 ( 
.A(n_3069),
.B(n_2689),
.Y(n_3267)
);

NOR2xp33_ASAP7_75t_L g3268 ( 
.A(n_3076),
.B(n_3098),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_3073),
.A2(n_2920),
.B1(n_2516),
.B2(n_2916),
.Y(n_3269)
);

BUFx2_ASAP7_75t_L g3270 ( 
.A(n_3001),
.Y(n_3270)
);

O2A1O1Ixp33_ASAP7_75t_L g3271 ( 
.A1(n_3144),
.A2(n_2861),
.B(n_2802),
.C(n_2749),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3127),
.A2(n_2510),
.B(n_2902),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3051),
.B(n_2885),
.Y(n_3273)
);

BUFx6f_ASAP7_75t_L g3274 ( 
.A(n_3161),
.Y(n_3274)
);

INVx2_ASAP7_75t_SL g3275 ( 
.A(n_2971),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3053),
.B(n_2895),
.Y(n_3276)
);

O2A1O1Ixp33_ASAP7_75t_L g3277 ( 
.A1(n_3123),
.A2(n_2869),
.B(n_2761),
.C(n_2884),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3130),
.A2(n_2907),
.B(n_2887),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3175),
.B(n_2863),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3163),
.B(n_2863),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_3025),
.A2(n_2462),
.B1(n_2439),
.B2(n_2867),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_3031),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2981),
.A2(n_2908),
.B(n_2909),
.Y(n_3283)
);

AOI221xp5_ASAP7_75t_L g3284 ( 
.A1(n_3191),
.A2(n_2733),
.B1(n_2936),
.B2(n_2784),
.C(n_2446),
.Y(n_3284)
);

NOR3xp33_ASAP7_75t_L g3285 ( 
.A(n_3179),
.B(n_2964),
.C(n_2936),
.Y(n_3285)
);

AOI31xp33_ASAP7_75t_L g3286 ( 
.A1(n_3155),
.A2(n_2841),
.A3(n_2812),
.B(n_2628),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_2981),
.A2(n_2924),
.B(n_2441),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3045),
.B(n_2784),
.Y(n_3288)
);

OAI21xp33_ASAP7_75t_L g3289 ( 
.A1(n_3191),
.A2(n_2429),
.B(n_2323),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2979),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2982),
.Y(n_3291)
);

OAI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3131),
.A2(n_2439),
.B(n_2462),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3151),
.B(n_2462),
.Y(n_3293)
);

BUFx6f_ASAP7_75t_L g3294 ( 
.A(n_3173),
.Y(n_3294)
);

OAI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3135),
.A2(n_2439),
.B(n_2462),
.Y(n_3295)
);

O2A1O1Ixp5_ASAP7_75t_L g3296 ( 
.A1(n_3074),
.A2(n_2440),
.B(n_2441),
.C(n_2638),
.Y(n_3296)
);

OAI22xp5_ASAP7_75t_L g3297 ( 
.A1(n_3050),
.A2(n_2516),
.B1(n_2788),
.B2(n_2729),
.Y(n_3297)
);

O2A1O1Ixp33_ASAP7_75t_L g3298 ( 
.A1(n_3159),
.A2(n_2647),
.B(n_2644),
.C(n_2462),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3036),
.Y(n_3299)
);

AOI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_3038),
.A2(n_3037),
.B(n_3156),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3190),
.B(n_2729),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_3038),
.A2(n_2841),
.B(n_2812),
.Y(n_3302)
);

A2O1A1Ixp33_ASAP7_75t_L g3303 ( 
.A1(n_3020),
.A2(n_2729),
.B(n_2788),
.C(n_2439),
.Y(n_3303)
);

OAI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3062),
.A2(n_2612),
.B(n_2439),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3037),
.A2(n_2841),
.B(n_2812),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3180),
.B(n_2788),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_3116),
.A2(n_2841),
.B(n_2812),
.Y(n_3307)
);

NOR2x1p5_ASAP7_75t_L g3308 ( 
.A(n_2988),
.B(n_2812),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3116),
.A2(n_2841),
.B(n_2612),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_3185),
.B(n_3172),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3039),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3022),
.A2(n_2841),
.B(n_2612),
.Y(n_3312)
);

AND2x2_ASAP7_75t_L g3313 ( 
.A(n_3089),
.B(n_21),
.Y(n_3313)
);

OAI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3046),
.A2(n_2612),
.B(n_22),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3047),
.B(n_2612),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_3067),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3114),
.B(n_22),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2984),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3022),
.A2(n_23),
.B(n_24),
.Y(n_3319)
);

CKINVDCx5p33_ASAP7_75t_R g3320 ( 
.A(n_2986),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3058),
.A2(n_3164),
.B(n_3141),
.Y(n_3321)
);

AOI21xp5_ASAP7_75t_L g3322 ( 
.A1(n_3058),
.A2(n_23),
.B(n_24),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3133),
.B(n_25),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3141),
.A2(n_25),
.B(n_26),
.Y(n_3324)
);

BUFx2_ASAP7_75t_SL g3325 ( 
.A(n_3009),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_3164),
.A2(n_26),
.B(n_27),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3004),
.A2(n_27),
.B(n_28),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3138),
.B(n_28),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2985),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3140),
.B(n_29),
.Y(n_3330)
);

NAND3xp33_ASAP7_75t_L g3331 ( 
.A(n_3150),
.B(n_29),
.C(n_30),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_2974),
.B(n_30),
.Y(n_3332)
);

OAI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_3056),
.A2(n_31),
.B(n_32),
.Y(n_3333)
);

INVx3_ASAP7_75t_L g3334 ( 
.A(n_3173),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3004),
.A2(n_31),
.B(n_32),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3048),
.A2(n_33),
.B(n_34),
.Y(n_3336)
);

HB1xp67_ASAP7_75t_L g3337 ( 
.A(n_2994),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3091),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_2989),
.B(n_35),
.Y(n_3339)
);

AOI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3048),
.A2(n_36),
.B(n_37),
.Y(n_3340)
);

OA22x2_ASAP7_75t_L g3341 ( 
.A1(n_3112),
.A2(n_3121),
.B1(n_3106),
.B2(n_3105),
.Y(n_3341)
);

A2O1A1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_2995),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_2989),
.A2(n_38),
.B(n_39),
.Y(n_3343)
);

O2A1O1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_2996),
.A2(n_701),
.B(n_702),
.C(n_700),
.Y(n_3344)
);

HB1xp67_ASAP7_75t_L g3345 ( 
.A(n_3052),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2997),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3034),
.B(n_40),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3195),
.A2(n_3103),
.B(n_3182),
.Y(n_3348)
);

O2A1O1Ixp33_ASAP7_75t_L g3349 ( 
.A1(n_2999),
.A2(n_702),
.B(n_43),
.C(n_41),
.Y(n_3349)
);

INVxp67_ASAP7_75t_L g3350 ( 
.A(n_3029),
.Y(n_3350)
);

BUFx12f_ASAP7_75t_L g3351 ( 
.A(n_3104),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3195),
.A2(n_41),
.B(n_42),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3003),
.Y(n_3353)
);

OAI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3072),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3354)
);

A2O1A1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_3015),
.A2(n_47),
.B(n_44),
.C(n_46),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3103),
.A2(n_46),
.B(n_47),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3182),
.A2(n_48),
.B(n_49),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3057),
.B(n_48),
.Y(n_3358)
);

OAI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3065),
.A2(n_49),
.B(n_50),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3034),
.B(n_3066),
.Y(n_3360)
);

INVx2_ASAP7_75t_SL g3361 ( 
.A(n_3083),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_3158),
.B(n_50),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3117),
.A2(n_51),
.B(n_52),
.Y(n_3363)
);

NOR2x1_ASAP7_75t_L g3364 ( 
.A(n_3077),
.B(n_694),
.Y(n_3364)
);

AOI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_3091),
.A2(n_3086),
.B1(n_3099),
.B2(n_3082),
.Y(n_3365)
);

AO21x1_ASAP7_75t_L g3366 ( 
.A1(n_3017),
.A2(n_51),
.B(n_52),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3068),
.B(n_53),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3079),
.B(n_3081),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3117),
.A2(n_53),
.B(n_54),
.Y(n_3369)
);

AOI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_3194),
.A2(n_54),
.B(n_55),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3084),
.B(n_55),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_2991),
.B(n_56),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3018),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3194),
.A2(n_56),
.B(n_58),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3090),
.B(n_58),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_SL g3376 ( 
.A(n_3165),
.B(n_59),
.Y(n_3376)
);

BUFx8_ASAP7_75t_SL g3377 ( 
.A(n_3122),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3019),
.Y(n_3378)
);

OAI22xp5_ASAP7_75t_L g3379 ( 
.A1(n_3146),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3146),
.B(n_61),
.Y(n_3380)
);

OAI21x1_ASAP7_75t_L g3381 ( 
.A1(n_3024),
.A2(n_62),
.B(n_63),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3027),
.Y(n_3382)
);

INVx2_ASAP7_75t_SL g3383 ( 
.A(n_3059),
.Y(n_3383)
);

BUFx3_ASAP7_75t_L g3384 ( 
.A(n_3119),
.Y(n_3384)
);

AO21x1_ASAP7_75t_L g3385 ( 
.A1(n_3028),
.A2(n_63),
.B(n_64),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_3170),
.B(n_65),
.Y(n_3386)
);

NAND2xp33_ASAP7_75t_SL g3387 ( 
.A(n_2987),
.B(n_66),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3094),
.B(n_66),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3096),
.B(n_67),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_2983),
.A2(n_67),
.B(n_70),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_2983),
.A2(n_70),
.B(n_71),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_2978),
.A2(n_74),
.B1(n_71),
.B2(n_72),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3054),
.A2(n_72),
.B(n_74),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3032),
.Y(n_3394)
);

BUFx6f_ASAP7_75t_L g3395 ( 
.A(n_3110),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3040),
.Y(n_3396)
);

NAND2x1p5_ASAP7_75t_L g3397 ( 
.A(n_3041),
.B(n_75),
.Y(n_3397)
);

A2O1A1Ixp33_ASAP7_75t_L g3398 ( 
.A1(n_3044),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3100),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3101),
.B(n_76),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3107),
.B(n_77),
.Y(n_3401)
);

BUFx12f_ASAP7_75t_L g3402 ( 
.A(n_3010),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3075),
.A2(n_78),
.B(n_79),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3108),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3109),
.Y(n_3405)
);

AND2x2_ASAP7_75t_SL g3406 ( 
.A(n_3376),
.B(n_3014),
.Y(n_3406)
);

A2O1A1Ixp33_ASAP7_75t_L g3407 ( 
.A1(n_3235),
.A2(n_3129),
.B(n_3134),
.C(n_3128),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_3268),
.B(n_3113),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3318),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3220),
.B(n_3099),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3209),
.A2(n_3014),
.B(n_3184),
.Y(n_3411)
);

NAND2x1p5_ASAP7_75t_L g3412 ( 
.A(n_3334),
.B(n_3162),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3223),
.B(n_3225),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3213),
.B(n_3097),
.Y(n_3414)
);

AOI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_3204),
.A2(n_3192),
.B(n_3184),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3213),
.B(n_3097),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3222),
.B(n_2978),
.Y(n_3417)
);

AND2x6_ASAP7_75t_L g3418 ( 
.A(n_3365),
.B(n_3115),
.Y(n_3418)
);

O2A1O1Ixp33_ASAP7_75t_L g3419 ( 
.A1(n_3216),
.A2(n_3124),
.B(n_3136),
.C(n_3118),
.Y(n_3419)
);

INVxp67_ASAP7_75t_L g3420 ( 
.A(n_3255),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3219),
.B(n_3086),
.Y(n_3421)
);

CKINVDCx5p33_ASAP7_75t_R g3422 ( 
.A(n_3196),
.Y(n_3422)
);

AOI222xp33_ASAP7_75t_L g3423 ( 
.A1(n_3201),
.A2(n_3102),
.B1(n_2980),
.B2(n_3082),
.C1(n_3165),
.C2(n_3078),
.Y(n_3423)
);

O2A1O1Ixp33_ASAP7_75t_L g3424 ( 
.A1(n_3379),
.A2(n_3154),
.B(n_3160),
.C(n_3153),
.Y(n_3424)
);

OAI22x1_ASAP7_75t_L g3425 ( 
.A1(n_3338),
.A2(n_2980),
.B1(n_3149),
.B2(n_3148),
.Y(n_3425)
);

NOR2xp33_ASAP7_75t_L g3426 ( 
.A(n_3233),
.B(n_3120),
.Y(n_3426)
);

BUFx6f_ASAP7_75t_L g3427 ( 
.A(n_3212),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_3264),
.B(n_3092),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_3212),
.Y(n_3429)
);

OAI22xp5_ASAP7_75t_L g3430 ( 
.A1(n_3242),
.A2(n_3078),
.B1(n_3192),
.B2(n_3095),
.Y(n_3430)
);

INVx6_ASAP7_75t_L g3431 ( 
.A(n_3212),
.Y(n_3431)
);

AOI21xp33_ASAP7_75t_L g3432 ( 
.A1(n_3242),
.A2(n_3049),
.B(n_3165),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_3377),
.Y(n_3433)
);

AND2x4_ASAP7_75t_L g3434 ( 
.A(n_3334),
.B(n_78),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_SL g3435 ( 
.A(n_3257),
.B(n_79),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3198),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3436)
);

O2A1O1Ixp33_ASAP7_75t_L g3437 ( 
.A1(n_3342),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_3437)
);

AND2x4_ASAP7_75t_L g3438 ( 
.A(n_3308),
.B(n_83),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3215),
.B(n_86),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_3206),
.A2(n_697),
.B(n_695),
.Y(n_3440)
);

O2A1O1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_3355),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3396),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3230),
.A2(n_701),
.B(n_699),
.Y(n_3443)
);

O2A1O1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_3398),
.A2(n_90),
.B(n_87),
.C(n_89),
.Y(n_3444)
);

OAI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_3251),
.A2(n_90),
.B(n_91),
.Y(n_3445)
);

NOR2x1_ASAP7_75t_R g3446 ( 
.A(n_3351),
.B(n_91),
.Y(n_3446)
);

A2O1A1Ixp33_ASAP7_75t_L g3447 ( 
.A1(n_3376),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_3447)
);

BUFx12f_ASAP7_75t_L g3448 ( 
.A(n_3320),
.Y(n_3448)
);

OAI22xp5_ASAP7_75t_SL g3449 ( 
.A1(n_3380),
.A2(n_95),
.B1(n_92),
.B2(n_94),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3246),
.B(n_95),
.Y(n_3450)
);

AOI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_3228),
.A2(n_688),
.B(n_687),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3214),
.A2(n_3339),
.B1(n_3221),
.B2(n_3347),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_3271),
.B(n_96),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3286),
.A2(n_689),
.B(n_688),
.Y(n_3454)
);

AO21x1_ASAP7_75t_L g3455 ( 
.A1(n_3392),
.A2(n_96),
.B(n_97),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3256),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3265),
.A2(n_100),
.B1(n_97),
.B2(n_98),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3211),
.Y(n_3458)
);

BUFx4f_ASAP7_75t_L g3459 ( 
.A(n_3240),
.Y(n_3459)
);

BUFx2_ASAP7_75t_L g3460 ( 
.A(n_3270),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_3200),
.B(n_100),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3249),
.B(n_102),
.Y(n_3462)
);

HB1xp67_ASAP7_75t_L g3463 ( 
.A(n_3279),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3282),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_3281),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_3465)
);

BUFx2_ASAP7_75t_L g3466 ( 
.A(n_3306),
.Y(n_3466)
);

NAND3xp33_ASAP7_75t_L g3467 ( 
.A(n_3331),
.B(n_103),
.C(n_104),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3286),
.A2(n_3197),
.B(n_3259),
.Y(n_3468)
);

BUFx16f_ASAP7_75t_R g3469 ( 
.A(n_3205),
.Y(n_3469)
);

INVx1_ASAP7_75t_SL g3470 ( 
.A(n_3301),
.Y(n_3470)
);

A2O1A1Ixp33_ASAP7_75t_L g3471 ( 
.A1(n_3253),
.A2(n_3277),
.B(n_3314),
.C(n_3197),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3299),
.Y(n_3472)
);

O2A1O1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_3333),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3260),
.A2(n_679),
.B(n_678),
.Y(n_3474)
);

NOR2x1_ASAP7_75t_SL g3475 ( 
.A(n_3325),
.B(n_105),
.Y(n_3475)
);

OR2x6_ASAP7_75t_SL g3476 ( 
.A(n_3203),
.B(n_106),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3224),
.B(n_107),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3202),
.B(n_3227),
.Y(n_3478)
);

NAND3xp33_ASAP7_75t_SL g3479 ( 
.A(n_3359),
.B(n_108),
.C(n_109),
.Y(n_3479)
);

INVx2_ASAP7_75t_SL g3480 ( 
.A(n_3263),
.Y(n_3480)
);

AO21x2_ASAP7_75t_L g3481 ( 
.A1(n_3262),
.A2(n_109),
.B(n_110),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_3243),
.A2(n_685),
.B(n_684),
.Y(n_3482)
);

BUFx6f_ASAP7_75t_L g3483 ( 
.A(n_3263),
.Y(n_3483)
);

OR2x6_ASAP7_75t_L g3484 ( 
.A(n_3341),
.B(n_111),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3234),
.A2(n_114),
.B1(n_111),
.B2(n_112),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3341),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3250),
.B(n_115),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3243),
.A2(n_694),
.B(n_693),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3311),
.Y(n_3489)
);

BUFx2_ASAP7_75t_SL g3490 ( 
.A(n_3254),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3316),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3238),
.A2(n_698),
.B(n_116),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3273),
.B(n_116),
.Y(n_3493)
);

BUFx8_ASAP7_75t_L g3494 ( 
.A(n_3383),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_R g3495 ( 
.A(n_3229),
.B(n_3361),
.Y(n_3495)
);

INVx1_ASAP7_75t_SL g3496 ( 
.A(n_3345),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3280),
.B(n_3208),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3247),
.A2(n_117),
.B(n_118),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3248),
.A2(n_118),
.B(n_119),
.Y(n_3499)
);

BUFx2_ASAP7_75t_L g3500 ( 
.A(n_3294),
.Y(n_3500)
);

AND2x4_ASAP7_75t_L g3501 ( 
.A(n_3285),
.B(n_119),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3310),
.B(n_121),
.Y(n_3502)
);

O2A1O1Ixp5_ASAP7_75t_L g3503 ( 
.A1(n_3217),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3294),
.B(n_122),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3218),
.B(n_123),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3278),
.A2(n_680),
.B(n_679),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3337),
.B(n_124),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3276),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3404),
.Y(n_3509)
);

OAI21xp33_ASAP7_75t_SL g3510 ( 
.A1(n_3284),
.A2(n_125),
.B(n_127),
.Y(n_3510)
);

O2A1O1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_3344),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3397),
.B(n_128),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3231),
.Y(n_3513)
);

AND2x4_ASAP7_75t_L g3514 ( 
.A(n_3294),
.B(n_130),
.Y(n_3514)
);

AND2x4_ASAP7_75t_L g3515 ( 
.A(n_3266),
.B(n_132),
.Y(n_3515)
);

AOI22xp33_ASAP7_75t_SL g3516 ( 
.A1(n_3331),
.A2(n_698),
.B1(n_692),
.B2(n_134),
.Y(n_3516)
);

INVx2_ASAP7_75t_SL g3517 ( 
.A(n_3261),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3245),
.A2(n_132),
.B(n_133),
.Y(n_3518)
);

OAI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3267),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_3519)
);

A2O1A1Ixp33_ASAP7_75t_L g3520 ( 
.A1(n_3343),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_3520)
);

AND2x4_ASAP7_75t_L g3521 ( 
.A(n_3290),
.B(n_138),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3405),
.Y(n_3522)
);

A2O1A1Ixp33_ASAP7_75t_L g3523 ( 
.A1(n_3327),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_3523)
);

OR2x6_ASAP7_75t_L g3524 ( 
.A(n_3402),
.B(n_139),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3237),
.A2(n_682),
.B(n_681),
.Y(n_3525)
);

OAI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3303),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3239),
.A2(n_3244),
.B(n_3302),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3291),
.Y(n_3528)
);

A2O1A1Ixp33_ASAP7_75t_L g3529 ( 
.A1(n_3335),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_3529)
);

AOI21xp5_ASAP7_75t_L g3530 ( 
.A1(n_3272),
.A2(n_692),
.B(n_690),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3258),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3307),
.A2(n_3305),
.B(n_3295),
.Y(n_3532)
);

BUFx3_ASAP7_75t_L g3533 ( 
.A(n_3240),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3210),
.Y(n_3534)
);

OAI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3232),
.A2(n_148),
.B1(n_145),
.B2(n_147),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3399),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3199),
.B(n_149),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3329),
.Y(n_3538)
);

AOI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3292),
.A2(n_150),
.B(n_151),
.Y(n_3539)
);

OR2x6_ASAP7_75t_L g3540 ( 
.A(n_3240),
.B(n_3274),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3312),
.A2(n_150),
.B(n_151),
.Y(n_3541)
);

NOR2xp33_ASAP7_75t_L g3542 ( 
.A(n_3386),
.B(n_152),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_R g3543 ( 
.A(n_3274),
.B(n_152),
.Y(n_3543)
);

HB1xp67_ASAP7_75t_L g3544 ( 
.A(n_3360),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3236),
.B(n_153),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3309),
.A2(n_154),
.B(n_155),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3269),
.B(n_3293),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3288),
.B(n_690),
.Y(n_3548)
);

BUFx2_ASAP7_75t_L g3549 ( 
.A(n_3384),
.Y(n_3549)
);

NAND2x1p5_ASAP7_75t_L g3550 ( 
.A(n_3274),
.B(n_154),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_3241),
.B(n_155),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3304),
.A2(n_3283),
.B(n_3298),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3346),
.Y(n_3553)
);

AOI21x1_ASAP7_75t_L g3554 ( 
.A1(n_3226),
.A2(n_156),
.B(n_157),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3304),
.A2(n_156),
.B(n_157),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3353),
.Y(n_3556)
);

NOR2xp33_ASAP7_75t_L g3557 ( 
.A(n_3372),
.B(n_158),
.Y(n_3557)
);

O2A1O1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3349),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3373),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3313),
.B(n_159),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3287),
.A2(n_160),
.B(n_161),
.Y(n_3561)
);

AOI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3354),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_3562)
);

A2O1A1Ixp33_ASAP7_75t_L g3563 ( 
.A1(n_3336),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_3563)
);

INVx8_ASAP7_75t_L g3564 ( 
.A(n_3395),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_R g3565 ( 
.A(n_3387),
.B(n_164),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3378),
.Y(n_3566)
);

AOI21x1_ASAP7_75t_L g3567 ( 
.A1(n_3319),
.A2(n_165),
.B(n_166),
.Y(n_3567)
);

NOR3xp33_ASAP7_75t_L g3568 ( 
.A(n_3340),
.B(n_167),
.C(n_168),
.Y(n_3568)
);

OAI22xp5_ASAP7_75t_L g3569 ( 
.A1(n_3241),
.A2(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_3569)
);

CKINVDCx20_ASAP7_75t_R g3570 ( 
.A(n_3350),
.Y(n_3570)
);

NOR2x1_ASAP7_75t_L g3571 ( 
.A(n_3364),
.B(n_169),
.Y(n_3571)
);

OAI21xp5_ASAP7_75t_L g3572 ( 
.A1(n_3322),
.A2(n_170),
.B(n_171),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_SL g3573 ( 
.A(n_3297),
.B(n_171),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3382),
.Y(n_3574)
);

AOI21x1_ASAP7_75t_L g3575 ( 
.A1(n_3300),
.A2(n_172),
.B(n_173),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3289),
.A2(n_3321),
.B(n_3296),
.Y(n_3576)
);

HB1xp67_ASAP7_75t_L g3577 ( 
.A(n_3394),
.Y(n_3577)
);

AOI21xp5_ASAP7_75t_L g3578 ( 
.A1(n_3348),
.A2(n_172),
.B(n_174),
.Y(n_3578)
);

BUFx6f_ASAP7_75t_L g3579 ( 
.A(n_3395),
.Y(n_3579)
);

O2A1O1Ixp33_ASAP7_75t_L g3580 ( 
.A1(n_3397),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3368),
.A2(n_176),
.B(n_177),
.Y(n_3581)
);

CKINVDCx20_ASAP7_75t_R g3582 ( 
.A(n_3275),
.Y(n_3582)
);

AOI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_3362),
.A2(n_3332),
.B1(n_3330),
.B2(n_3403),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3358),
.B(n_178),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3395),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3367),
.B(n_178),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3370),
.A2(n_179),
.B(n_180),
.Y(n_3587)
);

AOI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3393),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3374),
.A2(n_181),
.B(n_183),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3371),
.B(n_184),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3375),
.B(n_184),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3352),
.A2(n_185),
.B(n_186),
.Y(n_3592)
);

NAND3xp33_ASAP7_75t_SL g3593 ( 
.A(n_3366),
.B(n_187),
.C(n_188),
.Y(n_3593)
);

AOI221xp5_ASAP7_75t_L g3594 ( 
.A1(n_3385),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_3594)
);

INVx4_ASAP7_75t_L g3595 ( 
.A(n_3252),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_SL g3596 ( 
.A(n_3315),
.B(n_189),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3390),
.A2(n_190),
.B(n_191),
.Y(n_3597)
);

INVxp67_ASAP7_75t_L g3598 ( 
.A(n_3317),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3391),
.A2(n_191),
.B(n_192),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3388),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3324),
.A2(n_192),
.B(n_193),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3389),
.Y(n_3602)
);

O2A1O1Ixp33_ASAP7_75t_SL g3603 ( 
.A1(n_3400),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3326),
.A2(n_194),
.B(n_195),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3401),
.B(n_196),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_L g3606 ( 
.A(n_3323),
.B(n_197),
.Y(n_3606)
);

AO21x1_ASAP7_75t_L g3607 ( 
.A1(n_3363),
.A2(n_197),
.B(n_198),
.Y(n_3607)
);

INVx3_ASAP7_75t_L g3608 ( 
.A(n_3381),
.Y(n_3608)
);

INVx5_ASAP7_75t_L g3609 ( 
.A(n_3207),
.Y(n_3609)
);

INVx2_ASAP7_75t_SL g3610 ( 
.A(n_3328),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_3356),
.B(n_198),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3357),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3369),
.A2(n_199),
.B(n_200),
.Y(n_3613)
);

A2O1A1Ixp33_ASAP7_75t_L g3614 ( 
.A1(n_3235),
.A2(n_203),
.B(n_200),
.C(n_201),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3233),
.B(n_201),
.Y(n_3615)
);

AOI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3545),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_3616)
);

INVx3_ASAP7_75t_L g3617 ( 
.A(n_3579),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3409),
.Y(n_3618)
);

AOI21xp33_ASAP7_75t_L g3619 ( 
.A1(n_3471),
.A2(n_204),
.B(n_206),
.Y(n_3619)
);

OAI22xp5_ASAP7_75t_L g3620 ( 
.A1(n_3452),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_3620)
);

INVx5_ASAP7_75t_L g3621 ( 
.A(n_3608),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3556),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3442),
.Y(n_3623)
);

BUFx8_ASAP7_75t_L g3624 ( 
.A(n_3517),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3534),
.Y(n_3625)
);

BUFx6f_ASAP7_75t_L g3626 ( 
.A(n_3427),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3538),
.Y(n_3627)
);

AND2x2_ASAP7_75t_L g3628 ( 
.A(n_3466),
.B(n_686),
.Y(n_3628)
);

BUFx3_ASAP7_75t_L g3629 ( 
.A(n_3582),
.Y(n_3629)
);

INVx5_ASAP7_75t_L g3630 ( 
.A(n_3608),
.Y(n_3630)
);

BUFx2_ASAP7_75t_SL g3631 ( 
.A(n_3609),
.Y(n_3631)
);

HB1xp67_ASAP7_75t_L g3632 ( 
.A(n_3463),
.Y(n_3632)
);

INVx1_ASAP7_75t_SL g3633 ( 
.A(n_3549),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3566),
.Y(n_3634)
);

BUFx2_ASAP7_75t_L g3635 ( 
.A(n_3460),
.Y(n_3635)
);

BUFx6f_ASAP7_75t_L g3636 ( 
.A(n_3427),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3577),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3458),
.Y(n_3638)
);

OAI21xp33_ASAP7_75t_SL g3639 ( 
.A1(n_3595),
.A2(n_208),
.B(n_209),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3513),
.Y(n_3640)
);

AND2x4_ASAP7_75t_L g3641 ( 
.A(n_3574),
.B(n_210),
.Y(n_3641)
);

INVx6_ASAP7_75t_SL g3642 ( 
.A(n_3540),
.Y(n_3642)
);

CKINVDCx16_ASAP7_75t_R g3643 ( 
.A(n_3495),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3536),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3527),
.A2(n_211),
.B(n_212),
.Y(n_3645)
);

BUFx3_ASAP7_75t_L g3646 ( 
.A(n_3431),
.Y(n_3646)
);

BUFx6f_ASAP7_75t_L g3647 ( 
.A(n_3427),
.Y(n_3647)
);

INVx8_ASAP7_75t_L g3648 ( 
.A(n_3564),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3528),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3553),
.Y(n_3650)
);

CKINVDCx5p33_ASAP7_75t_R g3651 ( 
.A(n_3422),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3559),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3544),
.Y(n_3653)
);

INVx2_ASAP7_75t_SL g3654 ( 
.A(n_3431),
.Y(n_3654)
);

INVx3_ASAP7_75t_L g3655 ( 
.A(n_3579),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3417),
.Y(n_3656)
);

INVx1_ASAP7_75t_SL g3657 ( 
.A(n_3470),
.Y(n_3657)
);

AOI22xp5_ASAP7_75t_L g3658 ( 
.A1(n_3461),
.A2(n_3479),
.B1(n_3583),
.B2(n_3453),
.Y(n_3658)
);

AND2x4_ASAP7_75t_SL g3659 ( 
.A(n_3483),
.B(n_212),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3413),
.B(n_3497),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3509),
.Y(n_3661)
);

AND2x4_ASAP7_75t_L g3662 ( 
.A(n_3500),
.B(n_213),
.Y(n_3662)
);

INVx1_ASAP7_75t_SL g3663 ( 
.A(n_3496),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3522),
.Y(n_3664)
);

CKINVDCx5p33_ASAP7_75t_R g3665 ( 
.A(n_3433),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3414),
.Y(n_3666)
);

BUFx6f_ASAP7_75t_L g3667 ( 
.A(n_3429),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3421),
.B(n_213),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3456),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_3579),
.Y(n_3670)
);

BUFx2_ASAP7_75t_L g3671 ( 
.A(n_3420),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3416),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3429),
.Y(n_3673)
);

INVx1_ASAP7_75t_SL g3674 ( 
.A(n_3478),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3410),
.B(n_686),
.Y(n_3675)
);

NAND3xp33_ASAP7_75t_L g3676 ( 
.A(n_3492),
.B(n_214),
.C(n_215),
.Y(n_3676)
);

BUFx2_ASAP7_75t_L g3677 ( 
.A(n_3540),
.Y(n_3677)
);

AND2x4_ASAP7_75t_L g3678 ( 
.A(n_3585),
.B(n_215),
.Y(n_3678)
);

OR2x6_ASAP7_75t_L g3679 ( 
.A(n_3484),
.B(n_216),
.Y(n_3679)
);

BUFx2_ASAP7_75t_L g3680 ( 
.A(n_3533),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_3426),
.B(n_216),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3464),
.Y(n_3682)
);

AO22x1_ASAP7_75t_L g3683 ( 
.A1(n_3445),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_3683)
);

AND2x6_ASAP7_75t_L g3684 ( 
.A(n_3438),
.B(n_219),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3564),
.Y(n_3685)
);

AOI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3554),
.A2(n_220),
.B(n_221),
.Y(n_3686)
);

O2A1O1Ixp5_ASAP7_75t_L g3687 ( 
.A1(n_3482),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3472),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3610),
.B(n_222),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3489),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3406),
.B(n_684),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3600),
.B(n_223),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3491),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3575),
.Y(n_3694)
);

BUFx2_ASAP7_75t_L g3695 ( 
.A(n_3484),
.Y(n_3695)
);

BUFx6f_ASAP7_75t_L g3696 ( 
.A(n_3429),
.Y(n_3696)
);

BUFx8_ASAP7_75t_SL g3697 ( 
.A(n_3448),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3602),
.B(n_224),
.Y(n_3698)
);

BUFx2_ASAP7_75t_L g3699 ( 
.A(n_3418),
.Y(n_3699)
);

OR2x6_ASAP7_75t_L g3700 ( 
.A(n_3595),
.B(n_224),
.Y(n_3700)
);

INVx1_ASAP7_75t_SL g3701 ( 
.A(n_3490),
.Y(n_3701)
);

BUFx6f_ASAP7_75t_L g3702 ( 
.A(n_3483),
.Y(n_3702)
);

BUFx2_ASAP7_75t_SL g3703 ( 
.A(n_3609),
.Y(n_3703)
);

INVx1_ASAP7_75t_SL g3704 ( 
.A(n_3408),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3612),
.Y(n_3705)
);

BUFx3_ASAP7_75t_L g3706 ( 
.A(n_3494),
.Y(n_3706)
);

INVx1_ASAP7_75t_SL g3707 ( 
.A(n_3504),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3481),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3598),
.B(n_225),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_3407),
.B(n_225),
.Y(n_3710)
);

INVx3_ASAP7_75t_L g3711 ( 
.A(n_3483),
.Y(n_3711)
);

INVx3_ASAP7_75t_L g3712 ( 
.A(n_3412),
.Y(n_3712)
);

INVx3_ASAP7_75t_L g3713 ( 
.A(n_3438),
.Y(n_3713)
);

NOR2xp33_ASAP7_75t_SL g3714 ( 
.A(n_3480),
.B(n_226),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3609),
.Y(n_3715)
);

INVx5_ASAP7_75t_L g3716 ( 
.A(n_3501),
.Y(n_3716)
);

BUFx2_ASAP7_75t_R g3717 ( 
.A(n_3476),
.Y(n_3717)
);

AND2x2_ASAP7_75t_SL g3718 ( 
.A(n_3568),
.B(n_226),
.Y(n_3718)
);

AND2x4_ASAP7_75t_L g3719 ( 
.A(n_3501),
.B(n_227),
.Y(n_3719)
);

OAI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3562),
.A2(n_3588),
.B1(n_3467),
.B2(n_3486),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3419),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3450),
.B(n_227),
.Y(n_3722)
);

BUFx12f_ASAP7_75t_L g3723 ( 
.A(n_3494),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3515),
.Y(n_3724)
);

INVx1_ASAP7_75t_SL g3725 ( 
.A(n_3504),
.Y(n_3725)
);

OR2x6_ASAP7_75t_L g3726 ( 
.A(n_3454),
.B(n_228),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3432),
.B(n_228),
.Y(n_3727)
);

INVx4_ASAP7_75t_L g3728 ( 
.A(n_3459),
.Y(n_3728)
);

HB1xp67_ASAP7_75t_L g3729 ( 
.A(n_3425),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3468),
.A2(n_230),
.B(n_231),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3548),
.B(n_230),
.Y(n_3731)
);

AOI33xp33_ASAP7_75t_L g3732 ( 
.A1(n_3516),
.A2(n_234),
.A3(n_236),
.B1(n_231),
.B2(n_232),
.B3(n_235),
.Y(n_3732)
);

BUFx2_ASAP7_75t_L g3733 ( 
.A(n_3418),
.Y(n_3733)
);

BUFx6f_ASAP7_75t_L g3734 ( 
.A(n_3434),
.Y(n_3734)
);

BUFx6f_ASAP7_75t_L g3735 ( 
.A(n_3434),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3439),
.B(n_232),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3411),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3418),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_3570),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3515),
.B(n_683),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3487),
.B(n_234),
.Y(n_3741)
);

BUFx2_ASAP7_75t_L g3742 ( 
.A(n_3418),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3576),
.Y(n_3743)
);

OAI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3614),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_3744)
);

BUFx2_ASAP7_75t_L g3745 ( 
.A(n_3521),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3430),
.Y(n_3746)
);

OAI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3447),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_3747)
);

BUFx6f_ASAP7_75t_L g3748 ( 
.A(n_3514),
.Y(n_3748)
);

CKINVDCx5p33_ASAP7_75t_R g3749 ( 
.A(n_3543),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3521),
.Y(n_3750)
);

BUFx8_ASAP7_75t_L g3751 ( 
.A(n_3514),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_L g3752 ( 
.A(n_3502),
.B(n_238),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3567),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3415),
.Y(n_3754)
);

INVx1_ASAP7_75t_SL g3755 ( 
.A(n_3507),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3547),
.Y(n_3756)
);

BUFx2_ASAP7_75t_L g3757 ( 
.A(n_3524),
.Y(n_3757)
);

BUFx5_ASAP7_75t_L g3758 ( 
.A(n_3512),
.Y(n_3758)
);

A2O1A1Ixp33_ASAP7_75t_L g3759 ( 
.A1(n_3473),
.A2(n_3511),
.B(n_3558),
.C(n_3488),
.Y(n_3759)
);

INVx2_ASAP7_75t_SL g3760 ( 
.A(n_3524),
.Y(n_3760)
);

BUFx3_ASAP7_75t_L g3761 ( 
.A(n_3505),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3449),
.A2(n_242),
.B1(n_239),
.B2(n_241),
.Y(n_3762)
);

INVx5_ASAP7_75t_L g3763 ( 
.A(n_3607),
.Y(n_3763)
);

OR2x2_ASAP7_75t_SL g3764 ( 
.A(n_3593),
.B(n_243),
.Y(n_3764)
);

AND2x4_ASAP7_75t_L g3765 ( 
.A(n_3428),
.B(n_243),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3590),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3477),
.B(n_244),
.Y(n_3767)
);

BUFx6f_ASAP7_75t_L g3768 ( 
.A(n_3550),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3423),
.B(n_683),
.Y(n_3769)
);

AND2x4_ASAP7_75t_L g3770 ( 
.A(n_3532),
.B(n_245),
.Y(n_3770)
);

AOI221x1_ASAP7_75t_L g3771 ( 
.A1(n_3578),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3503),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3560),
.B(n_249),
.Y(n_3773)
);

INVx5_ASAP7_75t_L g3774 ( 
.A(n_3474),
.Y(n_3774)
);

A2O1A1Ixp33_ASAP7_75t_SL g3775 ( 
.A1(n_3572),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_L g3776 ( 
.A(n_3615),
.B(n_250),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3594),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3596),
.B(n_682),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3584),
.Y(n_3779)
);

BUFx3_ASAP7_75t_L g3780 ( 
.A(n_3537),
.Y(n_3780)
);

BUFx2_ASAP7_75t_SL g3781 ( 
.A(n_3551),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3586),
.B(n_254),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3455),
.Y(n_3783)
);

NOR2xp67_ASAP7_75t_L g3784 ( 
.A(n_3591),
.B(n_255),
.Y(n_3784)
);

AND2x4_ASAP7_75t_L g3785 ( 
.A(n_3552),
.B(n_3541),
.Y(n_3785)
);

AOI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3561),
.A2(n_255),
.B(n_256),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3443),
.A2(n_256),
.B(n_258),
.Y(n_3787)
);

BUFx2_ASAP7_75t_SL g3788 ( 
.A(n_3493),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3606),
.B(n_678),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3605),
.Y(n_3790)
);

AOI221xp5_ASAP7_75t_L g3791 ( 
.A1(n_3436),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.C(n_261),
.Y(n_3791)
);

INVx3_ASAP7_75t_L g3792 ( 
.A(n_3424),
.Y(n_3792)
);

NOR2x1_ASAP7_75t_R g3793 ( 
.A(n_3469),
.B(n_3435),
.Y(n_3793)
);

AOI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3557),
.A2(n_263),
.B1(n_260),
.B2(n_262),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3462),
.B(n_263),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3542),
.B(n_265),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_SL g3797 ( 
.A(n_3446),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3526),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_3798)
);

BUFx6f_ASAP7_75t_L g3799 ( 
.A(n_3573),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3451),
.A2(n_266),
.B(n_267),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3603),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3457),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_3802)
);

BUFx2_ASAP7_75t_L g3803 ( 
.A(n_3510),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3581),
.B(n_269),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3539),
.B(n_270),
.Y(n_3805)
);

HB1xp67_ASAP7_75t_L g3806 ( 
.A(n_3611),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3485),
.B(n_271),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3546),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3571),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3530),
.Y(n_3810)
);

OR2x2_ASAP7_75t_L g3811 ( 
.A(n_3506),
.B(n_271),
.Y(n_3811)
);

AOI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3508),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3498),
.Y(n_3813)
);

INVxp67_ASAP7_75t_SL g3814 ( 
.A(n_3525),
.Y(n_3814)
);

O2A1O1Ixp33_ASAP7_75t_L g3815 ( 
.A1(n_3520),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_3815)
);

INVx4_ASAP7_75t_L g3816 ( 
.A(n_3565),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3518),
.A2(n_275),
.B(n_276),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_SL g3818 ( 
.A(n_3580),
.B(n_276),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3475),
.B(n_3555),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3440),
.A2(n_277),
.B(n_278),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3563),
.Y(n_3821)
);

INVxp67_ASAP7_75t_L g3822 ( 
.A(n_3569),
.Y(n_3822)
);

INVx1_ASAP7_75t_SL g3823 ( 
.A(n_3499),
.Y(n_3823)
);

BUFx3_ASAP7_75t_L g3824 ( 
.A(n_3519),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3523),
.Y(n_3825)
);

AOI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_3531),
.A2(n_3535),
.B1(n_3465),
.B2(n_3529),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3597),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3592),
.Y(n_3828)
);

BUFx12f_ASAP7_75t_L g3829 ( 
.A(n_3601),
.Y(n_3829)
);

INVx3_ASAP7_75t_SL g3830 ( 
.A(n_3604),
.Y(n_3830)
);

CKINVDCx5p33_ASAP7_75t_R g3831 ( 
.A(n_3599),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_L g3832 ( 
.A1(n_3587),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3589),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3437),
.A2(n_3444),
.B(n_3441),
.Y(n_3834)
);

BUFx6f_ASAP7_75t_L g3835 ( 
.A(n_3613),
.Y(n_3835)
);

AOI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3545),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3409),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3409),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3556),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3463),
.B(n_284),
.Y(n_3840)
);

INVx1_ASAP7_75t_SL g3841 ( 
.A(n_3549),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3471),
.A2(n_285),
.B(n_286),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3635),
.B(n_3632),
.Y(n_3843)
);

BUFx2_ASAP7_75t_SL g3844 ( 
.A(n_3706),
.Y(n_3844)
);

OAI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3658),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_3845)
);

NAND2xp33_ASAP7_75t_L g3846 ( 
.A(n_3831),
.B(n_287),
.Y(n_3846)
);

AND2x4_ASAP7_75t_L g3847 ( 
.A(n_3622),
.B(n_288),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3627),
.Y(n_3848)
);

OR2x2_ASAP7_75t_L g3849 ( 
.A(n_3656),
.B(n_289),
.Y(n_3849)
);

INVx2_ASAP7_75t_SL g3850 ( 
.A(n_3633),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3638),
.Y(n_3851)
);

BUFx6f_ASAP7_75t_L g3852 ( 
.A(n_3626),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3634),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3710),
.A2(n_289),
.B(n_290),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3671),
.B(n_291),
.Y(n_3855)
);

AOI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3759),
.A2(n_291),
.B(n_292),
.Y(n_3856)
);

AND2x4_ASAP7_75t_L g3857 ( 
.A(n_3637),
.B(n_292),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3777),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3674),
.B(n_3666),
.Y(n_3859)
);

HB1xp67_ASAP7_75t_L g3860 ( 
.A(n_3839),
.Y(n_3860)
);

OAI22xp5_ASAP7_75t_L g3861 ( 
.A1(n_3679),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_3861)
);

AND2x6_ASAP7_75t_L g3862 ( 
.A(n_3770),
.B(n_296),
.Y(n_3862)
);

NAND2x1p5_ASAP7_75t_L g3863 ( 
.A(n_3657),
.B(n_296),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_SL g3864 ( 
.A(n_3643),
.B(n_297),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3644),
.Y(n_3865)
);

CKINVDCx20_ASAP7_75t_R g3866 ( 
.A(n_3651),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3640),
.Y(n_3867)
);

NOR2xp33_ASAP7_75t_L g3868 ( 
.A(n_3816),
.B(n_3793),
.Y(n_3868)
);

HAxp5_ASAP7_75t_L g3869 ( 
.A(n_3776),
.B(n_297),
.CON(n_3869),
.SN(n_3869)
);

AO21x2_ASAP7_75t_L g3870 ( 
.A1(n_3708),
.A2(n_298),
.B(n_299),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3653),
.B(n_298),
.Y(n_3871)
);

BUFx10_ASAP7_75t_L g3872 ( 
.A(n_3665),
.Y(n_3872)
);

BUFx6f_ASAP7_75t_L g3873 ( 
.A(n_3626),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3649),
.Y(n_3874)
);

AO22x2_ASAP7_75t_L g3875 ( 
.A1(n_3672),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3875)
);

NOR2xp33_ASAP7_75t_L g3876 ( 
.A(n_3816),
.B(n_301),
.Y(n_3876)
);

BUFx6f_ASAP7_75t_L g3877 ( 
.A(n_3626),
.Y(n_3877)
);

A2O1A1Ixp33_ASAP7_75t_SL g3878 ( 
.A1(n_3783),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3834),
.A2(n_303),
.B(n_304),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3660),
.B(n_305),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3818),
.A2(n_305),
.B(n_306),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3650),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3652),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3814),
.A2(n_306),
.B(n_307),
.Y(n_3884)
);

BUFx12f_ASAP7_75t_L g3885 ( 
.A(n_3739),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3704),
.B(n_308),
.Y(n_3886)
);

AOI221xp5_ASAP7_75t_L g3887 ( 
.A1(n_3842),
.A2(n_312),
.B1(n_308),
.B2(n_310),
.C(n_313),
.Y(n_3887)
);

OR2x2_ASAP7_75t_L g3888 ( 
.A(n_3737),
.B(n_312),
.Y(n_3888)
);

AOI22xp33_ASAP7_75t_L g3889 ( 
.A1(n_3829),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3625),
.B(n_314),
.Y(n_3890)
);

OR2x2_ASAP7_75t_L g3891 ( 
.A(n_3766),
.B(n_315),
.Y(n_3891)
);

CKINVDCx20_ASAP7_75t_R g3892 ( 
.A(n_3697),
.Y(n_3892)
);

BUFx6f_ASAP7_75t_L g3893 ( 
.A(n_3636),
.Y(n_3893)
);

AOI22xp33_ASAP7_75t_L g3894 ( 
.A1(n_3720),
.A2(n_319),
.B1(n_316),
.B2(n_318),
.Y(n_3894)
);

INVx3_ASAP7_75t_SL g3895 ( 
.A(n_3749),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3754),
.B(n_316),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3785),
.A2(n_3645),
.B(n_3683),
.Y(n_3897)
);

NOR2xp33_ASAP7_75t_L g3898 ( 
.A(n_3755),
.B(n_320),
.Y(n_3898)
);

INVx3_ASAP7_75t_L g3899 ( 
.A(n_3636),
.Y(n_3899)
);

AOI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_3785),
.A2(n_320),
.B(n_321),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3636),
.Y(n_3901)
);

BUFx2_ASAP7_75t_L g3902 ( 
.A(n_3758),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3661),
.B(n_321),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3775),
.A2(n_322),
.B(n_323),
.Y(n_3904)
);

INVx8_ASAP7_75t_L g3905 ( 
.A(n_3723),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3705),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3774),
.A2(n_322),
.B(n_324),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3664),
.B(n_324),
.Y(n_3908)
);

A2O1A1Ixp33_ASAP7_75t_L g3909 ( 
.A1(n_3732),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_3774),
.A2(n_325),
.B(n_327),
.Y(n_3910)
);

INVx5_ASAP7_75t_L g3911 ( 
.A(n_3684),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3690),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3618),
.Y(n_3913)
);

O2A1O1Ixp33_ASAP7_75t_L g3914 ( 
.A1(n_3744),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_3914)
);

INVxp67_ASAP7_75t_L g3915 ( 
.A(n_3790),
.Y(n_3915)
);

BUFx6f_ASAP7_75t_L g3916 ( 
.A(n_3647),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3746),
.B(n_329),
.Y(n_3917)
);

NOR2xp33_ASAP7_75t_L g3918 ( 
.A(n_3780),
.B(n_330),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3623),
.Y(n_3919)
);

CKINVDCx5p33_ASAP7_75t_R g3920 ( 
.A(n_3624),
.Y(n_3920)
);

INVxp33_ASAP7_75t_L g3921 ( 
.A(n_3629),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3837),
.Y(n_3922)
);

AOI22xp33_ASAP7_75t_SL g3923 ( 
.A1(n_3718),
.A2(n_677),
.B1(n_333),
.B2(n_331),
.Y(n_3923)
);

OR2x2_ASAP7_75t_SL g3924 ( 
.A(n_3729),
.B(n_3676),
.Y(n_3924)
);

OR2x6_ASAP7_75t_L g3925 ( 
.A(n_3770),
.B(n_331),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3756),
.B(n_332),
.Y(n_3926)
);

BUFx2_ASAP7_75t_SL g3927 ( 
.A(n_3701),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3838),
.B(n_334),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3779),
.B(n_335),
.Y(n_3929)
);

AOI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_3826),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3669),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3682),
.Y(n_3932)
);

OAI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_3730),
.A2(n_3800),
.B(n_3787),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3688),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_L g3935 ( 
.A1(n_3619),
.A2(n_339),
.B1(n_336),
.B2(n_337),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3663),
.B(n_3743),
.Y(n_3936)
);

AOI21xp5_ASAP7_75t_L g3937 ( 
.A1(n_3774),
.A2(n_340),
.B(n_341),
.Y(n_3937)
);

AND2x4_ASAP7_75t_L g3938 ( 
.A(n_3738),
.B(n_341),
.Y(n_3938)
);

NOR2xp67_ASAP7_75t_SL g3939 ( 
.A(n_3768),
.B(n_342),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3823),
.A2(n_342),
.B(n_344),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3693),
.B(n_3758),
.Y(n_3941)
);

NOR2xp33_ASAP7_75t_L g3942 ( 
.A(n_3761),
.B(n_345),
.Y(n_3942)
);

OAI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_3679),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3694),
.Y(n_3944)
);

AOI22xp5_ASAP7_75t_L g3945 ( 
.A1(n_3819),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3945)
);

AOI22xp33_ASAP7_75t_L g3946 ( 
.A1(n_3752),
.A2(n_3799),
.B1(n_3824),
.B2(n_3830),
.Y(n_3946)
);

INVx2_ASAP7_75t_SL g3947 ( 
.A(n_3841),
.Y(n_3947)
);

INVx2_ASAP7_75t_SL g3948 ( 
.A(n_3680),
.Y(n_3948)
);

A2O1A1Ixp33_ASAP7_75t_L g3949 ( 
.A1(n_3815),
.A2(n_350),
.B(n_348),
.C(n_349),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3715),
.Y(n_3950)
);

INVx2_ASAP7_75t_SL g3951 ( 
.A(n_3647),
.Y(n_3951)
);

INVx2_ASAP7_75t_SL g3952 ( 
.A(n_3647),
.Y(n_3952)
);

AOI21xp5_ASAP7_75t_L g3953 ( 
.A1(n_3721),
.A2(n_351),
.B(n_352),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3753),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3806),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3758),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3762),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3758),
.B(n_354),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3809),
.Y(n_3959)
);

OR2x2_ASAP7_75t_L g3960 ( 
.A(n_3745),
.B(n_354),
.Y(n_3960)
);

BUFx2_ASAP7_75t_L g3961 ( 
.A(n_3642),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3716),
.B(n_355),
.Y(n_3962)
);

BUFx6f_ASAP7_75t_L g3963 ( 
.A(n_3667),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3713),
.B(n_355),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3675),
.B(n_356),
.Y(n_3965)
);

BUFx3_ASAP7_75t_L g3966 ( 
.A(n_3624),
.Y(n_3966)
);

AOI21xp5_ASAP7_75t_L g3967 ( 
.A1(n_3810),
.A2(n_357),
.B(n_358),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3840),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3813),
.A2(n_360),
.B(n_361),
.Y(n_3969)
);

BUFx3_ASAP7_75t_L g3970 ( 
.A(n_3646),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3792),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3833),
.A2(n_360),
.B(n_362),
.Y(n_3972)
);

BUFx2_ASAP7_75t_R g3973 ( 
.A(n_3757),
.Y(n_3973)
);

INVx2_ASAP7_75t_SL g3974 ( 
.A(n_3667),
.Y(n_3974)
);

AOI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3808),
.A2(n_364),
.B(n_365),
.Y(n_3975)
);

O2A1O1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3747),
.A2(n_3805),
.B(n_3804),
.C(n_3807),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3817),
.A2(n_364),
.B(n_365),
.Y(n_3977)
);

O2A1O1Ixp33_ASAP7_75t_L g3978 ( 
.A1(n_3727),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_3978)
);

BUFx2_ASAP7_75t_R g3979 ( 
.A(n_3788),
.Y(n_3979)
);

NAND2xp33_ASAP7_75t_L g3980 ( 
.A(n_3684),
.B(n_366),
.Y(n_3980)
);

NOR2x1p5_ASAP7_75t_L g3981 ( 
.A(n_3728),
.B(n_367),
.Y(n_3981)
);

INVx3_ASAP7_75t_L g3982 ( 
.A(n_3667),
.Y(n_3982)
);

OR2x6_ASAP7_75t_SL g3983 ( 
.A(n_3796),
.B(n_368),
.Y(n_3983)
);

NOR2xp67_ASAP7_75t_L g3984 ( 
.A(n_3621),
.B(n_369),
.Y(n_3984)
);

CKINVDCx20_ASAP7_75t_R g3985 ( 
.A(n_3751),
.Y(n_3985)
);

BUFx6f_ASAP7_75t_L g3986 ( 
.A(n_3673),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3668),
.B(n_370),
.Y(n_3987)
);

INVx3_ASAP7_75t_SL g3988 ( 
.A(n_3648),
.Y(n_3988)
);

BUFx2_ASAP7_75t_L g3989 ( 
.A(n_3642),
.Y(n_3989)
);

BUFx5_ASAP7_75t_L g3990 ( 
.A(n_3684),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3792),
.B(n_370),
.Y(n_3991)
);

CKINVDCx5p33_ASAP7_75t_R g3992 ( 
.A(n_3797),
.Y(n_3992)
);

HB1xp67_ASAP7_75t_L g3993 ( 
.A(n_3699),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_3835),
.A2(n_371),
.B(n_372),
.Y(n_3994)
);

AOI222xp33_ASAP7_75t_L g3995 ( 
.A1(n_3791),
.A2(n_677),
.B1(n_375),
.B2(n_376),
.C1(n_377),
.C2(n_378),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3724),
.B(n_371),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3750),
.B(n_375),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3835),
.A2(n_376),
.B(n_378),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3733),
.Y(n_3999)
);

BUFx3_ASAP7_75t_L g4000 ( 
.A(n_3685),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3716),
.B(n_3799),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3695),
.B(n_379),
.Y(n_4002)
);

OR2x2_ASAP7_75t_L g4003 ( 
.A(n_3707),
.B(n_380),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3742),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3788),
.B(n_3722),
.Y(n_4005)
);

OA21x2_ASAP7_75t_L g4006 ( 
.A1(n_3772),
.A2(n_380),
.B(n_381),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3725),
.B(n_381),
.Y(n_4007)
);

BUFx12f_ASAP7_75t_L g4008 ( 
.A(n_3728),
.Y(n_4008)
);

AOI22xp5_ASAP7_75t_L g4009 ( 
.A1(n_3726),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3835),
.A2(n_382),
.B(n_384),
.Y(n_4010)
);

BUFx2_ASAP7_75t_L g4011 ( 
.A(n_3677),
.Y(n_4011)
);

AO21x1_ASAP7_75t_L g4012 ( 
.A1(n_3801),
.A2(n_385),
.B(n_387),
.Y(n_4012)
);

NAND2xp33_ASAP7_75t_L g4013 ( 
.A(n_3684),
.B(n_385),
.Y(n_4013)
);

BUFx2_ASAP7_75t_L g4014 ( 
.A(n_3713),
.Y(n_4014)
);

OAI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3616),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3734),
.B(n_388),
.Y(n_4016)
);

NAND2x1p5_ASAP7_75t_L g4017 ( 
.A(n_3716),
.B(n_389),
.Y(n_4017)
);

O2A1O1Ixp5_ASAP7_75t_L g4018 ( 
.A1(n_3687),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_3820),
.A2(n_390),
.B(n_391),
.Y(n_4019)
);

OAI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3726),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_4020)
);

AOI221x1_ASAP7_75t_L g4021 ( 
.A1(n_3620),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.C(n_396),
.Y(n_4021)
);

INVx3_ASAP7_75t_L g4022 ( 
.A(n_3673),
.Y(n_4022)
);

INVx3_ASAP7_75t_SL g4023 ( 
.A(n_3648),
.Y(n_4023)
);

INVx1_ASAP7_75t_SL g4024 ( 
.A(n_3971),
.Y(n_4024)
);

BUFx3_ASAP7_75t_L g4025 ( 
.A(n_3885),
.Y(n_4025)
);

BUFx12f_ASAP7_75t_L g4026 ( 
.A(n_3992),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3856),
.A2(n_3763),
.B1(n_3825),
.B2(n_3821),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3944),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3851),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3959),
.Y(n_4030)
);

OAI22xp33_ASAP7_75t_L g4031 ( 
.A1(n_3911),
.A2(n_3763),
.B1(n_3771),
.B2(n_3803),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3950),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3955),
.B(n_3763),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3867),
.Y(n_4034)
);

OAI21xp5_ASAP7_75t_SL g4035 ( 
.A1(n_3923),
.A2(n_3794),
.B(n_3812),
.Y(n_4035)
);

AOI22xp33_ASAP7_75t_L g4036 ( 
.A1(n_3980),
.A2(n_4013),
.B1(n_3933),
.B2(n_3846),
.Y(n_4036)
);

BUFx10_ASAP7_75t_L g4037 ( 
.A(n_3920),
.Y(n_4037)
);

INVx4_ASAP7_75t_L g4038 ( 
.A(n_3905),
.Y(n_4038)
);

OAI22xp33_ASAP7_75t_L g4039 ( 
.A1(n_3911),
.A2(n_3700),
.B1(n_3811),
.B2(n_3799),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_3874),
.Y(n_4040)
);

CKINVDCx11_ASAP7_75t_R g4041 ( 
.A(n_3892),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3882),
.Y(n_4042)
);

BUFx10_ASAP7_75t_L g4043 ( 
.A(n_3868),
.Y(n_4043)
);

AOI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_3887),
.A2(n_3798),
.B1(n_3769),
.B2(n_3691),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3883),
.Y(n_4045)
);

BUFx3_ASAP7_75t_L g4046 ( 
.A(n_3966),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3995),
.A2(n_3822),
.B1(n_3781),
.B2(n_3828),
.Y(n_4047)
);

CKINVDCx11_ASAP7_75t_R g4048 ( 
.A(n_3866),
.Y(n_4048)
);

BUFx3_ASAP7_75t_L g4049 ( 
.A(n_3905),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3954),
.Y(n_4050)
);

INVx3_ASAP7_75t_SL g4051 ( 
.A(n_3895),
.Y(n_4051)
);

BUFx6f_ASAP7_75t_L g4052 ( 
.A(n_3852),
.Y(n_4052)
);

BUFx2_ASAP7_75t_SL g4053 ( 
.A(n_3985),
.Y(n_4053)
);

INVx5_ASAP7_75t_L g4054 ( 
.A(n_3862),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3860),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3912),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3906),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3843),
.B(n_3734),
.Y(n_4058)
);

BUFx8_ASAP7_75t_L g4059 ( 
.A(n_4008),
.Y(n_4059)
);

BUFx12f_ASAP7_75t_L g4060 ( 
.A(n_3872),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3913),
.Y(n_4061)
);

OAI21xp5_ASAP7_75t_SL g4062 ( 
.A1(n_3894),
.A2(n_3836),
.B(n_3789),
.Y(n_4062)
);

OAI22xp33_ASAP7_75t_L g4063 ( 
.A1(n_3911),
.A2(n_3700),
.B1(n_3714),
.B2(n_3734),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3848),
.Y(n_4064)
);

OAI21xp5_ASAP7_75t_SL g4065 ( 
.A1(n_3930),
.A2(n_3767),
.B(n_3827),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3919),
.Y(n_4066)
);

CKINVDCx20_ASAP7_75t_R g4067 ( 
.A(n_3988),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3879),
.A2(n_3781),
.B1(n_3832),
.B2(n_3765),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3970),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3936),
.B(n_3709),
.Y(n_4070)
);

OAI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_4021),
.A2(n_3735),
.B1(n_3768),
.B2(n_3748),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3931),
.Y(n_4072)
);

OAI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_3909),
.A2(n_3717),
.B1(n_3764),
.B2(n_3802),
.Y(n_4073)
);

OAI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3897),
.A2(n_3639),
.B(n_3786),
.Y(n_4074)
);

CKINVDCx20_ASAP7_75t_R g4075 ( 
.A(n_4023),
.Y(n_4075)
);

BUFx6f_ASAP7_75t_L g4076 ( 
.A(n_3852),
.Y(n_4076)
);

OAI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3945),
.A2(n_3735),
.B1(n_3768),
.B2(n_3748),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3853),
.Y(n_4078)
);

HB1xp67_ASAP7_75t_L g4079 ( 
.A(n_3915),
.Y(n_4079)
);

AOI22xp33_ASAP7_75t_L g4080 ( 
.A1(n_3881),
.A2(n_3765),
.B1(n_3719),
.B2(n_3681),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3934),
.Y(n_4081)
);

INVx6_ASAP7_75t_L g4082 ( 
.A(n_3852),
.Y(n_4082)
);

AOI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_3862),
.A2(n_3719),
.B1(n_3760),
.B2(n_3773),
.Y(n_4083)
);

AOI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_3845),
.A2(n_3795),
.B1(n_3784),
.B2(n_3778),
.Y(n_4084)
);

OAI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_3925),
.A2(n_3735),
.B1(n_3748),
.B2(n_3712),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3865),
.Y(n_4086)
);

AOI22xp33_ASAP7_75t_L g4087 ( 
.A1(n_3862),
.A2(n_3751),
.B1(n_3741),
.B2(n_3736),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3922),
.Y(n_4088)
);

INVxp67_ASAP7_75t_SL g4089 ( 
.A(n_3941),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3977),
.A2(n_4019),
.B1(n_3858),
.B2(n_3990),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3932),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3990),
.A2(n_3731),
.B1(n_3641),
.B2(n_3782),
.Y(n_4092)
);

CKINVDCx20_ASAP7_75t_R g4093 ( 
.A(n_3961),
.Y(n_4093)
);

INVx4_ASAP7_75t_L g4094 ( 
.A(n_3925),
.Y(n_4094)
);

BUFx2_ASAP7_75t_L g4095 ( 
.A(n_3902),
.Y(n_4095)
);

OAI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_4009),
.A2(n_3712),
.B1(n_3702),
.B2(n_3711),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3859),
.Y(n_4097)
);

CKINVDCx20_ASAP7_75t_R g4098 ( 
.A(n_3989),
.Y(n_4098)
);

INVx3_ASAP7_75t_L g4099 ( 
.A(n_3956),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_4011),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3993),
.Y(n_4101)
);

BUFx10_ASAP7_75t_L g4102 ( 
.A(n_3876),
.Y(n_4102)
);

INVx1_ASAP7_75t_SL g4103 ( 
.A(n_3927),
.Y(n_4103)
);

AOI22xp33_ASAP7_75t_L g4104 ( 
.A1(n_3990),
.A2(n_3641),
.B1(n_3659),
.B2(n_3662),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4014),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3999),
.Y(n_4106)
);

AOI22xp33_ASAP7_75t_L g4107 ( 
.A1(n_3990),
.A2(n_3662),
.B1(n_3740),
.B2(n_3678),
.Y(n_4107)
);

INVx6_ASAP7_75t_L g4108 ( 
.A(n_3873),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_3948),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4004),
.Y(n_4110)
);

INVx4_ASAP7_75t_SL g4111 ( 
.A(n_3958),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3850),
.Y(n_4112)
);

NAND2x1p5_ASAP7_75t_L g4113 ( 
.A(n_4001),
.B(n_3621),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_4015),
.A2(n_3678),
.B1(n_3711),
.B2(n_3628),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_3947),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3968),
.Y(n_4116)
);

BUFx3_ASAP7_75t_L g4117 ( 
.A(n_4000),
.Y(n_4117)
);

INVx1_ASAP7_75t_SL g4118 ( 
.A(n_3973),
.Y(n_4118)
);

OAI22xp33_ASAP7_75t_L g4119 ( 
.A1(n_3900),
.A2(n_3702),
.B1(n_3686),
.B2(n_3698),
.Y(n_4119)
);

AOI22xp33_ASAP7_75t_L g4120 ( 
.A1(n_3935),
.A2(n_3702),
.B1(n_3631),
.B2(n_3703),
.Y(n_4120)
);

INVx2_ASAP7_75t_SL g4121 ( 
.A(n_3873),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_SL g4122 ( 
.A1(n_3875),
.A2(n_3703),
.B1(n_3631),
.B2(n_3689),
.Y(n_4122)
);

INVx6_ASAP7_75t_L g4123 ( 
.A(n_3873),
.Y(n_4123)
);

AOI22xp33_ASAP7_75t_SL g4124 ( 
.A1(n_3875),
.A2(n_3692),
.B1(n_3621),
.B2(n_3630),
.Y(n_4124)
);

INVx4_ASAP7_75t_L g4125 ( 
.A(n_4017),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_SL g4126 ( 
.A1(n_3957),
.A2(n_3630),
.B1(n_3655),
.B2(n_3617),
.Y(n_4126)
);

INVx1_ASAP7_75t_SL g4127 ( 
.A(n_3979),
.Y(n_4127)
);

BUFx2_ASAP7_75t_L g4128 ( 
.A(n_3899),
.Y(n_4128)
);

INVx6_ASAP7_75t_L g4129 ( 
.A(n_3877),
.Y(n_4129)
);

CKINVDCx20_ASAP7_75t_R g4130 ( 
.A(n_3844),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4006),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4006),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3871),
.Y(n_4133)
);

OAI22xp5_ASAP7_75t_SL g4134 ( 
.A1(n_3924),
.A2(n_3654),
.B1(n_3696),
.B2(n_3673),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_3949),
.A2(n_3655),
.B1(n_3670),
.B2(n_3617),
.Y(n_4135)
);

BUFx2_ASAP7_75t_SL g4136 ( 
.A(n_3984),
.Y(n_4136)
);

AOI22xp33_ASAP7_75t_L g4137 ( 
.A1(n_3904),
.A2(n_3884),
.B1(n_3953),
.B2(n_3940),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3903),
.Y(n_4138)
);

BUFx12f_ASAP7_75t_L g4139 ( 
.A(n_3981),
.Y(n_4139)
);

CKINVDCx11_ASAP7_75t_R g4140 ( 
.A(n_3983),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_3889),
.A2(n_3670),
.B1(n_3696),
.B2(n_3630),
.Y(n_4141)
);

OAI22xp33_ASAP7_75t_R g4142 ( 
.A1(n_3918),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3908),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_SL g4144 ( 
.A1(n_3870),
.A2(n_3696),
.B1(n_400),
.B2(n_398),
.Y(n_4144)
);

INVx1_ASAP7_75t_SL g4145 ( 
.A(n_4005),
.Y(n_4145)
);

INVx2_ASAP7_75t_SL g4146 ( 
.A(n_3877),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_3854),
.A2(n_401),
.B1(n_398),
.B2(n_399),
.Y(n_4147)
);

BUFx2_ASAP7_75t_L g4148 ( 
.A(n_3901),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3849),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3890),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3877),
.Y(n_4151)
);

CKINVDCx20_ASAP7_75t_R g4152 ( 
.A(n_3864),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3951),
.Y(n_4153)
);

BUFx3_ASAP7_75t_L g4154 ( 
.A(n_3893),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3952),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3891),
.Y(n_4156)
);

AOI22xp5_ASAP7_75t_L g4157 ( 
.A1(n_4020),
.A2(n_676),
.B1(n_403),
.B2(n_399),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3928),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3888),
.Y(n_4159)
);

INVx2_ASAP7_75t_SL g4160 ( 
.A(n_3893),
.Y(n_4160)
);

BUFx2_ASAP7_75t_L g4161 ( 
.A(n_3982),
.Y(n_4161)
);

AOI22xp33_ASAP7_75t_SL g4162 ( 
.A1(n_3861),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3974),
.Y(n_4163)
);

CKINVDCx20_ASAP7_75t_R g4164 ( 
.A(n_4016),
.Y(n_4164)
);

BUFx2_ASAP7_75t_SL g4165 ( 
.A(n_3847),
.Y(n_4165)
);

BUFx12f_ASAP7_75t_L g4166 ( 
.A(n_4003),
.Y(n_4166)
);

CKINVDCx20_ASAP7_75t_R g4167 ( 
.A(n_3987),
.Y(n_4167)
);

CKINVDCx20_ASAP7_75t_R g4168 ( 
.A(n_3855),
.Y(n_4168)
);

INVx1_ASAP7_75t_SL g4169 ( 
.A(n_3896),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_3847),
.Y(n_4170)
);

CKINVDCx11_ASAP7_75t_R g4171 ( 
.A(n_3893),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_4012),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_4172)
);

CKINVDCx20_ASAP7_75t_R g4173 ( 
.A(n_3965),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_SL g4174 ( 
.A1(n_3943),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4028),
.Y(n_4175)
);

OAI22xp33_ASAP7_75t_L g4176 ( 
.A1(n_4054),
.A2(n_3863),
.B1(n_3962),
.B2(n_3991),
.Y(n_4176)
);

AND2x4_ASAP7_75t_L g4177 ( 
.A(n_4111),
.B(n_4022),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_4024),
.Y(n_4178)
);

OAI21x1_ASAP7_75t_L g4179 ( 
.A1(n_4113),
.A2(n_3910),
.B(n_3907),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4050),
.Y(n_4180)
);

CKINVDCx5p33_ASAP7_75t_R g4181 ( 
.A(n_4041),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_4024),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4029),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4058),
.B(n_3921),
.Y(n_4184)
);

OAI21x1_ASAP7_75t_L g4185 ( 
.A1(n_4131),
.A2(n_3937),
.B(n_3994),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_4132),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_4145),
.B(n_3960),
.Y(n_4187)
);

AOI22xp33_ASAP7_75t_L g4188 ( 
.A1(n_4073),
.A2(n_3967),
.B1(n_3972),
.B2(n_3969),
.Y(n_4188)
);

BUFx2_ASAP7_75t_L g4189 ( 
.A(n_4130),
.Y(n_4189)
);

HB1xp67_ASAP7_75t_L g4190 ( 
.A(n_4079),
.Y(n_4190)
);

INVxp67_ASAP7_75t_L g4191 ( 
.A(n_4033),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_4169),
.Y(n_4192)
);

AO21x2_ASAP7_75t_L g4193 ( 
.A1(n_4031),
.A2(n_3878),
.B(n_4002),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4034),
.Y(n_4194)
);

AOI22xp33_ASAP7_75t_SL g4195 ( 
.A1(n_4054),
.A2(n_3942),
.B1(n_3898),
.B2(n_3998),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4040),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4045),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4030),
.Y(n_4198)
);

AOI22xp33_ASAP7_75t_L g4199 ( 
.A1(n_4073),
.A2(n_3975),
.B1(n_4010),
.B2(n_3946),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4145),
.B(n_3880),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4042),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4057),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4032),
.Y(n_4203)
);

AO22x1_ASAP7_75t_L g4204 ( 
.A1(n_4054),
.A2(n_3857),
.B1(n_3938),
.B2(n_3964),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4100),
.B(n_3857),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_4142),
.A2(n_4140),
.B1(n_4036),
.B2(n_4137),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_4056),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4061),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4066),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4072),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4081),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4116),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_4064),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4078),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4097),
.B(n_3886),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4055),
.Y(n_4216)
);

INVx3_ASAP7_75t_L g4217 ( 
.A(n_4099),
.Y(n_4217)
);

INVx4_ASAP7_75t_L g4218 ( 
.A(n_4038),
.Y(n_4218)
);

AOI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_4134),
.A2(n_3939),
.B1(n_3938),
.B2(n_3917),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4086),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_4150),
.B(n_3976),
.Y(n_4221)
);

AOI21x1_ASAP7_75t_L g4222 ( 
.A1(n_4070),
.A2(n_3926),
.B(n_3929),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4088),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_4158),
.B(n_3996),
.Y(n_4224)
);

OR2x2_ASAP7_75t_L g4225 ( 
.A(n_4169),
.B(n_4007),
.Y(n_4225)
);

BUFx4f_ASAP7_75t_SL g4226 ( 
.A(n_4026),
.Y(n_4226)
);

BUFx2_ASAP7_75t_L g4227 ( 
.A(n_4103),
.Y(n_4227)
);

INVx4_ASAP7_75t_L g4228 ( 
.A(n_4038),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4091),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4101),
.Y(n_4230)
);

OAI21x1_ASAP7_75t_L g4231 ( 
.A1(n_4099),
.A2(n_3997),
.B(n_4018),
.Y(n_4231)
);

AOI21x1_ASAP7_75t_L g4232 ( 
.A1(n_4138),
.A2(n_4143),
.B(n_4095),
.Y(n_4232)
);

INVx2_ASAP7_75t_SL g4233 ( 
.A(n_4037),
.Y(n_4233)
);

AO21x2_ASAP7_75t_L g4234 ( 
.A1(n_4074),
.A2(n_3914),
.B(n_3978),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4089),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4159),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4156),
.Y(n_4237)
);

BUFx2_ASAP7_75t_L g4238 ( 
.A(n_4103),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4133),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4149),
.Y(n_4240)
);

AOI22xp33_ASAP7_75t_L g4241 ( 
.A1(n_4027),
.A2(n_3869),
.B1(n_3963),
.B2(n_3916),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_4110),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4106),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4105),
.Y(n_4244)
);

HB1xp67_ASAP7_75t_L g4245 ( 
.A(n_4134),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4170),
.Y(n_4246)
);

INVx3_ASAP7_75t_L g4247 ( 
.A(n_4052),
.Y(n_4247)
);

INVx3_ASAP7_75t_L g4248 ( 
.A(n_4052),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4128),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4153),
.Y(n_4250)
);

AO21x2_ASAP7_75t_L g4251 ( 
.A1(n_4074),
.A2(n_3963),
.B(n_3916),
.Y(n_4251)
);

AOI22xp33_ASAP7_75t_L g4252 ( 
.A1(n_4162),
.A2(n_3963),
.B1(n_3986),
.B2(n_3916),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4148),
.B(n_3986),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4155),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_4112),
.B(n_3986),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4161),
.Y(n_4256)
);

OAI21x1_ASAP7_75t_L g4257 ( 
.A1(n_4163),
.A2(n_407),
.B(n_408),
.Y(n_4257)
);

OAI21x1_ASAP7_75t_L g4258 ( 
.A1(n_4109),
.A2(n_408),
.B(n_409),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_4115),
.B(n_410),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4121),
.Y(n_4260)
);

HB1xp67_ASAP7_75t_L g4261 ( 
.A(n_4111),
.Y(n_4261)
);

HB1xp67_ASAP7_75t_L g4262 ( 
.A(n_4052),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_4076),
.Y(n_4263)
);

HB1xp67_ASAP7_75t_L g4264 ( 
.A(n_4076),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4146),
.Y(n_4265)
);

BUFx2_ASAP7_75t_L g4266 ( 
.A(n_4093),
.Y(n_4266)
);

AO21x1_ASAP7_75t_SL g4267 ( 
.A1(n_4141),
.A2(n_410),
.B(n_411),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4151),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_4076),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4094),
.Y(n_4270)
);

OAI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_4035),
.A2(n_415),
.B1(n_412),
.B2(n_413),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4160),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4094),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4082),
.Y(n_4274)
);

BUFx3_ASAP7_75t_L g4275 ( 
.A(n_4059),
.Y(n_4275)
);

BUFx3_ASAP7_75t_L g4276 ( 
.A(n_4059),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4154),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4082),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_SL g4279 ( 
.A(n_4124),
.B(n_412),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4108),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4108),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4122),
.B(n_416),
.Y(n_4282)
);

INVx6_ASAP7_75t_L g4283 ( 
.A(n_4037),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4165),
.Y(n_4284)
);

HB1xp67_ASAP7_75t_L g4285 ( 
.A(n_4166),
.Y(n_4285)
);

INVx3_ASAP7_75t_L g4286 ( 
.A(n_4123),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4123),
.Y(n_4287)
);

HB1xp67_ASAP7_75t_L g4288 ( 
.A(n_4117),
.Y(n_4288)
);

HB1xp67_ASAP7_75t_L g4289 ( 
.A(n_4129),
.Y(n_4289)
);

OAI22xp33_ASAP7_75t_L g4290 ( 
.A1(n_4035),
.A2(n_420),
.B1(n_417),
.B2(n_418),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4129),
.Y(n_4291)
);

AOI22xp33_ASAP7_75t_SL g4292 ( 
.A1(n_4152),
.A2(n_420),
.B1(n_417),
.B2(n_418),
.Y(n_4292)
);

AOI22xp33_ASAP7_75t_L g4293 ( 
.A1(n_4174),
.A2(n_676),
.B1(n_423),
.B2(n_421),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4085),
.Y(n_4294)
);

AO21x2_ASAP7_75t_L g4295 ( 
.A1(n_4071),
.A2(n_421),
.B(n_422),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4039),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4136),
.Y(n_4297)
);

AOI22xp33_ASAP7_75t_L g4298 ( 
.A1(n_4044),
.A2(n_675),
.B1(n_424),
.B2(n_422),
.Y(n_4298)
);

OA21x2_ASAP7_75t_L g4299 ( 
.A1(n_4092),
.A2(n_423),
.B(n_424),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4069),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4125),
.Y(n_4301)
);

HB1xp67_ASAP7_75t_SL g4302 ( 
.A(n_4053),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4125),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4102),
.Y(n_4304)
);

HB1xp67_ASAP7_75t_L g4305 ( 
.A(n_4135),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4043),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4043),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4119),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4102),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4046),
.Y(n_4310)
);

OR2x2_ASAP7_75t_L g4311 ( 
.A(n_4118),
.B(n_425),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4171),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4047),
.B(n_425),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4135),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4098),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4096),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4168),
.Y(n_4317)
);

AOI22xp33_ASAP7_75t_L g4318 ( 
.A1(n_4044),
.A2(n_675),
.B1(n_428),
.B2(n_426),
.Y(n_4318)
);

BUFx3_ASAP7_75t_L g4319 ( 
.A(n_4067),
.Y(n_4319)
);

HB1xp67_ASAP7_75t_L g4320 ( 
.A(n_4118),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4164),
.Y(n_4321)
);

AO21x2_ASAP7_75t_L g4322 ( 
.A1(n_4305),
.A2(n_4063),
.B(n_4157),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4186),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4304),
.B(n_4127),
.Y(n_4324)
);

AND2x4_ASAP7_75t_L g4325 ( 
.A(n_4261),
.B(n_4270),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4192),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4192),
.Y(n_4327)
);

OR2x2_ASAP7_75t_L g4328 ( 
.A(n_4187),
.B(n_4127),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4180),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4304),
.B(n_4051),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4186),
.Y(n_4331)
);

OA21x2_ASAP7_75t_L g4332 ( 
.A1(n_4279),
.A2(n_4305),
.B(n_4245),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4208),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4227),
.B(n_4238),
.Y(n_4334)
);

OR2x2_ASAP7_75t_L g4335 ( 
.A(n_4225),
.B(n_4235),
.Y(n_4335)
);

BUFx2_ASAP7_75t_L g4336 ( 
.A(n_4261),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4270),
.B(n_4049),
.Y(n_4337)
);

AND2x4_ASAP7_75t_L g4338 ( 
.A(n_4273),
.B(n_4025),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4209),
.Y(n_4339)
);

OAI21x1_ASAP7_75t_L g4340 ( 
.A1(n_4232),
.A2(n_4083),
.B(n_4087),
.Y(n_4340)
);

AO21x2_ASAP7_75t_L g4341 ( 
.A1(n_4279),
.A2(n_4157),
.B(n_4077),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4211),
.Y(n_4342)
);

AND2x4_ASAP7_75t_L g4343 ( 
.A(n_4251),
.B(n_4075),
.Y(n_4343)
);

INVx2_ASAP7_75t_SL g4344 ( 
.A(n_4283),
.Y(n_4344)
);

OA21x2_ASAP7_75t_L g4345 ( 
.A1(n_4245),
.A2(n_4065),
.B(n_4090),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4210),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4273),
.B(n_4060),
.Y(n_4347)
);

HB1xp67_ASAP7_75t_L g4348 ( 
.A(n_4190),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4175),
.Y(n_4349)
);

AND2x4_ASAP7_75t_L g4350 ( 
.A(n_4297),
.B(n_4107),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4183),
.Y(n_4351)
);

AO21x2_ASAP7_75t_L g4352 ( 
.A1(n_4271),
.A2(n_4065),
.B(n_4084),
.Y(n_4352)
);

AO21x2_ASAP7_75t_L g4353 ( 
.A1(n_4271),
.A2(n_4084),
.B(n_4062),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4194),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_L g4355 ( 
.A(n_4221),
.B(n_4139),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4201),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4211),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4202),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4306),
.B(n_4126),
.Y(n_4359)
);

BUFx6f_ASAP7_75t_L g4360 ( 
.A(n_4275),
.Y(n_4360)
);

CKINVDCx20_ASAP7_75t_R g4361 ( 
.A(n_4181),
.Y(n_4361)
);

HB1xp67_ASAP7_75t_L g4362 ( 
.A(n_4190),
.Y(n_4362)
);

AND2x4_ASAP7_75t_SL g4363 ( 
.A(n_4320),
.B(n_4104),
.Y(n_4363)
);

INVx3_ASAP7_75t_L g4364 ( 
.A(n_4283),
.Y(n_4364)
);

INVxp67_ASAP7_75t_L g4365 ( 
.A(n_4295),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4207),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4212),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4307),
.B(n_4048),
.Y(n_4368)
);

HB1xp67_ASAP7_75t_L g4369 ( 
.A(n_4178),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4242),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4196),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4242),
.Y(n_4372)
);

NOR2xp33_ASAP7_75t_L g4373 ( 
.A(n_4320),
.B(n_4167),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4314),
.B(n_4144),
.Y(n_4374)
);

OR2x2_ASAP7_75t_L g4375 ( 
.A(n_4200),
.B(n_4114),
.Y(n_4375)
);

OAI21x1_ASAP7_75t_L g4376 ( 
.A1(n_4178),
.A2(n_4120),
.B(n_4080),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_4182),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4216),
.Y(n_4378)
);

INVx1_ASAP7_75t_SL g4379 ( 
.A(n_4302),
.Y(n_4379)
);

OR2x2_ASAP7_75t_L g4380 ( 
.A(n_4191),
.B(n_4308),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4316),
.B(n_4173),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4196),
.Y(n_4382)
);

OAI21x1_ASAP7_75t_L g4383 ( 
.A1(n_4182),
.A2(n_4068),
.B(n_4172),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4296),
.B(n_4062),
.Y(n_4384)
);

HB1xp67_ASAP7_75t_L g4385 ( 
.A(n_4251),
.Y(n_4385)
);

INVxp67_ASAP7_75t_R g4386 ( 
.A(n_4288),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_4197),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4197),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4236),
.Y(n_4389)
);

INVx2_ASAP7_75t_SL g4390 ( 
.A(n_4283),
.Y(n_4390)
);

OR2x2_ASAP7_75t_L g4391 ( 
.A(n_4215),
.B(n_4147),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4250),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4250),
.Y(n_4393)
);

INVx5_ASAP7_75t_L g4394 ( 
.A(n_4275),
.Y(n_4394)
);

AO21x2_ASAP7_75t_L g4395 ( 
.A1(n_4290),
.A2(n_426),
.B(n_427),
.Y(n_4395)
);

OR2x2_ASAP7_75t_L g4396 ( 
.A(n_4294),
.B(n_427),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4254),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4239),
.Y(n_4398)
);

INVx2_ASAP7_75t_L g4399 ( 
.A(n_4254),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_SL g4400 ( 
.A(n_4176),
.B(n_428),
.Y(n_4400)
);

OAI21x1_ASAP7_75t_L g4401 ( 
.A1(n_4217),
.A2(n_429),
.B(n_430),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_SL g4402 ( 
.A(n_4181),
.B(n_429),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4240),
.Y(n_4403)
);

HB1xp67_ASAP7_75t_L g4404 ( 
.A(n_4198),
.Y(n_4404)
);

AOI22xp33_ASAP7_75t_L g4405 ( 
.A1(n_4234),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4198),
.Y(n_4406)
);

HB1xp67_ASAP7_75t_L g4407 ( 
.A(n_4203),
.Y(n_4407)
);

INVx4_ASAP7_75t_L g4408 ( 
.A(n_4276),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4237),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4230),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4230),
.Y(n_4411)
);

OR2x6_ASAP7_75t_L g4412 ( 
.A(n_4204),
.B(n_431),
.Y(n_4412)
);

BUFx12f_ASAP7_75t_L g4413 ( 
.A(n_4276),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4203),
.Y(n_4414)
);

INVx3_ASAP7_75t_L g4415 ( 
.A(n_4177),
.Y(n_4415)
);

OA21x2_ASAP7_75t_L g4416 ( 
.A1(n_4206),
.A2(n_432),
.B(n_434),
.Y(n_4416)
);

HB1xp67_ASAP7_75t_L g4417 ( 
.A(n_4213),
.Y(n_4417)
);

BUFx2_ASAP7_75t_L g4418 ( 
.A(n_4177),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4213),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_4214),
.Y(n_4420)
);

HB1xp67_ASAP7_75t_L g4421 ( 
.A(n_4214),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4244),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4244),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_4312),
.Y(n_4424)
);

BUFx6f_ASAP7_75t_L g4425 ( 
.A(n_4218),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4303),
.B(n_434),
.Y(n_4426)
);

INVx3_ASAP7_75t_L g4427 ( 
.A(n_4177),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_SL g4428 ( 
.A(n_4176),
.B(n_673),
.Y(n_4428)
);

AO21x2_ASAP7_75t_L g4429 ( 
.A1(n_4290),
.A2(n_435),
.B(n_436),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4220),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4246),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4303),
.B(n_435),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4263),
.Y(n_4433)
);

AOI21x1_ASAP7_75t_L g4434 ( 
.A1(n_4285),
.A2(n_437),
.B(n_438),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_4263),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4309),
.B(n_438),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4262),
.Y(n_4437)
);

OA21x2_ASAP7_75t_L g4438 ( 
.A1(n_4206),
.A2(n_439),
.B(n_441),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4262),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4264),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_4264),
.Y(n_4441)
);

OAI21x1_ASAP7_75t_L g4442 ( 
.A1(n_4217),
.A2(n_441),
.B(n_442),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4289),
.B(n_443),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_4228),
.Y(n_4444)
);

INVx2_ASAP7_75t_SL g4445 ( 
.A(n_4312),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4269),
.Y(n_4446)
);

CKINVDCx5p33_ASAP7_75t_R g4447 ( 
.A(n_4319),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4223),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4229),
.Y(n_4449)
);

INVx1_ASAP7_75t_SL g4450 ( 
.A(n_4266),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4243),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4289),
.Y(n_4452)
);

INVx1_ASAP7_75t_SL g4453 ( 
.A(n_4189),
.Y(n_4453)
);

INVx3_ASAP7_75t_L g4454 ( 
.A(n_4228),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4269),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4224),
.Y(n_4456)
);

OR2x2_ASAP7_75t_L g4457 ( 
.A(n_4284),
.B(n_444),
.Y(n_4457)
);

OA21x2_ASAP7_75t_L g4458 ( 
.A1(n_4231),
.A2(n_445),
.B(n_446),
.Y(n_4458)
);

OAI21x1_ASAP7_75t_L g4459 ( 
.A1(n_4249),
.A2(n_4256),
.B(n_4301),
.Y(n_4459)
);

OAI21x1_ASAP7_75t_L g4460 ( 
.A1(n_4247),
.A2(n_445),
.B(n_446),
.Y(n_4460)
);

AOI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4285),
.A2(n_447),
.B(n_448),
.Y(n_4461)
);

HB1xp67_ASAP7_75t_L g4462 ( 
.A(n_4193),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_L g4463 ( 
.A(n_4218),
.B(n_4233),
.Y(n_4463)
);

INVx2_ASAP7_75t_SL g4464 ( 
.A(n_4319),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4288),
.Y(n_4465)
);

OAI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_4365),
.A2(n_4428),
.B(n_4400),
.Y(n_4466)
);

OAI22xp5_ASAP7_75t_SL g4467 ( 
.A1(n_4332),
.A2(n_4195),
.B1(n_4226),
.B2(n_4199),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4352),
.B(n_4193),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4348),
.Y(n_4469)
);

BUFx3_ASAP7_75t_L g4470 ( 
.A(n_4413),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4386),
.B(n_4286),
.Y(n_4471)
);

AO21x2_ASAP7_75t_L g4472 ( 
.A1(n_4462),
.A2(n_4282),
.B(n_4295),
.Y(n_4472)
);

NAND2xp33_ASAP7_75t_R g4473 ( 
.A(n_4332),
.B(n_4299),
.Y(n_4473)
);

A2O1A1Ixp33_ASAP7_75t_L g4474 ( 
.A1(n_4365),
.A2(n_4188),
.B(n_4219),
.C(n_4313),
.Y(n_4474)
);

INVx2_ASAP7_75t_SL g4475 ( 
.A(n_4394),
.Y(n_4475)
);

AND2x4_ASAP7_75t_L g4476 ( 
.A(n_4343),
.B(n_4218),
.Y(n_4476)
);

INVxp67_ASAP7_75t_L g4477 ( 
.A(n_4334),
.Y(n_4477)
);

OR2x2_ASAP7_75t_L g4478 ( 
.A(n_4380),
.B(n_4335),
.Y(n_4478)
);

AOI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4352),
.A2(n_4234),
.B1(n_4188),
.B2(n_4298),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4348),
.Y(n_4480)
);

AND2x4_ASAP7_75t_L g4481 ( 
.A(n_4343),
.B(n_4315),
.Y(n_4481)
);

INVxp67_ASAP7_75t_L g4482 ( 
.A(n_4373),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4343),
.B(n_4330),
.Y(n_4483)
);

INVx2_ASAP7_75t_L g4484 ( 
.A(n_4360),
.Y(n_4484)
);

AOI22xp5_ASAP7_75t_L g4485 ( 
.A1(n_4353),
.A2(n_4318),
.B1(n_4298),
.B2(n_4199),
.Y(n_4485)
);

AND2x4_ASAP7_75t_SL g4486 ( 
.A(n_4361),
.B(n_4315),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4347),
.B(n_4286),
.Y(n_4487)
);

INVx2_ASAP7_75t_SL g4488 ( 
.A(n_4394),
.Y(n_4488)
);

OA21x2_ASAP7_75t_L g4489 ( 
.A1(n_4462),
.A2(n_4278),
.B(n_4274),
.Y(n_4489)
);

INVx5_ASAP7_75t_L g4490 ( 
.A(n_4360),
.Y(n_4490)
);

AOI22xp5_ASAP7_75t_L g4491 ( 
.A1(n_4353),
.A2(n_4318),
.B1(n_4299),
.B2(n_4252),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4364),
.B(n_4274),
.Y(n_4492)
);

O2A1O1Ixp33_ASAP7_75t_SL g4493 ( 
.A1(n_4400),
.A2(n_4311),
.B(n_4317),
.C(n_4321),
.Y(n_4493)
);

OAI22xp5_ASAP7_75t_L g4494 ( 
.A1(n_4428),
.A2(n_4252),
.B1(n_4241),
.B2(n_4299),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4362),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4364),
.B(n_4278),
.Y(n_4496)
);

NAND3xp33_ASAP7_75t_L g4497 ( 
.A(n_4405),
.B(n_4292),
.C(n_4293),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4324),
.B(n_4280),
.Y(n_4498)
);

INVx5_ASAP7_75t_SL g4499 ( 
.A(n_4360),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4341),
.A2(n_4293),
.B1(n_4241),
.B2(n_4277),
.Y(n_4500)
);

NOR2xp33_ASAP7_75t_L g4501 ( 
.A(n_4413),
.B(n_4226),
.Y(n_4501)
);

AO32x2_ASAP7_75t_L g4502 ( 
.A1(n_4424),
.A2(n_4222),
.A3(n_4280),
.B1(n_4281),
.B2(n_4259),
.Y(n_4502)
);

BUFx3_ASAP7_75t_L g4503 ( 
.A(n_4361),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4418),
.B(n_4281),
.Y(n_4504)
);

O2A1O1Ixp33_ASAP7_75t_L g4505 ( 
.A1(n_4332),
.A2(n_4310),
.B(n_4321),
.C(n_4317),
.Y(n_4505)
);

AO32x2_ASAP7_75t_L g4506 ( 
.A1(n_4445),
.A2(n_4390),
.A3(n_4344),
.B1(n_4464),
.B2(n_4408),
.Y(n_4506)
);

HB1xp67_ASAP7_75t_L g4507 ( 
.A(n_4362),
.Y(n_4507)
);

A2O1A1Ixp33_ASAP7_75t_L g4508 ( 
.A1(n_4405),
.A2(n_4179),
.B(n_4185),
.C(n_4258),
.Y(n_4508)
);

AOI22xp33_ASAP7_75t_L g4509 ( 
.A1(n_4345),
.A2(n_4267),
.B1(n_4300),
.B2(n_4205),
.Y(n_4509)
);

NOR2xp33_ASAP7_75t_L g4510 ( 
.A(n_4408),
.B(n_4184),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4360),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4338),
.B(n_4253),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4431),
.Y(n_4513)
);

NOR2xp33_ASAP7_75t_L g4514 ( 
.A(n_4379),
.B(n_4287),
.Y(n_4514)
);

AOI221x1_ASAP7_75t_SL g4515 ( 
.A1(n_4374),
.A2(n_4291),
.B1(n_4272),
.B2(n_4268),
.C(n_4265),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4338),
.B(n_4247),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4345),
.B(n_4257),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4363),
.B(n_4248),
.Y(n_4518)
);

AND2x4_ASAP7_75t_L g4519 ( 
.A(n_4415),
.B(n_4248),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4363),
.B(n_4260),
.Y(n_4520)
);

AND2x2_ASAP7_75t_L g4521 ( 
.A(n_4337),
.B(n_4255),
.Y(n_4521)
);

AOI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_4341),
.A2(n_450),
.B1(n_447),
.B2(n_448),
.Y(n_4522)
);

BUFx3_ASAP7_75t_L g4523 ( 
.A(n_4394),
.Y(n_4523)
);

BUFx3_ASAP7_75t_L g4524 ( 
.A(n_4394),
.Y(n_4524)
);

OAI21xp5_ASAP7_75t_L g4525 ( 
.A1(n_4340),
.A2(n_450),
.B(n_451),
.Y(n_4525)
);

INVx3_ASAP7_75t_L g4526 ( 
.A(n_4415),
.Y(n_4526)
);

AO21x2_ASAP7_75t_L g4527 ( 
.A1(n_4385),
.A2(n_452),
.B(n_453),
.Y(n_4527)
);

AND2x4_ASAP7_75t_L g4528 ( 
.A(n_4427),
.B(n_4325),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4345),
.B(n_452),
.Y(n_4529)
);

NAND2xp33_ASAP7_75t_L g4530 ( 
.A(n_4447),
.B(n_454),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4430),
.Y(n_4531)
);

OAI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_4383),
.A2(n_454),
.B(n_455),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4427),
.Y(n_4533)
);

OR2x2_ASAP7_75t_L g4534 ( 
.A(n_4384),
.B(n_456),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4412),
.B(n_456),
.Y(n_4535)
);

AND2x2_ASAP7_75t_L g4536 ( 
.A(n_4412),
.B(n_457),
.Y(n_4536)
);

OAI211xp5_ASAP7_75t_L g4537 ( 
.A1(n_4416),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_4537)
);

AND2x2_ASAP7_75t_L g4538 ( 
.A(n_4412),
.B(n_458),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4430),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4465),
.B(n_459),
.Y(n_4540)
);

HB1xp67_ASAP7_75t_SL g4541 ( 
.A(n_4447),
.Y(n_4541)
);

BUFx2_ASAP7_75t_L g4542 ( 
.A(n_4336),
.Y(n_4542)
);

CKINVDCx5p33_ASAP7_75t_R g4543 ( 
.A(n_4453),
.Y(n_4543)
);

NOR2xp33_ASAP7_75t_L g4544 ( 
.A(n_4450),
.B(n_461),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4359),
.B(n_461),
.Y(n_4545)
);

AOI221xp5_ASAP7_75t_L g4546 ( 
.A1(n_4322),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.C(n_465),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4350),
.B(n_462),
.Y(n_4547)
);

AND2x4_ASAP7_75t_L g4548 ( 
.A(n_4325),
.B(n_672),
.Y(n_4548)
);

INVx3_ASAP7_75t_L g4549 ( 
.A(n_4425),
.Y(n_4549)
);

OR2x2_ASAP7_75t_L g4550 ( 
.A(n_4456),
.B(n_464),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4350),
.B(n_465),
.Y(n_4551)
);

OA21x2_ASAP7_75t_L g4552 ( 
.A1(n_4459),
.A2(n_466),
.B(n_467),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4368),
.B(n_466),
.Y(n_4553)
);

OR2x2_ASAP7_75t_L g4554 ( 
.A(n_4375),
.B(n_4326),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4329),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_4452),
.B(n_467),
.Y(n_4556)
);

OAI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_4376),
.A2(n_468),
.B(n_469),
.Y(n_4557)
);

O2A1O1Ixp33_ASAP7_75t_L g4558 ( 
.A1(n_4322),
.A2(n_471),
.B(n_469),
.C(n_470),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4333),
.Y(n_4559)
);

O2A1O1Ixp33_ASAP7_75t_L g4560 ( 
.A1(n_4402),
.A2(n_4438),
.B(n_4416),
.C(n_4429),
.Y(n_4560)
);

OR2x6_ASAP7_75t_L g4561 ( 
.A(n_4425),
.B(n_4416),
.Y(n_4561)
);

INVx8_ASAP7_75t_L g4562 ( 
.A(n_4425),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4463),
.B(n_470),
.Y(n_4563)
);

INVxp67_ASAP7_75t_L g4564 ( 
.A(n_4373),
.Y(n_4564)
);

OA21x2_ASAP7_75t_L g4565 ( 
.A1(n_4385),
.A2(n_471),
.B(n_472),
.Y(n_4565)
);

AO21x2_ASAP7_75t_L g4566 ( 
.A1(n_4437),
.A2(n_472),
.B(n_473),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4339),
.Y(n_4567)
);

A2O1A1Ixp33_ASAP7_75t_L g4568 ( 
.A1(n_4355),
.A2(n_476),
.B(n_474),
.C(n_475),
.Y(n_4568)
);

INVx5_ASAP7_75t_L g4569 ( 
.A(n_4425),
.Y(n_4569)
);

AO32x2_ASAP7_75t_L g4570 ( 
.A1(n_4328),
.A2(n_4451),
.A3(n_4327),
.B1(n_4440),
.B2(n_4441),
.Y(n_4570)
);

O2A1O1Ixp33_ASAP7_75t_L g4571 ( 
.A1(n_4438),
.A2(n_477),
.B(n_474),
.C(n_475),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4346),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4463),
.B(n_478),
.Y(n_4573)
);

OAI21xp5_ASAP7_75t_L g4574 ( 
.A1(n_4438),
.A2(n_479),
.B(n_480),
.Y(n_4574)
);

AOI22xp5_ASAP7_75t_L g4575 ( 
.A1(n_4395),
.A2(n_479),
.B1(n_480),
.B2(n_482),
.Y(n_4575)
);

NAND3xp33_ASAP7_75t_L g4576 ( 
.A(n_4458),
.B(n_482),
.C(n_483),
.Y(n_4576)
);

OAI22xp5_ASAP7_75t_L g4577 ( 
.A1(n_4391),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_4577)
);

AND2x2_ASAP7_75t_SL g4578 ( 
.A(n_4458),
.B(n_486),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4444),
.B(n_486),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4381),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_4580)
);

AOI21xp5_ASAP7_75t_L g4581 ( 
.A1(n_4395),
.A2(n_487),
.B(n_490),
.Y(n_4581)
);

OAI21xp5_ASAP7_75t_L g4582 ( 
.A1(n_4458),
.A2(n_4355),
.B(n_4434),
.Y(n_4582)
);

AND2x4_ASAP7_75t_L g4583 ( 
.A(n_4444),
.B(n_492),
.Y(n_4583)
);

AND2x4_ASAP7_75t_L g4584 ( 
.A(n_4454),
.B(n_492),
.Y(n_4584)
);

OAI21xp5_ASAP7_75t_L g4585 ( 
.A1(n_4461),
.A2(n_493),
.B(n_494),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4454),
.B(n_493),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4323),
.Y(n_4587)
);

AND2x2_ASAP7_75t_L g4588 ( 
.A(n_4439),
.B(n_494),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4433),
.B(n_495),
.Y(n_4589)
);

AND2x2_ASAP7_75t_L g4590 ( 
.A(n_4433),
.B(n_4435),
.Y(n_4590)
);

AND2x4_ASAP7_75t_L g4591 ( 
.A(n_4435),
.B(n_671),
.Y(n_4591)
);

OR2x2_ASAP7_75t_L g4592 ( 
.A(n_4396),
.B(n_495),
.Y(n_4592)
);

OA21x2_ASAP7_75t_L g4593 ( 
.A1(n_4323),
.A2(n_496),
.B(n_497),
.Y(n_4593)
);

OAI21xp5_ASAP7_75t_L g4594 ( 
.A1(n_4401),
.A2(n_497),
.B(n_498),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4446),
.B(n_499),
.Y(n_4595)
);

AOI22xp5_ASAP7_75t_L g4596 ( 
.A1(n_4429),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_4596)
);

AOI211xp5_ASAP7_75t_L g4597 ( 
.A1(n_4460),
.A2(n_4457),
.B(n_4442),
.C(n_4377),
.Y(n_4597)
);

OA21x2_ASAP7_75t_L g4598 ( 
.A1(n_4331),
.A2(n_500),
.B(n_501),
.Y(n_4598)
);

OA21x2_ASAP7_75t_L g4599 ( 
.A1(n_4331),
.A2(n_502),
.B(n_503),
.Y(n_4599)
);

CKINVDCx14_ASAP7_75t_R g4600 ( 
.A(n_4436),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4446),
.B(n_503),
.Y(n_4601)
);

HB1xp67_ASAP7_75t_L g4602 ( 
.A(n_4542),
.Y(n_4602)
);

AND2x4_ASAP7_75t_L g4603 ( 
.A(n_4528),
.B(n_4455),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4483),
.B(n_4481),
.Y(n_4604)
);

INVx3_ASAP7_75t_L g4605 ( 
.A(n_4528),
.Y(n_4605)
);

OR2x2_ASAP7_75t_L g4606 ( 
.A(n_4478),
.B(n_4554),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4481),
.B(n_4455),
.Y(n_4607)
);

BUFx3_ASAP7_75t_L g4608 ( 
.A(n_4503),
.Y(n_4608)
);

INVx2_ASAP7_75t_SL g4609 ( 
.A(n_4490),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4512),
.B(n_4443),
.Y(n_4610)
);

OR2x2_ASAP7_75t_L g4611 ( 
.A(n_4482),
.B(n_4369),
.Y(n_4611)
);

OR2x2_ASAP7_75t_L g4612 ( 
.A(n_4564),
.B(n_4369),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4506),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4507),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4471),
.B(n_4377),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4506),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4542),
.Y(n_4617)
);

AND2x4_ASAP7_75t_L g4618 ( 
.A(n_4569),
.B(n_4422),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4516),
.B(n_4426),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4487),
.B(n_4432),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4469),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4480),
.Y(n_4622)
);

HB1xp67_ASAP7_75t_L g4623 ( 
.A(n_4565),
.Y(n_4623)
);

INVxp67_ASAP7_75t_L g4624 ( 
.A(n_4541),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4498),
.B(n_4518),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_4470),
.Y(n_4626)
);

INVx1_ASAP7_75t_SL g4627 ( 
.A(n_4486),
.Y(n_4627)
);

BUFx2_ASAP7_75t_L g4628 ( 
.A(n_4506),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4495),
.Y(n_4629)
);

AOI22xp33_ASAP7_75t_L g4630 ( 
.A1(n_4467),
.A2(n_4378),
.B1(n_4449),
.B2(n_4448),
.Y(n_4630)
);

HB1xp67_ASAP7_75t_L g4631 ( 
.A(n_4565),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4492),
.B(n_4389),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4531),
.Y(n_4633)
);

HB1xp67_ASAP7_75t_L g4634 ( 
.A(n_4473),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4539),
.Y(n_4635)
);

OR2x2_ASAP7_75t_L g4636 ( 
.A(n_4477),
.B(n_4398),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4513),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4489),
.Y(n_4638)
);

BUFx3_ASAP7_75t_L g4639 ( 
.A(n_4490),
.Y(n_4639)
);

AND2x4_ASAP7_75t_L g4640 ( 
.A(n_4569),
.B(n_4422),
.Y(n_4640)
);

BUFx2_ASAP7_75t_SL g4641 ( 
.A(n_4490),
.Y(n_4641)
);

HB1xp67_ASAP7_75t_L g4642 ( 
.A(n_4468),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4476),
.B(n_4504),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4476),
.B(n_4484),
.Y(n_4644)
);

INVx5_ASAP7_75t_L g4645 ( 
.A(n_4499),
.Y(n_4645)
);

HB1xp67_ASAP7_75t_L g4646 ( 
.A(n_4489),
.Y(n_4646)
);

OR2x2_ASAP7_75t_L g4647 ( 
.A(n_4517),
.B(n_4403),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4555),
.Y(n_4648)
);

BUFx2_ASAP7_75t_L g4649 ( 
.A(n_4543),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4522),
.B(n_4409),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4526),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4526),
.Y(n_4652)
);

BUFx10_ASAP7_75t_L g4653 ( 
.A(n_4501),
.Y(n_4653)
);

INVx3_ASAP7_75t_L g4654 ( 
.A(n_4523),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4559),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_4524),
.Y(n_4656)
);

AND2x2_ASAP7_75t_L g4657 ( 
.A(n_4511),
.B(n_4392),
.Y(n_4657)
);

INVx3_ASAP7_75t_L g4658 ( 
.A(n_4499),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4567),
.Y(n_4659)
);

AO21x2_ASAP7_75t_L g4660 ( 
.A1(n_4466),
.A2(n_4407),
.B(n_4404),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4475),
.Y(n_4661)
);

OR2x2_ASAP7_75t_L g4662 ( 
.A(n_4534),
.B(n_4349),
.Y(n_4662)
);

BUFx2_ASAP7_75t_L g4663 ( 
.A(n_4488),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4569),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4548),
.Y(n_4665)
);

OAI322xp33_ASAP7_75t_L g4666 ( 
.A1(n_4479),
.A2(n_4366),
.A3(n_4351),
.B1(n_4354),
.B2(n_4356),
.C1(n_4358),
.C2(n_4367),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4496),
.B(n_4392),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4515),
.B(n_4393),
.Y(n_4668)
);

INVxp67_ASAP7_75t_SL g4669 ( 
.A(n_4560),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4520),
.B(n_4393),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4548),
.Y(n_4671)
);

INVx2_ASAP7_75t_SL g4672 ( 
.A(n_4562),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4572),
.Y(n_4673)
);

CKINVDCx8_ASAP7_75t_R g4674 ( 
.A(n_4583),
.Y(n_4674)
);

INVx8_ASAP7_75t_L g4675 ( 
.A(n_4562),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4546),
.B(n_4397),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4601),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4589),
.Y(n_4678)
);

BUFx6f_ASAP7_75t_L g4679 ( 
.A(n_4583),
.Y(n_4679)
);

HB1xp67_ASAP7_75t_L g4680 ( 
.A(n_4527),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4485),
.B(n_4397),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4595),
.Y(n_4682)
);

BUFx2_ASAP7_75t_L g4683 ( 
.A(n_4570),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4519),
.B(n_4399),
.Y(n_4684)
);

AOI221xp5_ASAP7_75t_L g4685 ( 
.A1(n_4558),
.A2(n_4414),
.B1(n_4410),
.B2(n_4411),
.C(n_4370),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4587),
.Y(n_4686)
);

BUFx2_ASAP7_75t_L g4687 ( 
.A(n_4570),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4533),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4593),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4521),
.B(n_4399),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4514),
.B(n_4423),
.Y(n_4691)
);

INVx2_ASAP7_75t_L g4692 ( 
.A(n_4570),
.Y(n_4692)
);

BUFx6f_ASAP7_75t_L g4693 ( 
.A(n_4584),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4552),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4510),
.B(n_4423),
.Y(n_4695)
);

BUFx4f_ASAP7_75t_L g4696 ( 
.A(n_4584),
.Y(n_4696)
);

HB1xp67_ASAP7_75t_L g4697 ( 
.A(n_4552),
.Y(n_4697)
);

OR2x2_ASAP7_75t_L g4698 ( 
.A(n_4472),
.B(n_4406),
.Y(n_4698)
);

OR2x2_ASAP7_75t_L g4699 ( 
.A(n_4500),
.B(n_4406),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4600),
.B(n_4371),
.Y(n_4700)
);

NOR2xp33_ASAP7_75t_L g4701 ( 
.A(n_4493),
.B(n_4372),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4593),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4598),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4547),
.B(n_4371),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4551),
.B(n_4382),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4519),
.B(n_4382),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4669),
.B(n_4474),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4669),
.B(n_4529),
.Y(n_4708)
);

OAI221xp5_ASAP7_75t_SL g4709 ( 
.A1(n_4630),
.A2(n_4491),
.B1(n_4505),
.B2(n_4497),
.C(n_4596),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4608),
.B(n_4545),
.Y(n_4710)
);

AOI221xp5_ASAP7_75t_L g4711 ( 
.A1(n_4666),
.A2(n_4494),
.B1(n_4582),
.B2(n_4532),
.C(n_4574),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4608),
.B(n_4578),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4604),
.B(n_4549),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4604),
.B(n_4561),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4617),
.B(n_4535),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4627),
.B(n_4561),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4665),
.B(n_4536),
.Y(n_4717)
);

OAI221xp5_ASAP7_75t_L g4718 ( 
.A1(n_4630),
.A2(n_4525),
.B1(n_4557),
.B2(n_4508),
.C(n_4575),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4649),
.B(n_4563),
.Y(n_4719)
);

NAND3xp33_ASAP7_75t_L g4720 ( 
.A(n_4680),
.B(n_4634),
.C(n_4683),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4643),
.B(n_4573),
.Y(n_4721)
);

NAND2xp5_ASAP7_75t_L g4722 ( 
.A(n_4665),
.B(n_4538),
.Y(n_4722)
);

NAND2xp33_ASAP7_75t_SL g4723 ( 
.A(n_4680),
.B(n_4566),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4643),
.B(n_4553),
.Y(n_4724)
);

NAND3xp33_ASAP7_75t_L g4725 ( 
.A(n_4634),
.B(n_4576),
.C(n_4530),
.Y(n_4725)
);

OAI21xp33_ASAP7_75t_SL g4726 ( 
.A1(n_4623),
.A2(n_4509),
.B(n_4590),
.Y(n_4726)
);

OAI21xp33_ASAP7_75t_SL g4727 ( 
.A1(n_4623),
.A2(n_4585),
.B(n_4502),
.Y(n_4727)
);

OAI22xp5_ASAP7_75t_L g4728 ( 
.A1(n_4687),
.A2(n_4581),
.B1(n_4537),
.B2(n_4597),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4625),
.B(n_4579),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4610),
.B(n_4586),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_SL g4731 ( 
.A(n_4628),
.B(n_4571),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4671),
.B(n_4663),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4615),
.B(n_4588),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4671),
.B(n_4591),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4661),
.B(n_4591),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_L g4736 ( 
.A(n_4624),
.B(n_4556),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4700),
.B(n_4544),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4661),
.B(n_4540),
.Y(n_4738)
);

OAI21xp5_ASAP7_75t_SL g4739 ( 
.A1(n_4676),
.A2(n_4568),
.B(n_4580),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4704),
.B(n_4550),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4605),
.B(n_4502),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4605),
.B(n_4502),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_4626),
.B(n_4592),
.Y(n_4743)
);

NAND3xp33_ASAP7_75t_L g4744 ( 
.A(n_4631),
.B(n_4577),
.C(n_4594),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4705),
.B(n_4598),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_SL g4746 ( 
.A(n_4631),
.B(n_4404),
.Y(n_4746)
);

AOI22xp33_ASAP7_75t_SL g4747 ( 
.A1(n_4697),
.A2(n_4599),
.B1(n_4421),
.B2(n_4417),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4602),
.B(n_4599),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4602),
.B(n_4407),
.Y(n_4749)
);

OAI21xp5_ASAP7_75t_SL g4750 ( 
.A1(n_4650),
.A2(n_4421),
.B(n_4417),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4677),
.B(n_4387),
.Y(n_4751)
);

AOI221xp5_ASAP7_75t_L g4752 ( 
.A1(n_4668),
.A2(n_4701),
.B1(n_4681),
.B2(n_4697),
.C(n_4692),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4620),
.B(n_4387),
.Y(n_4753)
);

OAI21xp5_ASAP7_75t_SL g4754 ( 
.A1(n_4658),
.A2(n_4419),
.B(n_4420),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4678),
.B(n_4388),
.Y(n_4755)
);

NOR2xp67_ASAP7_75t_L g4756 ( 
.A(n_4645),
.B(n_4342),
.Y(n_4756)
);

NAND3xp33_ASAP7_75t_L g4757 ( 
.A(n_4642),
.B(n_4420),
.C(n_4419),
.Y(n_4757)
);

NAND3xp33_ASAP7_75t_L g4758 ( 
.A(n_4642),
.B(n_4388),
.C(n_4357),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4658),
.B(n_4342),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4658),
.B(n_4357),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4682),
.B(n_504),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4619),
.B(n_4644),
.Y(n_4762)
);

AOI221xp5_ASAP7_75t_L g4763 ( 
.A1(n_4701),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.C(n_508),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_L g4764 ( 
.A(n_4644),
.B(n_505),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4605),
.B(n_508),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4696),
.B(n_4607),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4653),
.B(n_509),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4656),
.B(n_510),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4746),
.Y(n_4769)
);

INVx2_ASAP7_75t_SL g4770 ( 
.A(n_4714),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4746),
.Y(n_4771)
);

INVx1_ASAP7_75t_SL g4772 ( 
.A(n_4723),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4714),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4716),
.B(n_4653),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4731),
.B(n_4692),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4749),
.Y(n_4776)
);

NAND2x1p5_ASAP7_75t_L g4777 ( 
.A(n_4756),
.B(n_4645),
.Y(n_4777)
);

OAI22xp5_ASAP7_75t_L g4778 ( 
.A1(n_4709),
.A2(n_4616),
.B1(n_4613),
.B2(n_4674),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4765),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4768),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4732),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_4716),
.B(n_4653),
.Y(n_4782)
);

INVx1_ASAP7_75t_SL g4783 ( 
.A(n_4723),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4762),
.Y(n_4784)
);

AND2x2_ASAP7_75t_L g4785 ( 
.A(n_4713),
.B(n_4696),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4713),
.B(n_4696),
.Y(n_4786)
);

HB1xp67_ASAP7_75t_L g4787 ( 
.A(n_4741),
.Y(n_4787)
);

AOI221xp5_ASAP7_75t_L g4788 ( 
.A1(n_4731),
.A2(n_4694),
.B1(n_4616),
.B2(n_4613),
.C(n_4614),
.Y(n_4788)
);

OR2x2_ASAP7_75t_L g4789 ( 
.A(n_4712),
.B(n_4611),
.Y(n_4789)
);

NOR2xp67_ASAP7_75t_L g4790 ( 
.A(n_4725),
.B(n_4645),
.Y(n_4790)
);

NOR2xp33_ASAP7_75t_L g4791 ( 
.A(n_4707),
.B(n_4626),
.Y(n_4791)
);

OAI22xp33_ASAP7_75t_L g4792 ( 
.A1(n_4718),
.A2(n_4694),
.B1(n_4699),
.B2(n_4646),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4734),
.Y(n_4793)
);

INVx3_ASAP7_75t_L g4794 ( 
.A(n_4766),
.Y(n_4794)
);

AND2x4_ASAP7_75t_L g4795 ( 
.A(n_4724),
.B(n_4645),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4717),
.Y(n_4796)
);

BUFx3_ASAP7_75t_L g4797 ( 
.A(n_4767),
.Y(n_4797)
);

NAND3xp33_ASAP7_75t_L g4798 ( 
.A(n_4727),
.B(n_4656),
.C(n_4612),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4722),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4751),
.Y(n_4800)
);

OR2x2_ASAP7_75t_L g4801 ( 
.A(n_4715),
.B(n_4606),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4752),
.B(n_4689),
.Y(n_4802)
);

AND2x4_ASAP7_75t_L g4803 ( 
.A(n_4766),
.B(n_4639),
.Y(n_4803)
);

AND2x2_ASAP7_75t_L g4804 ( 
.A(n_4719),
.B(n_4672),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4728),
.B(n_4702),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4755),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4721),
.B(n_4733),
.Y(n_4807)
);

OAI22xp5_ASAP7_75t_L g4808 ( 
.A1(n_4744),
.A2(n_4674),
.B1(n_4646),
.B2(n_4703),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4735),
.Y(n_4809)
);

AND2x4_ASAP7_75t_L g4810 ( 
.A(n_4729),
.B(n_4639),
.Y(n_4810)
);

HB1xp67_ASAP7_75t_L g4811 ( 
.A(n_4741),
.Y(n_4811)
);

AND2x2_ASAP7_75t_L g4812 ( 
.A(n_4730),
.B(n_4672),
.Y(n_4812)
);

INVx4_ASAP7_75t_L g4813 ( 
.A(n_4759),
.Y(n_4813)
);

OR2x2_ASAP7_75t_L g4814 ( 
.A(n_4710),
.B(n_4662),
.Y(n_4814)
);

INVx4_ASAP7_75t_L g4815 ( 
.A(n_4760),
.Y(n_4815)
);

BUFx2_ASAP7_75t_L g4816 ( 
.A(n_4742),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4737),
.B(n_4691),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4764),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_4743),
.B(n_4679),
.Y(n_4819)
);

OR2x2_ASAP7_75t_L g4820 ( 
.A(n_4740),
.B(n_4636),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4748),
.Y(n_4821)
);

BUFx2_ASAP7_75t_L g4822 ( 
.A(n_4742),
.Y(n_4822)
);

AOI211xp5_ASAP7_75t_L g4823 ( 
.A1(n_4711),
.A2(n_4685),
.B(n_4609),
.C(n_4622),
.Y(n_4823)
);

AND2x2_ASAP7_75t_L g4824 ( 
.A(n_4743),
.B(n_4679),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4720),
.Y(n_4825)
);

AND2x2_ASAP7_75t_L g4826 ( 
.A(n_4774),
.B(n_4654),
.Y(n_4826)
);

AND2x2_ASAP7_75t_L g4827 ( 
.A(n_4782),
.B(n_4654),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4787),
.Y(n_4828)
);

OR2x2_ASAP7_75t_L g4829 ( 
.A(n_4816),
.B(n_4822),
.Y(n_4829)
);

NOR2xp33_ASAP7_75t_L g4830 ( 
.A(n_4802),
.B(n_4739),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_4777),
.Y(n_4831)
);

NAND5xp2_ASAP7_75t_L g4832 ( 
.A(n_4823),
.B(n_4750),
.C(n_4736),
.D(n_4708),
.E(n_4763),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4787),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4777),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4813),
.B(n_4679),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4804),
.B(n_4654),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_SL g4837 ( 
.A(n_4792),
.B(n_4747),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4811),
.Y(n_4838)
);

OR2x2_ASAP7_75t_L g4839 ( 
.A(n_4805),
.B(n_4745),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4813),
.B(n_4679),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4819),
.B(n_4641),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4811),
.Y(n_4842)
);

NOR2x1_ASAP7_75t_R g4843 ( 
.A(n_4797),
.B(n_4803),
.Y(n_4843)
);

OR2x2_ASAP7_75t_L g4844 ( 
.A(n_4805),
.B(n_4808),
.Y(n_4844)
);

NOR2xp33_ASAP7_75t_L g4845 ( 
.A(n_4802),
.B(n_4693),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4779),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_4824),
.B(n_4693),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4797),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_SL g4849 ( 
.A(n_4790),
.B(n_4693),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4785),
.B(n_4693),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4815),
.B(n_4736),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4815),
.B(n_4664),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4814),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4786),
.B(n_4695),
.Y(n_4854)
);

INVx2_ASAP7_75t_L g4855 ( 
.A(n_4771),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4807),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4771),
.Y(n_4857)
);

AND2x4_ASAP7_75t_L g4858 ( 
.A(n_4795),
.B(n_4609),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4794),
.B(n_4664),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4784),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4789),
.Y(n_4861)
);

AND2x2_ASAP7_75t_L g4862 ( 
.A(n_4812),
.B(n_4670),
.Y(n_4862)
);

AND2x2_ASAP7_75t_L g4863 ( 
.A(n_4795),
.B(n_4817),
.Y(n_4863)
);

AND2x4_ASAP7_75t_L g4864 ( 
.A(n_4803),
.B(n_4660),
.Y(n_4864)
);

OR2x2_ASAP7_75t_L g4865 ( 
.A(n_4808),
.B(n_4738),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4810),
.B(n_4688),
.Y(n_4866)
);

OR2x2_ASAP7_75t_L g4867 ( 
.A(n_4775),
.B(n_4801),
.Y(n_4867)
);

AND2x2_ASAP7_75t_L g4868 ( 
.A(n_4810),
.B(n_4688),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4820),
.Y(n_4869)
);

AND2x2_ASAP7_75t_L g4870 ( 
.A(n_4770),
.B(n_4651),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4828),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4837),
.B(n_4788),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4836),
.Y(n_4873)
);

OR2x2_ASAP7_75t_L g4874 ( 
.A(n_4829),
.B(n_4775),
.Y(n_4874)
);

OR2x2_ASAP7_75t_L g4875 ( 
.A(n_4867),
.B(n_4825),
.Y(n_4875)
);

INVxp67_ASAP7_75t_SL g4876 ( 
.A(n_4843),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4833),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4836),
.B(n_4794),
.Y(n_4878)
);

NAND2xp67_ASAP7_75t_L g4879 ( 
.A(n_4841),
.B(n_4825),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_4870),
.B(n_4845),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4837),
.B(n_4788),
.Y(n_4881)
);

NAND2x1p5_ASAP7_75t_L g4882 ( 
.A(n_4831),
.B(n_4772),
.Y(n_4882)
);

NOR2xp33_ASAP7_75t_L g4883 ( 
.A(n_4849),
.B(n_4791),
.Y(n_4883)
);

NOR2xp33_ASAP7_75t_L g4884 ( 
.A(n_4841),
.B(n_4791),
.Y(n_4884)
);

NOR2x1_ASAP7_75t_L g4885 ( 
.A(n_4844),
.B(n_4772),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4830),
.B(n_4792),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4838),
.Y(n_4887)
);

AND2x2_ASAP7_75t_L g4888 ( 
.A(n_4847),
.B(n_4773),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4870),
.B(n_4778),
.Y(n_4889)
);

INVx2_ASAP7_75t_L g4890 ( 
.A(n_4842),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_4859),
.Y(n_4891)
);

NOR2xp33_ASAP7_75t_L g4892 ( 
.A(n_4847),
.B(n_4781),
.Y(n_4892)
);

OAI21xp33_ASAP7_75t_L g4893 ( 
.A1(n_4830),
.A2(n_4778),
.B(n_4726),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4826),
.B(n_4793),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4845),
.B(n_4769),
.Y(n_4895)
);

INVxp67_ASAP7_75t_SL g4896 ( 
.A(n_4826),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4827),
.B(n_4809),
.Y(n_4897)
);

OR2x2_ASAP7_75t_L g4898 ( 
.A(n_4856),
.B(n_4798),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4848),
.B(n_4783),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4827),
.B(n_4796),
.Y(n_4900)
);

HB1xp67_ASAP7_75t_L g4901 ( 
.A(n_4858),
.Y(n_4901)
);

OAI332xp33_ASAP7_75t_L g4902 ( 
.A1(n_4872),
.A2(n_4783),
.A3(n_4865),
.B1(n_4839),
.B2(n_4821),
.B3(n_4855),
.C1(n_4857),
.C2(n_4851),
.Y(n_4902)
);

HB1xp67_ASAP7_75t_L g4903 ( 
.A(n_4901),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4896),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4882),
.Y(n_4905)
);

OR2x2_ASAP7_75t_L g4906 ( 
.A(n_4889),
.B(n_4852),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4872),
.B(n_4855),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4873),
.Y(n_4908)
);

HB1xp67_ASAP7_75t_L g4909 ( 
.A(n_4882),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4881),
.B(n_4857),
.Y(n_4910)
);

OAI31xp33_ASAP7_75t_L g4911 ( 
.A1(n_4881),
.A2(n_4832),
.A3(n_4864),
.B(n_4858),
.Y(n_4911)
);

HB1xp67_ASAP7_75t_L g4912 ( 
.A(n_4879),
.Y(n_4912)
);

INVx2_ASAP7_75t_SL g4913 ( 
.A(n_4888),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4899),
.Y(n_4914)
);

OAI322xp33_ASAP7_75t_L g4915 ( 
.A1(n_4886),
.A2(n_4898),
.A3(n_4875),
.B1(n_4874),
.B2(n_4895),
.C1(n_4899),
.C2(n_4880),
.Y(n_4915)
);

OAI31xp67_ASAP7_75t_L g4916 ( 
.A1(n_4890),
.A2(n_4831),
.A3(n_4834),
.B(n_4754),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4876),
.B(n_4866),
.Y(n_4917)
);

INVxp67_ASAP7_75t_SL g4918 ( 
.A(n_4885),
.Y(n_4918)
);

INVx1_ASAP7_75t_SL g4919 ( 
.A(n_4886),
.Y(n_4919)
);

NOR2x1p5_ASAP7_75t_L g4920 ( 
.A(n_4878),
.B(n_4835),
.Y(n_4920)
);

OR2x2_ASAP7_75t_L g4921 ( 
.A(n_4891),
.B(n_4861),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4900),
.Y(n_4922)
);

INVx2_ASAP7_75t_L g4923 ( 
.A(n_4894),
.Y(n_4923)
);

AOI22xp5_ASAP7_75t_L g4924 ( 
.A1(n_4893),
.A2(n_4850),
.B1(n_4863),
.B2(n_4862),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4903),
.Y(n_4925)
);

XOR2x2_ASAP7_75t_L g4926 ( 
.A(n_4924),
.B(n_4884),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4909),
.Y(n_4927)
);

INVxp67_ASAP7_75t_SL g4928 ( 
.A(n_4912),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4913),
.B(n_4866),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4918),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4917),
.Y(n_4931)
);

XOR2x2_ASAP7_75t_L g4932 ( 
.A(n_4906),
.B(n_4883),
.Y(n_4932)
);

BUFx12f_ASAP7_75t_L g4933 ( 
.A(n_4920),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4904),
.Y(n_4934)
);

XOR2xp5_ASAP7_75t_L g4935 ( 
.A(n_4922),
.B(n_4850),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4923),
.Y(n_4936)
);

XNOR2x2_ASAP7_75t_L g4937 ( 
.A(n_4919),
.B(n_4892),
.Y(n_4937)
);

INVx2_ASAP7_75t_L g4938 ( 
.A(n_4905),
.Y(n_4938)
);

NOR2xp33_ASAP7_75t_SL g4939 ( 
.A(n_4915),
.B(n_4897),
.Y(n_4939)
);

OA22x2_ASAP7_75t_L g4940 ( 
.A1(n_4919),
.A2(n_4858),
.B1(n_4834),
.B2(n_4840),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4908),
.Y(n_4941)
);

AO22x1_ASAP7_75t_L g4942 ( 
.A1(n_4907),
.A2(n_4910),
.B1(n_4864),
.B2(n_4877),
.Y(n_4942)
);

INVxp67_ASAP7_75t_L g4943 ( 
.A(n_4907),
.Y(n_4943)
);

XOR2x2_ASAP7_75t_L g4944 ( 
.A(n_4910),
.B(n_4854),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4942),
.Y(n_4945)
);

AND2x2_ASAP7_75t_L g4946 ( 
.A(n_4938),
.B(n_4868),
.Y(n_4946)
);

AND2x2_ASAP7_75t_L g4947 ( 
.A(n_4927),
.B(n_4868),
.Y(n_4947)
);

INVx1_ASAP7_75t_SL g4948 ( 
.A(n_4937),
.Y(n_4948)
);

BUFx2_ASAP7_75t_L g4949 ( 
.A(n_4933),
.Y(n_4949)
);

OR2x2_ASAP7_75t_L g4950 ( 
.A(n_4929),
.B(n_4853),
.Y(n_4950)
);

AND2x2_ASAP7_75t_L g4951 ( 
.A(n_4936),
.B(n_4869),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4928),
.B(n_4911),
.Y(n_4952)
);

OR2x2_ASAP7_75t_L g4953 ( 
.A(n_4925),
.B(n_4860),
.Y(n_4953)
);

HB1xp67_ASAP7_75t_L g4954 ( 
.A(n_4940),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4935),
.Y(n_4955)
);

CKINVDCx16_ASAP7_75t_R g4956 ( 
.A(n_4939),
.Y(n_4956)
);

INVx3_ASAP7_75t_L g4957 ( 
.A(n_4925),
.Y(n_4957)
);

OR2x2_ASAP7_75t_L g4958 ( 
.A(n_4930),
.B(n_4846),
.Y(n_4958)
);

INVxp67_ASAP7_75t_SL g4959 ( 
.A(n_4957),
.Y(n_4959)
);

AOI31xp33_ASAP7_75t_L g4960 ( 
.A1(n_4948),
.A2(n_4943),
.A3(n_4921),
.B(n_4914),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4947),
.Y(n_4961)
);

AOI21xp5_ASAP7_75t_L g4962 ( 
.A1(n_4945),
.A2(n_4902),
.B(n_4942),
.Y(n_4962)
);

AOI22xp33_ASAP7_75t_L g4963 ( 
.A1(n_4949),
.A2(n_4660),
.B1(n_4864),
.B2(n_4931),
.Y(n_4963)
);

AO22x1_ASAP7_75t_L g4964 ( 
.A1(n_4945),
.A2(n_4887),
.B1(n_4871),
.B2(n_4934),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4946),
.B(n_4951),
.Y(n_4965)
);

AOI22xp5_ASAP7_75t_L g4966 ( 
.A1(n_4956),
.A2(n_4675),
.B1(n_4944),
.B2(n_4926),
.Y(n_4966)
);

AOI211xp5_ASAP7_75t_L g4967 ( 
.A1(n_4954),
.A2(n_4941),
.B(n_4799),
.C(n_4776),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4959),
.B(n_4957),
.Y(n_4968)
);

OAI22xp33_ASAP7_75t_L g4969 ( 
.A1(n_4960),
.A2(n_4675),
.B1(n_4952),
.B2(n_4950),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_L g4970 ( 
.A(n_4964),
.B(n_4818),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4965),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_L g4972 ( 
.A(n_4962),
.B(n_4955),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4961),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4966),
.Y(n_4974)
);

AOI22xp5_ASAP7_75t_L g4975 ( 
.A1(n_4967),
.A2(n_4675),
.B1(n_4932),
.B2(n_4780),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4963),
.Y(n_4976)
);

AND2x4_ASAP7_75t_L g4977 ( 
.A(n_4965),
.B(n_4953),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4959),
.Y(n_4978)
);

AOI221xp5_ASAP7_75t_L g4979 ( 
.A1(n_4962),
.A2(n_4800),
.B1(n_4806),
.B2(n_4958),
.C(n_4629),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4959),
.B(n_4621),
.Y(n_4980)
);

AOI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4966),
.A2(n_4675),
.B1(n_4633),
.B2(n_4635),
.Y(n_4981)
);

NOR2x1_ASAP7_75t_L g4982 ( 
.A(n_4968),
.B(n_4761),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4977),
.B(n_4637),
.Y(n_4983)
);

INVx1_ASAP7_75t_SL g4984 ( 
.A(n_4970),
.Y(n_4984)
);

INVx3_ASAP7_75t_SL g4985 ( 
.A(n_4971),
.Y(n_4985)
);

NOR2xp33_ASAP7_75t_L g4986 ( 
.A(n_4978),
.B(n_4916),
.Y(n_4986)
);

NAND2x1_ASAP7_75t_SL g4987 ( 
.A(n_4975),
.B(n_4618),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4973),
.B(n_4648),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4981),
.B(n_4753),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4969),
.B(n_4655),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4979),
.B(n_4659),
.Y(n_4991)
);

NOR2x1_ASAP7_75t_L g4992 ( 
.A(n_4980),
.B(n_4638),
.Y(n_4992)
);

AND2x2_ASAP7_75t_L g4993 ( 
.A(n_4974),
.B(n_4651),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4972),
.Y(n_4994)
);

AND2x2_ASAP7_75t_L g4995 ( 
.A(n_4976),
.B(n_4652),
.Y(n_4995)
);

INVx2_ASAP7_75t_SL g4996 ( 
.A(n_4977),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4977),
.B(n_4673),
.Y(n_4997)
);

OR2x2_ASAP7_75t_L g4998 ( 
.A(n_4968),
.B(n_4647),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4968),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4977),
.B(n_4652),
.Y(n_5000)
);

NOR2xp33_ASAP7_75t_L g5001 ( 
.A(n_4971),
.B(n_4686),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4977),
.B(n_4684),
.Y(n_5002)
);

NOR2xp33_ASAP7_75t_L g5003 ( 
.A(n_4971),
.B(n_4618),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4977),
.B(n_4684),
.Y(n_5004)
);

AOI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_4996),
.A2(n_4618),
.B1(n_4640),
.B2(n_4747),
.Y(n_5005)
);

AND4x1_ASAP7_75t_L g5006 ( 
.A(n_4986),
.B(n_4757),
.C(n_4758),
.D(n_4706),
.Y(n_5006)
);

AOI22xp5_ASAP7_75t_L g5007 ( 
.A1(n_5003),
.A2(n_5004),
.B1(n_5002),
.B2(n_4993),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_5000),
.Y(n_5008)
);

OA22x2_ASAP7_75t_L g5009 ( 
.A1(n_4985),
.A2(n_4638),
.B1(n_4640),
.B2(n_4603),
.Y(n_5009)
);

INVx2_ASAP7_75t_L g5010 ( 
.A(n_4998),
.Y(n_5010)
);

HB1xp67_ASAP7_75t_L g5011 ( 
.A(n_4992),
.Y(n_5011)
);

OAI22xp5_ASAP7_75t_L g5012 ( 
.A1(n_4984),
.A2(n_4698),
.B1(n_4640),
.B2(n_4603),
.Y(n_5012)
);

INVx3_ASAP7_75t_L g5013 ( 
.A(n_4995),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4989),
.Y(n_5014)
);

INVx1_ASAP7_75t_SL g5015 ( 
.A(n_4987),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4983),
.Y(n_5016)
);

OAI22xp5_ASAP7_75t_L g5017 ( 
.A1(n_4994),
.A2(n_4603),
.B1(n_4657),
.B2(n_4706),
.Y(n_5017)
);

AOI22xp5_ASAP7_75t_L g5018 ( 
.A1(n_4999),
.A2(n_4657),
.B1(n_4667),
.B2(n_4632),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4997),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4982),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_5001),
.Y(n_5021)
);

INVx2_ASAP7_75t_L g5022 ( 
.A(n_4999),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4988),
.Y(n_5023)
);

AOI221xp5_ASAP7_75t_L g5024 ( 
.A1(n_4991),
.A2(n_4690),
.B1(n_511),
.B2(n_512),
.C(n_513),
.Y(n_5024)
);

NAND4xp25_ASAP7_75t_L g5025 ( 
.A(n_4990),
.B(n_510),
.C(n_511),
.D(n_512),
.Y(n_5025)
);

OAI22x1_ASAP7_75t_L g5026 ( 
.A1(n_4985),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_5026)
);

NAND4xp25_ASAP7_75t_L g5027 ( 
.A(n_4986),
.B(n_516),
.C(n_517),
.D(n_518),
.Y(n_5027)
);

AOI22xp5_ASAP7_75t_L g5028 ( 
.A1(n_4996),
.A2(n_516),
.B1(n_517),
.B2(n_520),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_5002),
.Y(n_5029)
);

OAI222xp33_ASAP7_75t_L g5030 ( 
.A1(n_4996),
.A2(n_671),
.B1(n_521),
.B2(n_522),
.C1(n_523),
.C2(n_525),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_5005),
.B(n_520),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_5018),
.B(n_521),
.Y(n_5032)
);

NOR3x1_ASAP7_75t_L g5033 ( 
.A(n_5025),
.B(n_5027),
.C(n_5008),
.Y(n_5033)
);

AOI22xp5_ASAP7_75t_L g5034 ( 
.A1(n_5017),
.A2(n_522),
.B1(n_523),
.B2(n_526),
.Y(n_5034)
);

AOI21xp5_ASAP7_75t_L g5035 ( 
.A1(n_5015),
.A2(n_526),
.B(n_527),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_5009),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_5011),
.Y(n_5037)
);

NOR3xp33_ASAP7_75t_L g5038 ( 
.A(n_5014),
.B(n_528),
.C(n_529),
.Y(n_5038)
);

HB1xp67_ASAP7_75t_L g5039 ( 
.A(n_5026),
.Y(n_5039)
);

AO22x2_ASAP7_75t_L g5040 ( 
.A1(n_5029),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_5040)
);

OAI211xp5_ASAP7_75t_SL g5041 ( 
.A1(n_5007),
.A2(n_5013),
.B(n_5020),
.C(n_5021),
.Y(n_5041)
);

NOR2x1_ASAP7_75t_L g5042 ( 
.A(n_5030),
.B(n_531),
.Y(n_5042)
);

AOI211xp5_ASAP7_75t_L g5043 ( 
.A1(n_5012),
.A2(n_531),
.B(n_532),
.C(n_533),
.Y(n_5043)
);

AOI22xp5_ASAP7_75t_L g5044 ( 
.A1(n_5010),
.A2(n_533),
.B1(n_534),
.B2(n_535),
.Y(n_5044)
);

AOI22xp5_ASAP7_75t_SL g5045 ( 
.A1(n_5013),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.Y(n_5045)
);

AOI22xp5_ASAP7_75t_L g5046 ( 
.A1(n_5022),
.A2(n_537),
.B1(n_538),
.B2(n_540),
.Y(n_5046)
);

NOR3xp33_ASAP7_75t_L g5047 ( 
.A(n_5016),
.B(n_537),
.C(n_538),
.Y(n_5047)
);

AOI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_5019),
.A2(n_540),
.B(n_541),
.Y(n_5048)
);

AOI211xp5_ASAP7_75t_L g5049 ( 
.A1(n_5024),
.A2(n_5023),
.B(n_5028),
.C(n_5006),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_5005),
.B(n_542),
.Y(n_5050)
);

OAI22xp5_ASAP7_75t_L g5051 ( 
.A1(n_5005),
.A2(n_542),
.B1(n_543),
.B2(n_544),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_5005),
.B(n_543),
.Y(n_5052)
);

OA22x2_ASAP7_75t_L g5053 ( 
.A1(n_5005),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_5009),
.Y(n_5054)
);

XNOR2x1_ASAP7_75t_SL g5055 ( 
.A(n_5036),
.B(n_545),
.Y(n_5055)
);

NOR3xp33_ASAP7_75t_L g5056 ( 
.A(n_5041),
.B(n_546),
.C(n_548),
.Y(n_5056)
);

NOR4xp25_ASAP7_75t_L g5057 ( 
.A(n_5031),
.B(n_549),
.C(n_550),
.D(n_551),
.Y(n_5057)
);

NOR4xp25_ASAP7_75t_L g5058 ( 
.A(n_5050),
.B(n_551),
.C(n_552),
.D(n_553),
.Y(n_5058)
);

NOR4xp75_ASAP7_75t_L g5059 ( 
.A(n_5052),
.B(n_553),
.C(n_554),
.D(n_555),
.Y(n_5059)
);

NOR2xp33_ASAP7_75t_L g5060 ( 
.A(n_5039),
.B(n_554),
.Y(n_5060)
);

NOR2x1_ASAP7_75t_L g5061 ( 
.A(n_5054),
.B(n_555),
.Y(n_5061)
);

OAI22xp33_ASAP7_75t_L g5062 ( 
.A1(n_5034),
.A2(n_556),
.B1(n_557),
.B2(n_558),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_5038),
.B(n_556),
.Y(n_5063)
);

AOI22xp5_ASAP7_75t_L g5064 ( 
.A1(n_5037),
.A2(n_557),
.B1(n_558),
.B2(n_560),
.Y(n_5064)
);

NAND3xp33_ASAP7_75t_SL g5065 ( 
.A(n_5043),
.B(n_5035),
.C(n_5049),
.Y(n_5065)
);

NOR2xp67_ASAP7_75t_L g5066 ( 
.A(n_5048),
.B(n_560),
.Y(n_5066)
);

NOR2x1p5_ASAP7_75t_L g5067 ( 
.A(n_5032),
.B(n_561),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_5053),
.Y(n_5068)
);

AOI211x1_ASAP7_75t_L g5069 ( 
.A1(n_5051),
.A2(n_561),
.B(n_562),
.C(n_563),
.Y(n_5069)
);

NAND3xp33_ASAP7_75t_L g5070 ( 
.A(n_5047),
.B(n_562),
.C(n_564),
.Y(n_5070)
);

NOR3xp33_ASAP7_75t_L g5071 ( 
.A(n_5042),
.B(n_565),
.C(n_566),
.Y(n_5071)
);

OAI211xp5_ASAP7_75t_SL g5072 ( 
.A1(n_5068),
.A2(n_5033),
.B(n_5044),
.C(n_5046),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_5060),
.Y(n_5073)
);

NOR3xp33_ASAP7_75t_L g5074 ( 
.A(n_5065),
.B(n_5045),
.C(n_5040),
.Y(n_5074)
);

NAND4xp75_ASAP7_75t_L g5075 ( 
.A(n_5061),
.B(n_565),
.C(n_567),
.D(n_568),
.Y(n_5075)
);

NOR3xp33_ASAP7_75t_L g5076 ( 
.A(n_5056),
.B(n_567),
.C(n_568),
.Y(n_5076)
);

AND2x2_ASAP7_75t_SL g5077 ( 
.A(n_5071),
.B(n_569),
.Y(n_5077)
);

AOI22xp5_ASAP7_75t_L g5078 ( 
.A1(n_5067),
.A2(n_670),
.B1(n_571),
.B2(n_573),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_5055),
.B(n_570),
.Y(n_5079)
);

NOR2x1p5_ASAP7_75t_L g5080 ( 
.A(n_5063),
.B(n_574),
.Y(n_5080)
);

OR2x2_ASAP7_75t_L g5081 ( 
.A(n_5057),
.B(n_575),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_5058),
.B(n_575),
.Y(n_5082)
);

AND3x1_ASAP7_75t_L g5083 ( 
.A(n_5064),
.B(n_576),
.C(n_577),
.Y(n_5083)
);

NAND4xp25_ASAP7_75t_L g5084 ( 
.A(n_5069),
.B(n_576),
.C(n_577),
.D(n_578),
.Y(n_5084)
);

NOR4xp25_ASAP7_75t_L g5085 ( 
.A(n_5070),
.B(n_579),
.C(n_580),
.D(n_581),
.Y(n_5085)
);

INVx2_ASAP7_75t_L g5086 ( 
.A(n_5059),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_5079),
.Y(n_5087)
);

AOI21xp33_ASAP7_75t_L g5088 ( 
.A1(n_5081),
.A2(n_5082),
.B(n_5077),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_5078),
.B(n_5066),
.Y(n_5089)
);

INVxp33_ASAP7_75t_SL g5090 ( 
.A(n_5074),
.Y(n_5090)
);

AOI221x1_ASAP7_75t_L g5091 ( 
.A1(n_5072),
.A2(n_5062),
.B1(n_584),
.B2(n_586),
.C(n_587),
.Y(n_5091)
);

AOI22xp5_ASAP7_75t_L g5092 ( 
.A1(n_5076),
.A2(n_583),
.B1(n_584),
.B2(n_587),
.Y(n_5092)
);

AOI211xp5_ASAP7_75t_L g5093 ( 
.A1(n_5085),
.A2(n_588),
.B(n_590),
.C(n_591),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_5075),
.Y(n_5094)
);

OAI21xp33_ASAP7_75t_L g5095 ( 
.A1(n_5086),
.A2(n_588),
.B(n_591),
.Y(n_5095)
);

AOI221xp5_ASAP7_75t_L g5096 ( 
.A1(n_5083),
.A2(n_592),
.B1(n_593),
.B2(n_594),
.C(n_595),
.Y(n_5096)
);

OAI22xp5_ASAP7_75t_L g5097 ( 
.A1(n_5073),
.A2(n_593),
.B1(n_596),
.B2(n_598),
.Y(n_5097)
);

OAI211xp5_ASAP7_75t_L g5098 ( 
.A1(n_5084),
.A2(n_596),
.B(n_599),
.C(n_601),
.Y(n_5098)
);

OAI221xp5_ASAP7_75t_L g5099 ( 
.A1(n_5080),
.A2(n_602),
.B1(n_603),
.B2(n_604),
.C(n_605),
.Y(n_5099)
);

INVx2_ASAP7_75t_SL g5100 ( 
.A(n_5079),
.Y(n_5100)
);

HB1xp67_ASAP7_75t_L g5101 ( 
.A(n_5079),
.Y(n_5101)
);

HB1xp67_ASAP7_75t_L g5102 ( 
.A(n_5079),
.Y(n_5102)
);

OAI21xp5_ASAP7_75t_L g5103 ( 
.A1(n_5079),
.A2(n_602),
.B(n_604),
.Y(n_5103)
);

OAI21xp33_ASAP7_75t_SL g5104 ( 
.A1(n_5079),
.A2(n_605),
.B(n_606),
.Y(n_5104)
);

NOR2x1_ASAP7_75t_L g5105 ( 
.A(n_5103),
.B(n_606),
.Y(n_5105)
);

INVx2_ASAP7_75t_L g5106 ( 
.A(n_5100),
.Y(n_5106)
);

OAI211xp5_ASAP7_75t_SL g5107 ( 
.A1(n_5088),
.A2(n_607),
.B(n_608),
.C(n_609),
.Y(n_5107)
);

AOI22xp5_ASAP7_75t_L g5108 ( 
.A1(n_5090),
.A2(n_5094),
.B1(n_5098),
.B2(n_5087),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_5101),
.Y(n_5109)
);

AOI22xp5_ASAP7_75t_L g5110 ( 
.A1(n_5096),
.A2(n_607),
.B1(n_610),
.B2(n_611),
.Y(n_5110)
);

AOI22xp5_ASAP7_75t_L g5111 ( 
.A1(n_5102),
.A2(n_610),
.B1(n_611),
.B2(n_612),
.Y(n_5111)
);

INVx2_ASAP7_75t_L g5112 ( 
.A(n_5099),
.Y(n_5112)
);

INVxp67_ASAP7_75t_L g5113 ( 
.A(n_5095),
.Y(n_5113)
);

AOI22xp5_ASAP7_75t_L g5114 ( 
.A1(n_5104),
.A2(n_612),
.B1(n_613),
.B2(n_614),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_5091),
.Y(n_5115)
);

AOI22xp33_ASAP7_75t_SL g5116 ( 
.A1(n_5089),
.A2(n_613),
.B1(n_614),
.B2(n_615),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_5097),
.Y(n_5117)
);

NOR2x1_ASAP7_75t_L g5118 ( 
.A(n_5093),
.B(n_616),
.Y(n_5118)
);

INVx2_ASAP7_75t_L g5119 ( 
.A(n_5092),
.Y(n_5119)
);

INVx2_ASAP7_75t_L g5120 ( 
.A(n_5100),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_SL g5121 ( 
.A(n_5096),
.B(n_616),
.Y(n_5121)
);

OR2x2_ASAP7_75t_L g5122 ( 
.A(n_5115),
.B(n_5114),
.Y(n_5122)
);

NAND4xp25_ASAP7_75t_L g5123 ( 
.A(n_5108),
.B(n_618),
.C(n_619),
.D(n_620),
.Y(n_5123)
);

NOR3xp33_ASAP7_75t_L g5124 ( 
.A(n_5109),
.B(n_618),
.C(n_619),
.Y(n_5124)
);

NAND4xp75_ASAP7_75t_L g5125 ( 
.A(n_5105),
.B(n_620),
.C(n_621),
.D(n_622),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_5118),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5110),
.Y(n_5127)
);

NOR3xp33_ASAP7_75t_L g5128 ( 
.A(n_5106),
.B(n_5120),
.C(n_5113),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_5121),
.A2(n_622),
.B(n_623),
.Y(n_5129)
);

NOR3xp33_ASAP7_75t_L g5130 ( 
.A(n_5117),
.B(n_623),
.C(n_624),
.Y(n_5130)
);

AOI22xp5_ASAP7_75t_L g5131 ( 
.A1(n_5107),
.A2(n_624),
.B1(n_626),
.B2(n_627),
.Y(n_5131)
);

OR2x2_ASAP7_75t_L g5132 ( 
.A(n_5119),
.B(n_626),
.Y(n_5132)
);

AND2x4_ASAP7_75t_L g5133 ( 
.A(n_5128),
.B(n_5112),
.Y(n_5133)
);

NAND4xp75_ASAP7_75t_L g5134 ( 
.A(n_5126),
.B(n_5111),
.C(n_5116),
.D(n_630),
.Y(n_5134)
);

NOR3xp33_ASAP7_75t_L g5135 ( 
.A(n_5122),
.B(n_628),
.C(n_629),
.Y(n_5135)
);

OAI21xp33_ASAP7_75t_SL g5136 ( 
.A1(n_5131),
.A2(n_628),
.B(n_629),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_5125),
.Y(n_5137)
);

NOR3xp33_ASAP7_75t_L g5138 ( 
.A(n_5127),
.B(n_630),
.C(n_631),
.Y(n_5138)
);

INVx3_ASAP7_75t_L g5139 ( 
.A(n_5133),
.Y(n_5139)
);

INVxp67_ASAP7_75t_L g5140 ( 
.A(n_5137),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5134),
.Y(n_5141)
);

AO21x1_ASAP7_75t_L g5142 ( 
.A1(n_5141),
.A2(n_5129),
.B(n_5130),
.Y(n_5142)
);

OAI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_5140),
.A2(n_5136),
.B(n_5123),
.Y(n_5143)
);

AO22x2_ASAP7_75t_L g5144 ( 
.A1(n_5143),
.A2(n_5139),
.B1(n_5135),
.B2(n_5124),
.Y(n_5144)
);

OAI221xp5_ASAP7_75t_SL g5145 ( 
.A1(n_5144),
.A2(n_5138),
.B1(n_5132),
.B2(n_5142),
.C(n_635),
.Y(n_5145)
);

INVxp67_ASAP7_75t_SL g5146 ( 
.A(n_5145),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_5146),
.B(n_632),
.Y(n_5147)
);

BUFx3_ASAP7_75t_L g5148 ( 
.A(n_5147),
.Y(n_5148)
);

AO22x2_ASAP7_75t_L g5149 ( 
.A1(n_5148),
.A2(n_633),
.B1(n_634),
.B2(n_636),
.Y(n_5149)
);

AOI21xp5_ASAP7_75t_L g5150 ( 
.A1(n_5149),
.A2(n_636),
.B(n_637),
.Y(n_5150)
);

AOI21xp5_ASAP7_75t_L g5151 ( 
.A1(n_5150),
.A2(n_637),
.B(n_638),
.Y(n_5151)
);

AOI22xp5_ASAP7_75t_L g5152 ( 
.A1(n_5151),
.A2(n_638),
.B1(n_639),
.B2(n_640),
.Y(n_5152)
);

OR2x6_ASAP7_75t_L g5153 ( 
.A(n_5152),
.B(n_639),
.Y(n_5153)
);

AOI221xp5_ASAP7_75t_L g5154 ( 
.A1(n_5153),
.A2(n_641),
.B1(n_643),
.B2(n_644),
.C(n_645),
.Y(n_5154)
);

OAI221xp5_ASAP7_75t_R g5155 ( 
.A1(n_5153),
.A2(n_644),
.B1(n_645),
.B2(n_646),
.C(n_647),
.Y(n_5155)
);

AOI22xp5_ASAP7_75t_L g5156 ( 
.A1(n_5155),
.A2(n_5154),
.B1(n_647),
.B2(n_649),
.Y(n_5156)
);

AOI211xp5_ASAP7_75t_L g5157 ( 
.A1(n_5156),
.A2(n_670),
.B(n_650),
.C(n_651),
.Y(n_5157)
);


endmodule