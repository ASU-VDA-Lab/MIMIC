module fake_ariane_349_n_289 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_54, n_25, n_289);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_54;
input n_25;

output n_289;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_288;
wire n_179;
wire n_64;
wire n_180;
wire n_160;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_110;
wire n_153;
wire n_197;
wire n_221;
wire n_86;
wire n_269;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_259;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_111;
wire n_242;
wire n_260;
wire n_274;
wire n_115;
wire n_272;
wire n_133;
wire n_66;
wire n_205;
wire n_236;
wire n_265;
wire n_71;
wire n_267;
wire n_208;
wire n_109;
wire n_245;
wire n_96;
wire n_156;
wire n_281;
wire n_209;
wire n_262;
wire n_286;
wire n_174;
wire n_275;
wire n_100;
wire n_283;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_235;
wire n_225;
wire n_200;
wire n_166;
wire n_253;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_246;
wire n_244;
wire n_226;
wire n_271;
wire n_220;
wire n_84;
wire n_247;
wire n_261;
wire n_199;
wire n_91;
wire n_189;
wire n_107;
wire n_159;
wire n_72;
wire n_105;
wire n_128;
wire n_217;
wire n_224;
wire n_240;
wire n_82;
wire n_178;
wire n_57;
wire n_131;
wire n_263;
wire n_201;
wire n_229;
wire n_70;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_287;
wire n_85;
wire n_130;
wire n_144;
wire n_256;
wire n_214;
wire n_227;
wire n_94;
wire n_101;
wire n_243;
wire n_284;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_162;
wire n_264;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_278;
wire n_122;
wire n_268;
wire n_257;
wire n_266;
wire n_198;
wire n_282;
wire n_148;
wire n_232;
wire n_164;
wire n_277;
wire n_157;
wire n_248;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_118;
wire n_93;
wire n_121;
wire n_276;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_87;
wire n_81;
wire n_206;
wire n_279;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_219;
wire n_140;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_270;
wire n_194;
wire n_97;
wire n_154;
wire n_280;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_285;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_63;
wire n_59;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_273;

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVxp33_ASAP7_75t_SL g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_29),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVxp33_ASAP7_75t_SL g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_5),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_0),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_0),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_1),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_1),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_2),
.Y(n_97)
);

AOI22x1_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_6),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_8),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_9),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NAND2x1_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_81),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_81),
.B1(n_80),
.B2(n_67),
.C(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_97),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_83),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_109),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_62),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_68),
.B1(n_70),
.B2(n_85),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_14),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_92),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_110),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_108),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_102),
.B1(n_91),
.B2(n_88),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_127),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

OR2x6_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_102),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_118),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_119),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_135),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_91),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_131),
.B1(n_111),
.B2(n_121),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_88),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_128),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_128),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_100),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_128),
.B(n_98),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_111),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_142),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2x1_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_141),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_144),
.B1(n_137),
.B2(n_146),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

AO31x2_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_141),
.A3(n_139),
.B(n_146),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_165),
.B(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_189),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_152),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_152),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

OAI221xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_150),
.B1(n_162),
.B2(n_159),
.C(n_166),
.Y(n_203)
);

AND2x4_ASAP7_75t_SL g204 ( 
.A(n_177),
.B(n_156),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_183),
.B1(n_196),
.B2(n_150),
.Y(n_211)
);

AO21x2_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_190),
.B(n_171),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_164),
.B1(n_172),
.B2(n_160),
.Y(n_214)
);

OAI211xp5_ASAP7_75t_SL g215 ( 
.A1(n_194),
.A2(n_167),
.B(n_174),
.C(n_160),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_174),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_195),
.B1(n_208),
.B2(n_199),
.Y(n_221)
);

OAI31xp33_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_201),
.A3(n_200),
.B(n_172),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

OAI33xp33_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_167),
.A3(n_187),
.B1(n_170),
.B2(n_156),
.B3(n_139),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_204),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_210),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_192),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_156),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_156),
.Y(n_230)
);

NOR2x1p5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_181),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_187),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_139),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_211),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_218),
.Y(n_242)
);

NOR2x1p5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_215),
.C(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_214),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_237),
.B(n_17),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_212),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_212),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_212),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_16),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_21),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_24),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_242),
.B(n_250),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_244),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_252),
.B(n_251),
.C(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_263),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

NOR4xp25_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_257),
.C(n_261),
.D(n_256),
.Y(n_276)
);

AOI211xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_257),
.B(n_255),
.C(n_254),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_259),
.C(n_254),
.Y(n_278)
);

AOI221xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_259),
.B1(n_139),
.B2(n_31),
.C(n_33),
.Y(n_279)
);

NOR2x1p5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_139),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_25),
.B(n_26),
.Y(n_281)
);

OR3x1_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_36),
.C(n_40),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_282),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_47),
.Y(n_286)
);

AOI311xp33_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_50),
.A3(n_51),
.B(n_52),
.C(n_53),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

AOI221xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_281),
.B1(n_285),
.B2(n_284),
.C(n_287),
.Y(n_289)
);


endmodule