module fake_jpeg_16753_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_5),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_22),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_1),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_21),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_2),
.B1(n_13),
.B2(n_10),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_7),
.B1(n_12),
.B2(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_8),
.B(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_12),
.B1(n_14),
.B2(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_12),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_26),
.B(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

OAI221xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_35),
.B2(n_33),
.C(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_40),
.C(n_38),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_42),
.Y(n_44)
);


endmodule