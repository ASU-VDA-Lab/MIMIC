module real_jpeg_28130_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_292;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_295;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

INVx11_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_0),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_55),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_4),
.A2(n_36),
.B1(n_45),
.B2(n_48),
.Y(n_184)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_6),
.A2(n_74),
.B1(n_75),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_6),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_122),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_122),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_6),
.A2(n_45),
.B1(n_48),
.B2(n_122),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_38),
.B1(n_45),
.B2(n_48),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_74),
.B1(n_75),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_170),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_170),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_8),
.A2(n_45),
.B1(n_48),
.B2(n_170),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_42),
.B1(n_74),
.B2(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_145)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_74),
.B1(n_75),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_11),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_149),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_149),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_11),
.A2(n_45),
.B1(n_48),
.B2(n_149),
.Y(n_250)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_13),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_14),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_70),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_27),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_14),
.A2(n_27),
.B(n_210),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_168),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_14),
.A2(n_45),
.B(n_49),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_14),
.B(n_116),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_14),
.A2(n_86),
.B1(n_141),
.B2(n_258),
.Y(n_260)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_99),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_19),
.B(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_83),
.B2(n_84),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_56),
.B2(n_57),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_23),
.A2(n_24),
.B(n_39),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_25),
.B(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_25),
.A2(n_31),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_31),
.B1(n_164),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_25),
.A2(n_31),
.B1(n_193),
.B2(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_28),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_27),
.B(n_71),
.Y(n_182)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_28),
.A2(n_78),
.B1(n_167),
.B2(n_182),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_28),
.A2(n_32),
.A3(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_31),
.B(n_145),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_33),
.B1(n_47),
.B2(n_49),
.Y(n_53)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_33),
.B(n_208),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_33),
.A2(n_47),
.B(n_168),
.C(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_35),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_40),
.A2(n_52),
.B(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_43),
.B(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_52),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_44),
.A2(n_52),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_44),
.A2(n_50),
.B(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_44),
.A2(n_52),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_44),
.A2(n_52),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_44),
.A2(n_52),
.B1(n_217),
.B2(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_44),
.B(n_168),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_48),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_52),
.A2(n_61),
.B(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_64),
.A2(n_66),
.B(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_64),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_76),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_80),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_69),
.A2(n_120),
.B1(n_121),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_69),
.A2(n_120),
.B1(n_148),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.C(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_70),
.B(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_70),
.A2(n_77),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_75),
.Y(n_78)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_75),
.B(n_168),
.CON(n_167),
.SN(n_167)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_92),
.B(n_96),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_93),
.B1(n_103),
.B2(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B(n_90),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_86),
.A2(n_89),
.B1(n_138),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_86),
.A2(n_112),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_86),
.A2(n_141),
.B1(n_250),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_87),
.A2(n_91),
.B(n_140),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_87),
.A2(n_88),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_91),
.Y(n_112)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_105),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_104),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_105),
.A2(n_106),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.C(n_118),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_108),
.B(n_113),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_109),
.A2(n_184),
.B(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_123),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_153),
.B(n_301),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_150),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_128),
.B(n_150),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.C(n_135),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_133),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_135),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.C(n_146),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_136),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_142),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_141),
.B(n_168),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_143),
.Y(n_291)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_295),
.B(n_300),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_198),
.B(n_281),
.C(n_294),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_185),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_156),
.B(n_185),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_171),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_158),
.B(n_159),
.C(n_171),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_173),
.B(n_177),
.C(n_180),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_186),
.A2(n_187),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_280),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_273),
.B(n_279),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_228),
.B(n_272),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_219),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_202),
.B(n_219),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_212),
.C(n_215),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_203),
.A2(n_204),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_206),
.Y(n_226)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_226),
.C(n_227),
.Y(n_274)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_266),
.B(n_271),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_246),
.B(n_265),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_238),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_254),
.B(n_264),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_252),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_259),
.B(n_263),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_257),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_292),
.B2(n_293),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.C(n_293),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);


endmodule