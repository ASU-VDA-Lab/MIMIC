module fake_jpeg_3360_n_625 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_625);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_625;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_69),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_9),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_71),
.B(n_109),
.Y(n_174)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_31),
.B(n_9),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_78),
.B(n_87),
.Y(n_166)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_31),
.B(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_33),
.B(n_11),
.Y(n_96)
);

AND2x4_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_45),
.Y(n_124)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_19),
.C(n_18),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_37),
.C(n_54),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_33),
.B(n_19),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_32),
.B1(n_55),
.B2(n_45),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_114),
.A2(n_133),
.B1(n_158),
.B2(n_165),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_124),
.B(n_58),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_51),
.B1(n_42),
.B2(n_39),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_164),
.B1(n_169),
.B2(n_179),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_32),
.B1(n_55),
.B2(n_45),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_59),
.A2(n_37),
.B1(n_54),
.B2(n_20),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_138),
.A2(n_20),
.B1(n_37),
.B2(n_26),
.Y(n_204)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_98),
.A2(n_32),
.B1(n_55),
.B2(n_42),
.Y(n_158)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_103),
.A2(n_52),
.B1(n_39),
.B2(n_51),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_112),
.A2(n_55),
.B1(n_51),
.B2(n_42),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_86),
.A2(n_55),
.B1(n_99),
.B2(n_66),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_55),
.Y(n_183)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_110),
.A2(n_51),
.B1(n_42),
.B2(n_34),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_181),
.B(n_183),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_182),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g276 ( 
.A(n_185),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_97),
.B1(n_85),
.B2(n_106),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_186),
.A2(n_208),
.B1(n_225),
.B2(n_147),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_91),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_189),
.B(n_197),
.Y(n_273)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_20),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_192),
.B(n_212),
.Y(n_257)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_41),
.B1(n_47),
.B2(n_40),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_194),
.A2(n_205),
.B1(n_231),
.B2(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_105),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_117),
.B(n_79),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_198),
.B(n_234),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_124),
.A2(n_111),
.B1(n_88),
.B2(n_101),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g254 ( 
.A1(n_199),
.A2(n_157),
.B1(n_120),
.B2(n_126),
.Y(n_254)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_200),
.Y(n_267)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_115),
.A2(n_60),
.B1(n_84),
.B2(n_104),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_243),
.B(n_204),
.Y(n_246)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_215),
.B1(n_218),
.B2(n_220),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_149),
.A2(n_47),
.B1(n_27),
.B2(n_40),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_34),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_206),
.B(n_213),
.Y(n_293)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_125),
.B(n_26),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_131),
.B(n_49),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_143),
.B(n_26),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_216),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_65),
.B1(n_62),
.B2(n_67),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_48),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_129),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_127),
.A2(n_57),
.B1(n_80),
.B2(n_82),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_48),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_222),
.B(n_227),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g292 ( 
.A(n_223),
.Y(n_292)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_115),
.Y(n_224)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_114),
.A2(n_107),
.B1(n_52),
.B2(n_48),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_146),
.B(n_43),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_120),
.Y(n_228)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_118),
.Y(n_229)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

CKINVDCx12_ASAP7_75t_R g291 ( 
.A(n_230),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_160),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_153),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_108),
.Y(n_235)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_178),
.A2(n_43),
.B1(n_47),
.B2(n_41),
.Y(n_238)
);

AO22x1_ASAP7_75t_SL g239 ( 
.A1(n_133),
.A2(n_108),
.B1(n_102),
.B2(n_90),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_239),
.A2(n_139),
.B1(n_155),
.B2(n_134),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_121),
.Y(n_241)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_140),
.B(n_43),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_159),
.A2(n_57),
.B1(n_100),
.B2(n_83),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_63),
.B1(n_94),
.B2(n_159),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_246),
.B(n_235),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_251),
.A2(n_270),
.B1(n_275),
.B2(n_235),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_254),
.A2(n_262),
.B1(n_280),
.B2(n_50),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_187),
.B(n_52),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_256),
.B(n_260),
.Y(n_309)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_126),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_184),
.A2(n_177),
.B1(n_171),
.B2(n_162),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_183),
.A2(n_145),
.B1(n_134),
.B2(n_139),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_268),
.A2(n_294),
.B1(n_225),
.B2(n_218),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_208),
.A2(n_177),
.B1(n_171),
.B2(n_162),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_186),
.A2(n_242),
.B1(n_227),
.B2(n_239),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_183),
.B(n_207),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_277),
.B(n_283),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_214),
.A2(n_142),
.B1(n_147),
.B2(n_155),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_242),
.A2(n_29),
.B(n_50),
.C(n_145),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_281),
.A2(n_240),
.B(n_236),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_193),
.B(n_156),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_189),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_286),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_289),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_212),
.B(n_156),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_189),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_300),
.Y(n_374)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_242),
.B1(n_222),
.B2(n_216),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_303),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_305),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_200),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

AOI32xp33_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_242),
.A3(n_226),
.B1(n_228),
.B2(n_239),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_320),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_312),
.A2(n_334),
.B1(n_341),
.B2(n_342),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_313),
.A2(n_333),
.B(n_230),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_314),
.A2(n_321),
.B1(n_322),
.B2(n_340),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_273),
.A2(n_237),
.B1(n_229),
.B2(n_221),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_326),
.Y(n_366)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_317),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_255),
.A2(n_201),
.B1(n_217),
.B2(n_185),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_211),
.B1(n_191),
.B2(n_188),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_254),
.B1(n_265),
.B2(n_258),
.Y(n_350)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_327),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_195),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_328),
.B(n_329),
.Y(n_351)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_257),
.B(n_210),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_331),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_188),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_269),
.A2(n_286),
.B(n_253),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_269),
.A2(n_202),
.B1(n_142),
.B2(n_233),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_335),
.B(n_258),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_293),
.B(n_195),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_337),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_180),
.A3(n_191),
.B1(n_241),
.B2(n_50),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_263),
.B(n_180),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_343),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_296),
.A2(n_185),
.B1(n_209),
.B2(n_203),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_246),
.A2(n_232),
.B1(n_50),
.B2(n_29),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_263),
.B(n_288),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_344),
.A2(n_290),
.B1(n_274),
.B2(n_297),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_281),
.A2(n_50),
.B1(n_21),
.B2(n_223),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_345),
.A2(n_348),
.B1(n_276),
.B2(n_252),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_249),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_346),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_288),
.B(n_279),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_274),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_250),
.A2(n_50),
.B1(n_21),
.B2(n_230),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_282),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_349),
.B(n_367),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_368),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_291),
.C(n_248),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_352),
.B(n_392),
.C(n_0),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_347),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_355),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_343),
.Y(n_356)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_303),
.A2(n_254),
.B1(n_289),
.B2(n_285),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_360),
.A2(n_372),
.B1(n_378),
.B2(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_379),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_313),
.A2(n_252),
.B(n_261),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_385),
.B(n_315),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_279),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_339),
.A2(n_289),
.B1(n_276),
.B2(n_271),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_289),
.B1(n_295),
.B2(n_285),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_312),
.A2(n_295),
.B1(n_297),
.B2(n_264),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_305),
.B(n_248),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_380),
.A2(n_391),
.B1(n_316),
.B2(n_323),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_387),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_308),
.A2(n_264),
.B1(n_290),
.B2(n_245),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_390),
.B1(n_311),
.B2(n_302),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_338),
.Y(n_386)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_331),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_245),
.B1(n_271),
.B2(n_261),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_259),
.B1(n_21),
.B2(n_2),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_330),
.B(n_21),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_375),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_394),
.B(n_398),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_332),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_332),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_426),
.C(n_428),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_351),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_400),
.B(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_401),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_388),
.A2(n_316),
.B1(n_345),
.B2(n_334),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_404),
.A2(n_408),
.B(n_409),
.Y(n_438)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_405),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_364),
.Y(n_464)
);

XNOR2x2_ASAP7_75t_SL g407 ( 
.A(n_361),
.B(n_373),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_429),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_371),
.A2(n_309),
.B1(n_342),
.B2(n_348),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_336),
.C(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_321),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_421),
.Y(n_461)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_415),
.B1(n_427),
.B2(n_431),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_358),
.A2(n_329),
.B1(n_335),
.B2(n_320),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_352),
.B(n_369),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_430),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_371),
.A2(n_300),
.B1(n_317),
.B2(n_310),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_383),
.Y(n_453)
);

AO21x2_ASAP7_75t_SL g419 ( 
.A1(n_368),
.A2(n_337),
.B(n_301),
.Y(n_419)
);

AO22x1_ASAP7_75t_SL g444 ( 
.A1(n_419),
.A2(n_372),
.B1(n_390),
.B2(n_350),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_319),
.Y(n_420)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_420),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_374),
.B(n_325),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_307),
.C(n_306),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_422),
.B(n_376),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_386),
.B(n_328),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_424),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_358),
.A2(n_327),
.B1(n_325),
.B2(n_324),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_425),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_18),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_373),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_366),
.B(n_17),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_392),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_360),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_389),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_432),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_407),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_416),
.C(n_430),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_449),
.C(n_451),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_414),
.A2(n_387),
.B1(n_355),
.B2(n_376),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_437),
.A2(n_442),
.B1(n_452),
.B2(n_459),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_413),
.Y(n_440)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_415),
.A2(n_377),
.B1(n_391),
.B2(n_384),
.Y(n_442)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_379),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_448),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_399),
.B(n_382),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_357),
.C(n_382),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_406),
.A2(n_381),
.B(n_357),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_L g495 ( 
.A1(n_450),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_359),
.C(n_370),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_417),
.B1(n_419),
.B2(n_403),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_453),
.B(n_464),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_408),
.A2(n_374),
.B(n_362),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_458),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_411),
.A2(n_419),
.B1(n_403),
.B2(n_397),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_419),
.A2(n_370),
.B1(n_362),
.B2(n_359),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_460),
.A2(n_397),
.B1(n_395),
.B2(n_401),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_354),
.C(n_353),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_463),
.C(n_448),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_402),
.B(n_354),
.C(n_353),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_431),
.A2(n_378),
.B1(n_17),
.B2(n_16),
.Y(n_465)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_420),
.Y(n_468)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_470),
.A2(n_427),
.B1(n_404),
.B2(n_409),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_393),
.Y(n_474)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_475),
.B(n_502),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_396),
.Y(n_477)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_396),
.Y(n_478)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_450),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_479),
.Y(n_527)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_481),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_459),
.A2(n_403),
.B1(n_425),
.B2(n_418),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_483),
.A2(n_489),
.B1(n_497),
.B2(n_440),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_436),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_494),
.Y(n_520)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_488),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_395),
.Y(n_490)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_490),
.Y(n_526)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_457),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_492),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_437),
.B(n_426),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_499),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_428),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_495),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_503),
.C(n_433),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_439),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_455),
.B(n_13),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_461),
.B(n_13),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_449),
.B(n_1),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_456),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_441),
.B(n_3),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_441),
.B(n_3),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_473),
.A2(n_452),
.B1(n_460),
.B2(n_439),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_505),
.A2(n_518),
.B1(n_529),
.B2(n_501),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g542 ( 
.A(n_506),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_508),
.B(n_511),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_509),
.A2(n_513),
.B1(n_524),
.B2(n_472),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_462),
.C(n_451),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_445),
.C(n_458),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_512),
.B(n_514),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_482),
.A2(n_468),
.B1(n_467),
.B2(n_447),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_485),
.A2(n_438),
.B(n_453),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_484),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_515),
.B(n_516),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_433),
.C(n_438),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_434),
.B1(n_467),
.B2(n_453),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_482),
.A2(n_447),
.B1(n_456),
.B2(n_464),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_496),
.B(n_435),
.C(n_469),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_471),
.C(n_494),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_484),
.A2(n_489),
.B1(n_488),
.B2(n_485),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_518),
.B1(n_505),
.B2(n_483),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_532),
.A2(n_534),
.B1(n_537),
.B2(n_510),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_521),
.B(n_490),
.Y(n_533)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_533),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_472),
.Y(n_535)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_535),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_536),
.A2(n_546),
.B1(n_492),
.B2(n_444),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_529),
.A2(n_510),
.B1(n_526),
.B2(n_523),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_516),
.B(n_471),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g572 ( 
.A(n_538),
.B(n_531),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_513),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_543),
.Y(n_561)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_517),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_525),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g557 ( 
.A(n_544),
.B(n_553),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_520),
.B(n_501),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_552),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_509),
.A2(n_493),
.B1(n_442),
.B2(n_481),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_547),
.B(n_549),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_506),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_524),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_522),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_501),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_511),
.B(n_503),
.C(n_502),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_556),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_551),
.A2(n_514),
.B(n_523),
.Y(n_556)
);

BUFx24_ASAP7_75t_SL g558 ( 
.A(n_550),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_558),
.B(n_4),
.Y(n_589)
);

AOI21xp33_ASAP7_75t_L g559 ( 
.A1(n_548),
.A2(n_519),
.B(n_504),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_559),
.A2(n_542),
.B(n_507),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_539),
.B(n_528),
.C(n_512),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_569),
.Y(n_574)
);

FAx1_ASAP7_75t_SL g563 ( 
.A(n_534),
.B(n_475),
.CI(n_531),
.CON(n_563),
.SN(n_563)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_563),
.B(n_565),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_566),
.A2(n_536),
.B1(n_546),
.B2(n_547),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_508),
.C(n_444),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_532),
.A2(n_537),
.B1(n_540),
.B2(n_533),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_570),
.A2(n_491),
.B1(n_497),
.B2(n_530),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_552),
.C(n_538),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_553),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_572),
.B(n_495),
.Y(n_585)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_573),
.Y(n_593)
);

AOI31xp33_ASAP7_75t_L g590 ( 
.A1(n_576),
.A2(n_579),
.A3(n_571),
.B(n_574),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_577),
.B(n_583),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_567),
.A2(n_549),
.B1(n_535),
.B2(n_541),
.Y(n_578)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_578),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_560),
.A2(n_504),
.B(n_530),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_569),
.B(n_491),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_580),
.B(n_588),
.Y(n_602)
);

AOI22x1_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_584),
.B1(n_563),
.B2(n_572),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_480),
.Y(n_583)
);

XOR2x2_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_470),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_585),
.B(n_557),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_568),
.B(n_480),
.Y(n_586)
);

AO21x1_ASAP7_75t_L g594 ( 
.A1(n_586),
.A2(n_556),
.B(n_561),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_555),
.B(n_3),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_587),
.B(n_589),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_3),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_590),
.B(n_594),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_580),
.B(n_554),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_595),
.B(n_596),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_581),
.B(n_566),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_581),
.A2(n_563),
.B(n_562),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_597),
.A2(n_575),
.B(n_578),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_599),
.B(n_600),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_575),
.B(n_4),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_601),
.B(n_4),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_603),
.A2(n_608),
.B1(n_592),
.B2(n_602),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_593),
.A2(n_584),
.B1(n_586),
.B2(n_573),
.Y(n_606)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_606),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_597),
.A2(n_585),
.B(n_588),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_609),
.A2(n_610),
.B(n_599),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_5),
.C(n_6),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_604),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_612),
.B(n_613),
.C(n_614),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_607),
.A2(n_598),
.B1(n_594),
.B2(n_600),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_615),
.B(n_607),
.C(n_605),
.Y(n_617)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_617),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_611),
.B(n_602),
.C(n_6),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_618),
.B(n_5),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_620),
.A2(n_616),
.B(n_7),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_621),
.A2(n_619),
.B(n_7),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_622),
.B(n_6),
.C(n_8),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_8),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g625 ( 
.A1(n_624),
.A2(n_8),
.B(n_477),
.Y(n_625)
);


endmodule