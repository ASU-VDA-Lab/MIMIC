module fake_jpeg_30960_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_4),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_0),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_19),
.B(n_37),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_59),
.A3(n_54),
.B1(n_46),
.B2(n_49),
.Y(n_63)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_17),
.B(n_35),
.C(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_50),
.B1(n_43),
.B2(n_40),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_42),
.B1(n_22),
.B2(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_49),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_51),
.B(n_53),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_3),
.B(n_6),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_21),
.B1(n_31),
.B2(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_7),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_8),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_73),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_97),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_14),
.C(n_15),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_16),
.C(n_20),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_76),
.B(n_75),
.C(n_26),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_103),
.B1(n_94),
.B2(n_30),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_99),
.C(n_90),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_105),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_109),
.B(n_110),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_102),
.C(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_38),
.Y(n_114)
);


endmodule