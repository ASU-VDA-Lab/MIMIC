module fake_netlist_6_2064_n_2441 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2441);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2441;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_2127;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g226 ( 
.A(n_76),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_182),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_122),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_102),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_99),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_65),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_83),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_30),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_171),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_92),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_10),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_98),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_13),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_196),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_170),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_223),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_162),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_115),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_103),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_109),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_72),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_184),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_66),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_117),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_46),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_27),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_138),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_80),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_59),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_63),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_78),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_67),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_202),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_67),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_66),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_150),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_125),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_76),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_68),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_10),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_84),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_103),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_126),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_83),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_166),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_85),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_70),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_136),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_177),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_190),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_62),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_132),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_199),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_78),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_215),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_218),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_119),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_130),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_174),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_18),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_207),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_208),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_33),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_95),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_169),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_146),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_55),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_121),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_189),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_62),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_53),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_29),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_20),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_68),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_71),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_188),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_6),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_172),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_157),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_42),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_158),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_60),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_106),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_159),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_13),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_71),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_133),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_197),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_183),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_79),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_19),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_75),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_53),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_37),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_96),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_113),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_41),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_141),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_154),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_191),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_35),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_225),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_107),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_120),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_28),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_44),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_0),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_23),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_54),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_142),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_161),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_101),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_3),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_212),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_211),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_40),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_73),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_93),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_43),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_8),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_128),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_144),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_40),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_31),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_137),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_143),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_23),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_18),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_99),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_155),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_59),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_69),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_153),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_28),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_206),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_114),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_135),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_112),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_60),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_145),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_43),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_34),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_193),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_6),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_8),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_14),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_95),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_85),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_33),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_131),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_179),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_15),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_57),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_14),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_92),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_100),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_42),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_147),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_31),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_1),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_149),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_65),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_106),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_35),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_178),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_198),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_209),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_201),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_57),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_2),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_186),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_25),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_140),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_4),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_217),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_101),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_84),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_164),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_24),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_74),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_185),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_15),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_118),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_221),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_17),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_58),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_80),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_216),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_11),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_192),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_16),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_24),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_316),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_228),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_229),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_316),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_234),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_316),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_362),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_316),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_245),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_246),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_227),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_316),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_249),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_226),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_251),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_252),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_360),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_253),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_254),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_269),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_257),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_226),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_259),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_398),
.B(n_0),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_227),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_261),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_360),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_264),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_265),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_316),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_316),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_267),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_316),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_269),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_316),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_316),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_226),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_275),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_270),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_304),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_279),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_289),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_395),
.B(n_2),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_270),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_270),
.Y(n_493)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_247),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_280),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_288),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_445),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_232),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_278),
.B(n_5),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_293),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_347),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_294),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_233),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_243),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_230),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_295),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_244),
.B(n_5),
.Y(n_508)
);

BUFx2_ASAP7_75t_SL g509 ( 
.A(n_244),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_347),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_347),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_365),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_227),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_365),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_296),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_365),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_299),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_304),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_400),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_304),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_300),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_355),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_305),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_308),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_278),
.B(n_7),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_355),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_355),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_230),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_371),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_310),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_371),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_277),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_371),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_236),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_314),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_317),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_232),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_319),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_335),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_439),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_236),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_338),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_266),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_266),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_340),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_268),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_351),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_315),
.B(n_9),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_268),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_271),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_R g555 ( 
.A(n_352),
.B(n_11),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_271),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_324),
.B(n_12),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_274),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_274),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_276),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_356),
.Y(n_561)
);

INVxp33_ASAP7_75t_SL g562 ( 
.A(n_235),
.Y(n_562)
);

BUFx6f_ASAP7_75t_SL g563 ( 
.A(n_247),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_363),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_276),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_447),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_545),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_456),
.B(n_315),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_490),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_452),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_454),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_545),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_465),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_547),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_459),
.B(n_467),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_448),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_548),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_479),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_456),
.B(n_378),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_490),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_548),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_456),
.B(n_378),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_480),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_470),
.B(n_418),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_557),
.B(n_324),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_534),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_550),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_550),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_490),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_488),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_446),
.A2(n_298),
.B(n_239),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_459),
.B(n_467),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_450),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_455),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_446),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_R g601 ( 
.A(n_494),
.B(n_366),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_470),
.B(n_418),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_468),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_495),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_509),
.B(n_508),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_470),
.B(n_367),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_500),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_502),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_553),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_458),
.B(n_373),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_513),
.B(n_374),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_488),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_465),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_513),
.B(n_377),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_449),
.Y(n_617)
);

AND3x2_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_552),
.C(n_491),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_519),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_449),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_R g621 ( 
.A(n_462),
.B(n_444),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_513),
.B(n_382),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_554),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_469),
.B(n_358),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_460),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_461),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_451),
.Y(n_627)
);

OA21x2_ASAP7_75t_L g628 ( 
.A1(n_484),
.A2(n_298),
.B(n_239),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_522),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_498),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_451),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_463),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_453),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_453),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_457),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_509),
.B(n_286),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_457),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_506),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_475),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_464),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_558),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_508),
.B(n_286),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_475),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_532),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_558),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_483),
.B(n_385),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_476),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_R g650 ( 
.A(n_466),
.B(n_389),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_476),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_478),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_522),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_472),
.A2(n_242),
.B1(n_250),
.B2(n_241),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_559),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_504),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_504),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_538),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_R g659 ( 
.A(n_503),
.B(n_237),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_524),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_600),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_570),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_631),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_593),
.B(n_472),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_600),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_576),
.B(n_483),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_631),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_636),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_573),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_562),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_576),
.B(n_524),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_600),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_624),
.B(n_471),
.Y(n_673)
);

BUFx4f_ASAP7_75t_L g674 ( 
.A(n_636),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_631),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_593),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_636),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_617),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_573),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_576),
.B(n_528),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_605),
.B(n_473),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_644),
.A2(n_527),
.B1(n_499),
.B2(n_312),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_624),
.A2(n_555),
.B1(n_358),
.B2(n_469),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_605),
.B(n_474),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_571),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_573),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_631),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_617),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_595),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_617),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_620),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_620),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_595),
.B(n_528),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_566),
.B(n_546),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_573),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_587),
.A2(n_321),
.B1(n_341),
.B2(n_301),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_595),
.B(n_529),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_620),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_648),
.B(n_477),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_640),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_627),
.Y(n_702)
);

AND3x2_ASAP7_75t_L g703 ( 
.A(n_638),
.B(n_309),
.C(n_306),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_573),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_630),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_570),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_648),
.B(n_486),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_573),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_630),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_606),
.B(n_489),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_640),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_627),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_627),
.Y(n_713)
);

AND2x6_ASAP7_75t_SL g714 ( 
.A(n_638),
.B(n_281),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_636),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_587),
.B(n_339),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_632),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_636),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_635),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_606),
.B(n_496),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_636),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_630),
.B(n_339),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_653),
.B(n_339),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_601),
.B(n_515),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_653),
.B(n_231),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_635),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_574),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_578),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_601),
.B(n_518),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_653),
.B(n_231),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_596),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_660),
.B(n_529),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_628),
.B(n_307),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_596),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_611),
.B(n_523),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_636),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_611),
.B(n_525),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_571),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_612),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_596),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_621),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_616),
.B(n_526),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_616),
.B(n_622),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_621),
.A2(n_429),
.B1(n_399),
.B2(n_238),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_635),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_612),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_641),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_622),
.B(n_537),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_641),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_660),
.B(n_531),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_596),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_641),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_645),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_568),
.B(n_239),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_596),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_574),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_598),
.B(n_541),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_645),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_625),
.B(n_543),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_568),
.B(n_549),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_SL g766 ( 
.A(n_657),
.B(n_563),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_651),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_596),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_615),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_651),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_610),
.B(n_564),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_651),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_652),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_581),
.B(n_478),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_652),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_581),
.B(n_481),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_610),
.B(n_551),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_584),
.B(n_481),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_657),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_652),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_637),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_596),
.Y(n_782)
);

AO22x2_ASAP7_75t_L g783 ( 
.A1(n_618),
.A2(n_312),
.B1(n_313),
.B2(n_243),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_615),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_660),
.B(n_248),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_626),
.B(n_561),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_637),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_603),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_584),
.B(n_482),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_619),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_594),
.B(n_248),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_613),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_637),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_654),
.A2(n_240),
.B1(n_256),
.B2(n_255),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_637),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_657),
.B(n_531),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_586),
.B(n_482),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_637),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_637),
.Y(n_800)
);

AND2x2_ASAP7_75t_SL g801 ( 
.A(n_628),
.B(n_298),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_650),
.B(n_247),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_639),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_594),
.B(n_272),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_639),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_619),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_SL g807 ( 
.A(n_656),
.B(n_563),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_613),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_633),
.B(n_642),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_639),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_586),
.B(n_348),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_639),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_L g813 ( 
.A(n_650),
.B(n_602),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_639),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_580),
.B(n_507),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_639),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_588),
.A2(n_260),
.B1(n_262),
.B2(n_258),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_639),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_618),
.A2(n_313),
.B1(n_536),
.B2(n_530),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_656),
.B(n_247),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_649),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_567),
.B(n_533),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_649),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_822),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_670),
.B(n_588),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_747),
.B(n_602),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_666),
.B(n_530),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_801),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_711),
.Y(n_829)
);

OAI221xp5_ASAP7_75t_L g830 ( 
.A1(n_683),
.A2(n_536),
.B1(n_654),
.B2(n_507),
.C(n_384),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_822),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_666),
.B(n_585),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_717),
.A2(n_582),
.B(n_569),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_690),
.B(n_649),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_718),
.A2(n_659),
.B1(n_585),
.B2(n_580),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_700),
.B(n_649),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_736),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_707),
.B(n_649),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_690),
.B(n_649),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_801),
.B(n_649),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_682),
.B(n_585),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_671),
.B(n_533),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_791),
.A2(n_354),
.B1(n_387),
.B2(n_348),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_659),
.C(n_273),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_736),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_664),
.B(n_603),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_791),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_801),
.B(n_289),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_671),
.B(n_569),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_685),
.A2(n_307),
.B1(n_330),
.B2(n_311),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_724),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_754),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_680),
.B(n_535),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_754),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_705),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_680),
.B(n_535),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_745),
.B(n_604),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_694),
.B(n_569),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_791),
.B(n_348),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_684),
.A2(n_572),
.B(n_575),
.C(n_567),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_791),
.A2(n_387),
.B1(n_354),
.B2(n_628),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_705),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_765),
.B(n_604),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_694),
.B(n_582),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_698),
.B(n_582),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_804),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_774),
.B(n_289),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_699),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_710),
.B(n_607),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_813),
.A2(n_330),
.B1(n_311),
.B2(n_390),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_716),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_709),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_718),
.A2(n_272),
.B1(n_327),
.B2(n_323),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_779),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_804),
.A2(n_387),
.B(n_354),
.C(n_327),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_709),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_698),
.B(n_591),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_716),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_812),
.A2(n_592),
.B(n_591),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_722),
.B(n_607),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_724),
.Y(n_882)
);

NOR2x1p5_ASAP7_75t_L g883 ( 
.A(n_815),
.B(n_608),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_739),
.B(n_591),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_779),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_724),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_741),
.B(n_608),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_776),
.B(n_289),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_746),
.B(n_752),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_724),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_804),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_778),
.B(n_592),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_789),
.B(n_592),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_798),
.B(n_289),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_673),
.B(n_658),
.C(n_646),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_718),
.A2(n_402),
.B1(n_403),
.B2(n_392),
.Y(n_896)
);

BUFx5_ASAP7_75t_L g897 ( 
.A(n_823),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_804),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_762),
.B(n_646),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_718),
.B(n_323),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_725),
.B(n_332),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_719),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_725),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_797),
.B(n_540),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_719),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_764),
.B(n_658),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_718),
.B(n_332),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_725),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_725),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_727),
.B(n_572),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_662),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_816),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_737),
.B(n_388),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_721),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_797),
.B(n_540),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_820),
.B(n_563),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_727),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_737),
.B(n_289),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_737),
.B(n_388),
.Y(n_920)
);

AND2x6_ASAP7_75t_SL g921 ( 
.A(n_786),
.B(n_281),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_721),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_664),
.B(n_563),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_687),
.Y(n_924)
);

BUFx8_ASAP7_75t_L g925 ( 
.A(n_743),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_727),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_743),
.B(n_542),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_733),
.B(n_785),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_750),
.B(n_542),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_733),
.B(n_785),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_733),
.B(n_417),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_758),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_783),
.A2(n_420),
.B1(n_424),
.B2(n_410),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_733),
.B(n_417),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_758),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_785),
.B(n_421),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_785),
.B(n_421),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_661),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_770),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_793),
.B(n_428),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_793),
.B(n_428),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_661),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_796),
.B(n_443),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_771),
.B(n_505),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_770),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_695),
.A2(n_302),
.B1(n_413),
.B2(n_350),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_665),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_750),
.B(n_263),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_761),
.B(n_544),
.C(n_283),
.Y(n_949)
);

NOR2x1p5_ASAP7_75t_L g950 ( 
.A(n_815),
.B(n_282),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_783),
.B(n_285),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_772),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_665),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_759),
.B(n_575),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_772),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_816),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_796),
.B(n_577),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_799),
.B(n_577),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_672),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_SL g960 ( 
.A(n_687),
.B(n_329),
.Y(n_960)
);

BUFx6f_ASAP7_75t_SL g961 ( 
.A(n_730),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_773),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_799),
.B(n_579),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_800),
.B(n_579),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_672),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_676),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_783),
.A2(n_431),
.B1(n_434),
.B2(n_426),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_678),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_781),
.B(n_329),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_781),
.B(n_329),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_730),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_800),
.B(n_583),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_759),
.A2(n_628),
.B1(n_329),
.B2(n_291),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_773),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_784),
.B(n_790),
.Y(n_975)
);

AND2x2_ASAP7_75t_SL g976 ( 
.A(n_748),
.B(n_329),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_784),
.B(n_284),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_759),
.A2(n_329),
.B1(n_232),
.B2(n_291),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_803),
.B(n_810),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_803),
.B(n_583),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_783),
.A2(n_441),
.B1(n_437),
.B2(n_436),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_810),
.B(n_814),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_L g983 ( 
.A(n_814),
.B(n_232),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_759),
.A2(n_232),
.B1(n_291),
.B2(n_405),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_811),
.A2(n_766),
.B1(n_802),
.B2(n_790),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_818),
.B(n_589),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_811),
.A2(n_232),
.B1(n_291),
.B2(n_405),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_806),
.B(n_232),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_678),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_794),
.A2(n_285),
.B(n_303),
.C(n_328),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_775),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_L g992 ( 
.A(n_794),
.B(n_290),
.C(n_287),
.Y(n_992)
);

INVx8_ASAP7_75t_L g993 ( 
.A(n_811),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_748),
.A2(n_328),
.B(n_432),
.C(n_427),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_689),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_818),
.B(n_589),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_687),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_858),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_875),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_828),
.B(n_730),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_829),
.Y(n_1001)
);

AND2x2_ASAP7_75t_SL g1002 ( 
.A(n_976),
.B(n_761),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_828),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_858),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_993),
.B(n_811),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_827),
.B(n_806),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_SL g1007 ( 
.A(n_830),
.B(n_742),
.C(n_686),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_867),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_869),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_971),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_911),
.B(n_811),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_825),
.B(n_792),
.C(n_729),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_SL g1013 ( 
.A(n_835),
.B(n_742),
.C(n_686),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_867),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_889),
.B(n_809),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_826),
.B(n_821),
.Y(n_1016)
);

INVx5_ASAP7_75t_L g1017 ( 
.A(n_828),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_911),
.B(n_855),
.Y(n_1018)
);

AO22x1_ASAP7_75t_L g1019 ( 
.A1(n_828),
.A2(n_769),
.B1(n_817),
.B2(n_337),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_829),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_910),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_976),
.A2(n_691),
.B1(n_692),
.B2(n_689),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_869),
.Y(n_1023)
);

CKINVDCx8_ASAP7_75t_R g1024 ( 
.A(n_921),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_828),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_827),
.B(n_735),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_872),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_918),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_926),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_925),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_911),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_832),
.B(n_735),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_882),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_925),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_885),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_842),
.B(n_821),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_971),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_925),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_898),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_872),
.Y(n_1040)
);

AOI22x1_ASAP7_75t_L g1041 ( 
.A1(n_842),
.A2(n_775),
.B1(n_692),
.B2(n_693),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_853),
.B(n_823),
.Y(n_1042)
);

AND2x2_ASAP7_75t_SL g1043 ( 
.A(n_978),
.B(n_697),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_966),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_832),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_863),
.B(n_777),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_879),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_853),
.B(n_691),
.Y(n_1048)
);

CKINVDCx8_ASAP7_75t_R g1049 ( 
.A(n_899),
.Y(n_1049)
);

OR2x2_ASAP7_75t_SL g1050 ( 
.A(n_844),
.B(n_992),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_841),
.B(n_808),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_890),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_898),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_898),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_908),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_856),
.B(n_735),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_909),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_856),
.B(n_904),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_898),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_961),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_944),
.B(n_726),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_904),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_938),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_879),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_916),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_942),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_898),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_947),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_916),
.B(n_693),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_997),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_953),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_959),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_997),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_951),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_985),
.B(n_732),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_837),
.B(n_702),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_902),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_965),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_873),
.B(n_703),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_902),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_997),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_SL g1082 ( 
.A1(n_906),
.A2(n_706),
.B1(n_788),
.B2(n_701),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_847),
.B(n_677),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_905),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_905),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_948),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_847),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_912),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_824),
.B(n_697),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_845),
.B(n_702),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_968),
.Y(n_1091)
);

AOI22x1_ASAP7_75t_L g1092 ( 
.A1(n_847),
.A2(n_713),
.B1(n_715),
.B2(n_712),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_877),
.B(n_787),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_SL g1094 ( 
.A(n_994),
.B(n_788),
.C(n_297),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_997),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_R g1096 ( 
.A(n_846),
.B(n_857),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_891),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_997),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_891),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_917),
.B(n_544),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_989),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_995),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_951),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_891),
.Y(n_1104)
);

BUFx4f_ASAP7_75t_L g1105 ( 
.A(n_993),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_SL g1106 ( 
.A(n_994),
.B(n_318),
.C(n_292),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_915),
.Y(n_1107)
);

AOI22x1_ASAP7_75t_L g1108 ( 
.A1(n_915),
.A2(n_713),
.B1(n_715),
.B2(n_712),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_951),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_852),
.B(n_728),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_922),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_854),
.B(n_728),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_836),
.B(n_749),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_961),
.B(n_807),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_961),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_922),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_870),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_831),
.B(n_749),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_927),
.B(n_751),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_954),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_932),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_993),
.B(n_590),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_932),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_851),
.A2(n_787),
.B1(n_753),
.B2(n_756),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_935),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_862),
.A2(n_674),
.B(n_677),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_927),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_851),
.A2(n_787),
.B1(n_753),
.B2(n_756),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_951),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_957),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_958),
.Y(n_1131)
);

AND2x6_ASAP7_75t_L g1132 ( 
.A(n_954),
.B(n_751),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_954),
.A2(n_763),
.B1(n_767),
.B2(n_757),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_977),
.Y(n_1134)
);

INVx6_ASAP7_75t_L g1135 ( 
.A(n_993),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_963),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_860),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_R g1138 ( 
.A(n_881),
.B(n_714),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_913),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_887),
.B(n_677),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_864),
.B(n_674),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_838),
.B(n_757),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_929),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_846),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_964),
.Y(n_1145)
);

AND2x6_ASAP7_75t_L g1146 ( 
.A(n_928),
.B(n_763),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_975),
.B(n_674),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_900),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_972),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_929),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_886),
.B(n_590),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_R g1152 ( 
.A(n_923),
.B(n_669),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_886),
.A2(n_780),
.B1(n_767),
.B2(n_723),
.Y(n_1153)
);

CKINVDCx11_ASAP7_75t_R g1154 ( 
.A(n_900),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_SL g1155 ( 
.A(n_848),
.B(n_687),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_900),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_861),
.A2(n_780),
.B(n_667),
.C(n_675),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_R g1158 ( 
.A(n_903),
.B(n_669),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_849),
.B(n_859),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_900),
.B(n_599),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_980),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_975),
.B(n_720),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_986),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_903),
.B(n_599),
.Y(n_1164)
);

AND2x6_ASAP7_75t_SL g1165 ( 
.A(n_907),
.B(n_303),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_850),
.A2(n_860),
.B1(n_848),
.B2(n_907),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_860),
.Y(n_1167)
);

OR2x2_ASAP7_75t_SL g1168 ( 
.A(n_946),
.B(n_337),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_860),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_950),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_L g1171 ( 
.A(n_860),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_L g1172 ( 
.A(n_883),
.B(n_669),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_871),
.A2(n_667),
.B(n_675),
.C(n_663),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_924),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_996),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_933),
.B(n_720),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_865),
.B(n_679),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_935),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_907),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_939),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_866),
.B(n_679),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_939),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_945),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_945),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_896),
.B(n_687),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_952),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_924),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_878),
.B(n_679),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_967),
.B(n_708),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_981),
.B(n_720),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_952),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_839),
.B(n_696),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1015),
.B(n_990),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1017),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1030),
.Y(n_1195)
);

AOI211x1_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_1019),
.B(n_1089),
.C(n_1075),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1017),
.B(n_840),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1006),
.B(n_990),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1113),
.A2(n_920),
.B(n_914),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_998),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_998),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1086),
.B(n_988),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1134),
.A2(n_930),
.B(n_884),
.C(n_901),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1030),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1043),
.A2(n_931),
.B(n_936),
.C(n_934),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1006),
.B(n_843),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1056),
.B(n_895),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1008),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1159),
.A2(n_840),
.B(n_919),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1004),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_999),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1041),
.A2(n_919),
.B(n_876),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1127),
.B(n_988),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1142),
.A2(n_888),
.B(n_868),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1041),
.A2(n_941),
.B(n_940),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1141),
.A2(n_937),
.B(n_943),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_SL g1217 ( 
.A(n_1117),
.B(n_949),
.C(n_322),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1014),
.Y(n_1218)
);

O2A1O1Ixp5_ASAP7_75t_SL g1219 ( 
.A1(n_1061),
.A2(n_888),
.B(n_894),
.C(n_868),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_1017),
.B(n_913),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1045),
.B(n_907),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1126),
.A2(n_924),
.B(n_913),
.Y(n_1222)
);

AO21x1_ASAP7_75t_L g1223 ( 
.A1(n_1155),
.A2(n_894),
.B(n_874),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1092),
.A2(n_982),
.B(n_979),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1174),
.A2(n_924),
.B(n_956),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1174),
.A2(n_924),
.B(n_956),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1092),
.A2(n_834),
.B(n_833),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1108),
.A2(n_834),
.B(n_880),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1120),
.B(n_860),
.Y(n_1229)
);

BUFx2_ASAP7_75t_SL g1230 ( 
.A(n_1017),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1045),
.B(n_1119),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1187),
.A2(n_893),
.B(n_892),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_1192),
.B(n_1181),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_999),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1107),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1127),
.B(n_955),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_SL g1237 ( 
.A(n_1017),
.B(n_955),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1025),
.A2(n_740),
.B(n_723),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1004),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1140),
.B(n_962),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1143),
.B(n_962),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1003),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1150),
.B(n_991),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_1003),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1187),
.A2(n_795),
.B(n_740),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1003),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1130),
.B(n_974),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1002),
.A2(n_973),
.B1(n_987),
.B2(n_984),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1024),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1003),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1144),
.B(n_974),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1003),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1051),
.A2(n_325),
.B(n_320),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1035),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1131),
.B(n_991),
.Y(n_1255)
);

NAND2x1_ASAP7_75t_L g1256 ( 
.A(n_1025),
.B(n_696),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1177),
.A2(n_970),
.B(n_969),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1136),
.B(n_897),
.Y(n_1258)
);

NOR2xp67_ASAP7_75t_SL g1259 ( 
.A(n_1059),
.B(n_969),
.Y(n_1259)
);

AND3x4_ASAP7_75t_L g1260 ( 
.A(n_1012),
.B(n_350),
.C(n_302),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1145),
.B(n_897),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1149),
.B(n_897),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1188),
.A2(n_970),
.B(n_704),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1083),
.A2(n_704),
.B(n_696),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1009),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1161),
.B(n_897),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1016),
.A2(n_983),
.B(n_681),
.Y(n_1267)
);

AOI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1117),
.A2(n_983),
.B(n_331),
.Y(n_1268)
);

NOR4xp25_ASAP7_75t_L g1269 ( 
.A(n_1049),
.B(n_343),
.C(n_407),
.D(n_404),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1066),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1039),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1083),
.A2(n_738),
.B(n_704),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1171),
.A2(n_805),
.B(n_795),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1083),
.A2(n_755),
.B(n_738),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_SL g1275 ( 
.A1(n_1025),
.A2(n_805),
.B(n_795),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1139),
.A2(n_755),
.B(n_738),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1119),
.B(n_1062),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1138),
.A2(n_333),
.B(n_326),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1163),
.B(n_897),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1010),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1139),
.A2(n_760),
.B(n_755),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1139),
.A2(n_1189),
.B(n_1042),
.Y(n_1282)
);

INVx5_ASAP7_75t_L g1283 ( 
.A(n_1039),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1175),
.B(n_897),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1035),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1173),
.B(n_1036),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1009),
.A2(n_760),
.B(n_681),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1039),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1010),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1023),
.A2(n_760),
.B(n_688),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1043),
.A2(n_346),
.B(n_432),
.C(n_427),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1001),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1065),
.B(n_897),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1056),
.B(n_663),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1118),
.B(n_688),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1039),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1118),
.B(n_609),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1171),
.A2(n_805),
.B(n_731),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1176),
.A2(n_343),
.B(n_425),
.C(n_422),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1023),
.A2(n_485),
.B(n_484),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1171),
.A2(n_731),
.B(n_708),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1089),
.B(n_609),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1027),
.A2(n_487),
.B(n_485),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1120),
.B(n_614),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1048),
.A2(n_960),
.B(n_539),
.Y(n_1305)
);

NOR2x1_ASAP7_75t_SL g1306 ( 
.A(n_1059),
.B(n_708),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1190),
.A2(n_353),
.A3(n_368),
.B(n_370),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1027),
.A2(n_1047),
.B(n_1040),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1040),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1155),
.A2(n_353),
.B(n_346),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1047),
.A2(n_492),
.B(n_487),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1066),
.B(n_1091),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1037),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1059),
.A2(n_731),
.B(n_708),
.Y(n_1314)
);

NAND2x1_ASAP7_75t_L g1315 ( 
.A(n_1095),
.B(n_708),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1059),
.A2(n_734),
.B(n_731),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1022),
.A2(n_960),
.B(n_539),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1064),
.A2(n_493),
.B(n_492),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_SL g1319 ( 
.A(n_1059),
.B(n_731),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_R g1320 ( 
.A(n_1001),
.B(n_334),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1091),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1044),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1063),
.B(n_614),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1185),
.A2(n_744),
.B(n_734),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1064),
.A2(n_497),
.B(n_493),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1077),
.A2(n_501),
.B(n_497),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1088),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1069),
.A2(n_744),
.B(n_734),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1068),
.B(n_623),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1077),
.A2(n_510),
.B(n_501),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1080),
.A2(n_511),
.B(n_510),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1054),
.A2(n_744),
.B(n_734),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1020),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1080),
.A2(n_512),
.B(n_511),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1007),
.B(n_342),
.C(n_336),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1147),
.A2(n_623),
.B(n_655),
.C(n_647),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1084),
.A2(n_514),
.B(n_512),
.Y(n_1337)
);

OAI22x1_ASAP7_75t_L g1338 ( 
.A1(n_1074),
.A2(n_383),
.B1(n_368),
.B2(n_425),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1049),
.B(n_344),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1162),
.A2(n_383),
.A3(n_422),
.B(n_416),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1166),
.A2(n_375),
.B(n_370),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1133),
.A2(n_1128),
.B(n_1124),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1037),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1002),
.B(n_629),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1071),
.B(n_629),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1084),
.A2(n_516),
.B(n_514),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1046),
.B(n_1011),
.Y(n_1347)
);

NAND2x1p5_ASAP7_75t_L g1348 ( 
.A(n_1105),
.B(n_668),
.Y(n_1348)
);

AOI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1076),
.A2(n_539),
.B(n_498),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1011),
.B(n_634),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1085),
.A2(n_517),
.B(n_516),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1085),
.A2(n_520),
.B(n_517),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1072),
.B(n_634),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1095),
.A2(n_744),
.B(n_734),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1095),
.A2(n_768),
.B(n_744),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1011),
.A2(n_782),
.B(n_768),
.Y(n_1356)
);

INVx5_ASAP7_75t_SL g1357 ( 
.A(n_1005),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1151),
.A2(n_498),
.B(n_643),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1107),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1111),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1287),
.A2(n_1000),
.B(n_1121),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1249),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1254),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1254),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1287),
.A2(n_1123),
.B(n_1121),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1260),
.A2(n_1024),
.B1(n_1168),
.B2(n_1020),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1290),
.A2(n_1272),
.B(n_1264),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1290),
.A2(n_1125),
.B(n_1123),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1194),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1233),
.A2(n_1110),
.B(n_1090),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1264),
.A2(n_1180),
.B(n_1125),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1339),
.B(n_1096),
.C(n_1013),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1277),
.B(n_1046),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1231),
.B(n_1151),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1272),
.A2(n_1182),
.B(n_1180),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1270),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1200),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1274),
.A2(n_1191),
.B(n_1182),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1200),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1230),
.B(n_1135),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1274),
.A2(n_1191),
.B(n_1112),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1308),
.A2(n_1116),
.B(n_1111),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1193),
.A2(n_1115),
.B1(n_1060),
.B2(n_1088),
.Y(n_1383)
);

NOR2x1_ASAP7_75t_R g1384 ( 
.A(n_1195),
.B(n_1034),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1231),
.B(n_1151),
.Y(n_1385)
);

CKINVDCx16_ASAP7_75t_R g1386 ( 
.A(n_1195),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1207),
.A2(n_1026),
.B(n_1032),
.C(n_1170),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1211),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1286),
.A2(n_1100),
.B(n_1152),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1310),
.A2(n_1153),
.B(n_1106),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1285),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1310),
.A2(n_1028),
.B(n_1021),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1321),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1211),
.Y(n_1394)
);

BUFx2_ASAP7_75t_SL g1395 ( 
.A(n_1271),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1209),
.A2(n_1029),
.B(n_1094),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1312),
.A2(n_1050),
.B1(n_1105),
.B2(n_1135),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1271),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1308),
.A2(n_1186),
.B(n_1116),
.Y(n_1399)
);

OR2x6_ASAP7_75t_L g1400 ( 
.A(n_1230),
.B(n_1135),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1341),
.A2(n_1067),
.B(n_1172),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1222),
.A2(n_1228),
.B(n_1227),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1235),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1201),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1341),
.A2(n_1067),
.B(n_1052),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1322),
.B(n_1234),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1208),
.Y(n_1407)
);

OAI222xp33_ASAP7_75t_L g1408 ( 
.A1(n_1248),
.A2(n_1082),
.B1(n_1198),
.B2(n_1347),
.C1(n_1344),
.C2(n_1302),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1344),
.B(n_1050),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1234),
.B(n_1168),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1277),
.B(n_1046),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1218),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1297),
.B(n_1018),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1260),
.A2(n_1031),
.B1(n_1018),
.B2(n_1074),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1228),
.A2(n_1186),
.B(n_1183),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1201),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1235),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1359),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1227),
.A2(n_1184),
.B(n_1178),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1221),
.A2(n_1018),
.B1(n_1109),
.B2(n_1129),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1276),
.A2(n_1097),
.B(n_1087),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1276),
.A2(n_1281),
.B(n_1212),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1292),
.A2(n_1115),
.B1(n_1060),
.B2(n_1160),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1280),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1359),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1281),
.A2(n_1097),
.B(n_1087),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1212),
.A2(n_1097),
.B(n_1087),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1205),
.A2(n_1164),
.B(n_1055),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1282),
.A2(n_1099),
.B(n_1057),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1350),
.B(n_1164),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1221),
.A2(n_1109),
.B1(n_1129),
.B2(n_1079),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1360),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1210),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1271),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1210),
.Y(n_1435)
);

OR2x6_ASAP7_75t_SL g1436 ( 
.A(n_1292),
.B(n_1333),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1268),
.A2(n_1079),
.B1(n_1103),
.B2(n_1156),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1282),
.A2(n_1099),
.B(n_1033),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1239),
.Y(n_1439)
);

INVx5_ASAP7_75t_L g1440 ( 
.A(n_1194),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1217),
.A2(n_1079),
.B1(n_1103),
.B2(n_1160),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1253),
.A2(n_1179),
.B1(n_1156),
.B2(n_1148),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1202),
.A2(n_1105),
.B1(n_1135),
.B2(n_1167),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1327),
.A2(n_1034),
.B1(n_1114),
.B2(n_1038),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1194),
.B(n_1067),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1239),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1229),
.B(n_1122),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1299),
.A2(n_1291),
.B(n_1342),
.C(n_1203),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1233),
.A2(n_1101),
.B(n_1078),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_L g1450 ( 
.A(n_1271),
.B(n_1039),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1304),
.B(n_1019),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1333),
.A2(n_1160),
.B1(n_1148),
.B2(n_1179),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1271),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1263),
.A2(n_1099),
.B(n_1053),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1263),
.A2(n_1053),
.B(n_1102),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1249),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1241),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1349),
.A2(n_1053),
.B(n_1146),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1199),
.A2(n_1164),
.B(n_1093),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1243),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1350),
.B(n_1304),
.Y(n_1461)
);

AOI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1199),
.A2(n_1093),
.B(n_1005),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1265),
.Y(n_1463)
);

CKINVDCx16_ASAP7_75t_R g1464 ( 
.A(n_1204),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1335),
.B(n_1160),
.C(n_1154),
.Y(n_1465)
);

INVx6_ASAP7_75t_L g1466 ( 
.A(n_1283),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1327),
.A2(n_1251),
.B1(n_1038),
.B2(n_1206),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1224),
.A2(n_521),
.B(n_520),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1265),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1251),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1349),
.A2(n_1146),
.B(n_521),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1300),
.A2(n_1146),
.B(n_647),
.Y(n_1472)
);

OAI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1278),
.A2(n_1122),
.B1(n_404),
.B2(n_407),
.C(n_408),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1280),
.B(n_1154),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1300),
.A2(n_1146),
.B(n_655),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1309),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1258),
.A2(n_1169),
.B1(n_1167),
.B2(n_1137),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1283),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1323),
.B(n_1132),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1269),
.A2(n_416),
.B(n_408),
.C(n_375),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1303),
.A2(n_1146),
.B(n_643),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1261),
.A2(n_1169),
.B1(n_1137),
.B2(n_1122),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1303),
.A2(n_1318),
.B(n_1311),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1289),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1240),
.A2(n_1073),
.B(n_1070),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1204),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1309),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1311),
.A2(n_1146),
.B(n_560),
.Y(n_1488)
);

AOI31xp67_ASAP7_75t_L g1489 ( 
.A1(n_1219),
.A2(n_1223),
.A3(n_1196),
.B(n_1294),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1319),
.B(n_1070),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1247),
.B(n_1093),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1295),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1318),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1255),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1329),
.B(n_349),
.C(n_345),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1236),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1213),
.B(n_1104),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1223),
.A2(n_1122),
.B(n_1005),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1345),
.B(n_1132),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1229),
.A2(n_1132),
.B1(n_1005),
.B2(n_1104),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1319),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1289),
.Y(n_1502)
);

NAND2x1_ASAP7_75t_L g1503 ( 
.A(n_1275),
.B(n_1070),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1224),
.A2(n_560),
.B(n_559),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1325),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1325),
.A2(n_565),
.B(n_386),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1326),
.A2(n_565),
.B(n_386),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1229),
.B(n_1104),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1353),
.B(n_1132),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1326),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1293),
.A2(n_1132),
.B1(n_1104),
.B2(n_413),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_SL g1512 ( 
.A1(n_1237),
.A2(n_396),
.B(n_384),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1338),
.A2(n_1132),
.B1(n_1104),
.B2(n_413),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1246),
.Y(n_1514)
);

AO31x2_ASAP7_75t_L g1515 ( 
.A1(n_1338),
.A2(n_394),
.A3(n_396),
.B(n_397),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1313),
.B(n_1165),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1330),
.A2(n_394),
.B(n_397),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1330),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1331),
.A2(n_1098),
.B(n_1081),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1313),
.B(n_1070),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1331),
.A2(n_1098),
.B(n_1081),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1336),
.A2(n_1073),
.B(n_1098),
.C(n_1081),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1334),
.A2(n_1098),
.B(n_1081),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1246),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1283),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1214),
.A2(n_1158),
.B(n_1098),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1343),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1334),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_R g1529 ( 
.A(n_1343),
.B(n_357),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1337),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1358),
.B(n_1250),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1346),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1346),
.Y(n_1533)
);

AOI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1214),
.A2(n_1073),
.B(n_782),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1351),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1262),
.B(n_359),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1283),
.B(n_668),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1266),
.A2(n_409),
.B1(n_364),
.B2(n_369),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1351),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1352),
.A2(n_232),
.B(n_291),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1407),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1362),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1505),
.A2(n_1237),
.A3(n_1232),
.B(n_1324),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1362),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1456),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1461),
.B(n_1320),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1363),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1409),
.A2(n_1279),
.B1(n_1284),
.B2(n_1317),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1380),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1456),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1450),
.A2(n_1273),
.B(n_1267),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1412),
.Y(n_1552)
);

CKINVDCx11_ASAP7_75t_R g1553 ( 
.A(n_1486),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1534),
.A2(n_1259),
.B(n_1215),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1376),
.Y(n_1555)
);

AND2x6_ASAP7_75t_L g1556 ( 
.A(n_1531),
.B(n_1357),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1380),
.B(n_1197),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1372),
.A2(n_1357),
.B1(n_1197),
.B2(n_350),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1470),
.B(n_1409),
.Y(n_1559)
);

OAI22x1_ASAP7_75t_L g1560 ( 
.A1(n_1441),
.A2(n_1197),
.B1(n_1242),
.B2(n_1244),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1457),
.B(n_1307),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1448),
.A2(n_1305),
.B(n_1259),
.C(n_1356),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1460),
.B(n_1307),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1393),
.Y(n_1564)
);

AND2x2_ASAP7_75t_SL g1565 ( 
.A(n_1450),
.B(n_1513),
.Y(n_1565)
);

OAI222xp33_ASAP7_75t_L g1566 ( 
.A1(n_1473),
.A2(n_440),
.B1(n_438),
.B2(n_435),
.C1(n_433),
.C2(n_430),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1483),
.A2(n_1521),
.B(n_1519),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1366),
.A2(n_413),
.B1(n_302),
.B2(n_350),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1461),
.A2(n_302),
.B1(n_401),
.B2(n_361),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1403),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1373),
.B(n_1307),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1410),
.A2(n_1357),
.B1(n_1283),
.B2(n_1306),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1389),
.A2(n_1238),
.B(n_1306),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1374),
.A2(n_406),
.B1(n_372),
.B2(n_376),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1437),
.A2(n_1357),
.B1(n_379),
.B2(n_380),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1374),
.B(n_1307),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1411),
.B(n_1307),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1483),
.A2(n_1352),
.B(n_1219),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1383),
.A2(n_442),
.B1(n_423),
.B2(n_381),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1377),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1385),
.B(n_1340),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1408),
.B(n_1250),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1424),
.Y(n_1583)
);

BUFx4f_ASAP7_75t_SL g1584 ( 
.A(n_1486),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1418),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1414),
.A2(n_1244),
.B1(n_1242),
.B2(n_1252),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1363),
.B(n_1340),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1385),
.A2(n_1467),
.B1(n_1430),
.B2(n_1451),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1406),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1494),
.B(n_1340),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1389),
.A2(n_1238),
.B(n_1298),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1380),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1430),
.B(n_1340),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1434),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1452),
.A2(n_391),
.B1(n_393),
.B2(n_411),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1494),
.B(n_1340),
.Y(n_1596)
);

BUFx4f_ASAP7_75t_L g1597 ( 
.A(n_1520),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1379),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1413),
.A2(n_412),
.B1(n_414),
.B2(n_415),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1387),
.A2(n_419),
.B1(n_1252),
.B2(n_1328),
.C(n_1250),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1492),
.A2(n_1216),
.B1(n_291),
.B2(n_232),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1379),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1492),
.A2(n_1465),
.B1(n_1428),
.B2(n_1496),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1496),
.A2(n_1288),
.B1(n_1296),
.B2(n_1220),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1508),
.B(n_1296),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1424),
.Y(n_1606)
);

INVx5_ASAP7_75t_L g1607 ( 
.A(n_1434),
.Y(n_1607)
);

O2A1O1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1480),
.A2(n_1288),
.B(n_1296),
.C(n_1275),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1364),
.B(n_1216),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1391),
.B(n_1216),
.Y(n_1610)
);

OAI222xp33_ASAP7_75t_L g1611 ( 
.A1(n_1431),
.A2(n_1420),
.B1(n_1442),
.B2(n_1364),
.C1(n_1538),
.C2(n_1536),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1389),
.A2(n_1301),
.B(n_1226),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1502),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1511),
.A2(n_1220),
.B1(n_1348),
.B2(n_1256),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1522),
.A2(n_1225),
.B(n_1220),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1508),
.B(n_232),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1495),
.B(n_1256),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1447),
.B(n_1315),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1398),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1380),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1390),
.A2(n_1491),
.B1(n_1396),
.B2(n_1447),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1491),
.B(n_1257),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1436),
.A2(n_1215),
.B1(n_1315),
.B2(n_1348),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1386),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1497),
.B(n_1257),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1514),
.B(n_1332),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1464),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1432),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1440),
.B(n_1354),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1500),
.A2(n_1348),
.B1(n_1355),
.B2(n_1316),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1390),
.A2(n_291),
.B1(n_1245),
.B2(n_19),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_R g1632 ( 
.A(n_1400),
.B(n_1314),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1497),
.B(n_12),
.Y(n_1633)
);

CKINVDCx11_ASAP7_75t_R g1634 ( 
.A(n_1436),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1404),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1432),
.Y(n_1636)
);

AND2x6_ASAP7_75t_SL g1637 ( 
.A(n_1474),
.B(n_16),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1400),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1484),
.B(n_20),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1527),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1479),
.A2(n_668),
.B(n_291),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1519),
.A2(n_291),
.B(n_668),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1417),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1397),
.B(n_291),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1425),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1388),
.B(n_21),
.Y(n_1646)
);

INVx4_ASAP7_75t_L g1647 ( 
.A(n_1398),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1524),
.B(n_21),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1398),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1527),
.Y(n_1650)
);

O2A1O1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1423),
.A2(n_22),
.B(n_25),
.C(n_26),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1388),
.B(n_22),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1390),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1499),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1404),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1463),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1444),
.A2(n_782),
.B1(n_768),
.B2(n_668),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1394),
.A2(n_782),
.B1(n_768),
.B2(n_668),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1469),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1396),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_1660)
);

AO31x2_ASAP7_75t_L g1661 ( 
.A1(n_1505),
.A2(n_38),
.A3(n_39),
.B(n_41),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1394),
.B(n_39),
.Y(n_1662)
);

BUFx4f_ASAP7_75t_SL g1663 ( 
.A(n_1520),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1521),
.A2(n_782),
.B(n_768),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1416),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1447),
.B(n_44),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1516),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1520),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1400),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1498),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.C(n_49),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1435),
.Y(n_1671)
);

OAI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1509),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.C(n_52),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1443),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1396),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1674)
);

AOI21xp33_ASAP7_75t_L g1675 ( 
.A1(n_1498),
.A2(n_56),
.B(n_58),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1405),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.C(n_69),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1523),
.A2(n_219),
.B(n_213),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1515),
.B(n_1435),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1392),
.A2(n_61),
.B1(n_70),
.B2(n_72),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1515),
.B(n_73),
.Y(n_1680)
);

CKINVDCx16_ASAP7_75t_R g1681 ( 
.A(n_1400),
.Y(n_1681)
);

AO31x2_ASAP7_75t_L g1682 ( 
.A1(n_1510),
.A2(n_74),
.A3(n_75),
.B(n_77),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1416),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1523),
.A2(n_210),
.B(n_200),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1440),
.B(n_195),
.Y(n_1685)
);

BUFx4f_ASAP7_75t_L g1686 ( 
.A(n_1434),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1485),
.A2(n_181),
.B(n_180),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1434),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1490),
.A2(n_175),
.B(n_173),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1529),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1433),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1398),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1446),
.B(n_77),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1531),
.A2(n_79),
.B(n_81),
.C(n_82),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1433),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1439),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1466),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1439),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1476),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1429),
.A2(n_81),
.B(n_82),
.Y(n_1700)
);

CKINVDCx14_ASAP7_75t_R g1701 ( 
.A(n_1384),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1466),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1515),
.B(n_86),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1476),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1482),
.B(n_87),
.C(n_88),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1487),
.Y(n_1706)
);

BUFx8_ASAP7_75t_L g1707 ( 
.A(n_1434),
.Y(n_1707)
);

AO31x2_ASAP7_75t_L g1708 ( 
.A1(n_1510),
.A2(n_1533),
.A3(n_1535),
.B(n_1539),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1487),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1392),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1477),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1382),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1440),
.B(n_168),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_SL g1714 ( 
.A1(n_1395),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1501),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_SL g1716 ( 
.A(n_1503),
.B(n_94),
.C(n_96),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1490),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1392),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1515),
.B(n_97),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1405),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_1720)
);

BUFx4f_ASAP7_75t_L g1721 ( 
.A(n_1453),
.Y(n_1721)
);

BUFx4f_ASAP7_75t_SL g1722 ( 
.A(n_1453),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1515),
.B(n_1449),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1382),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1401),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1453),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1399),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1401),
.A2(n_108),
.B1(n_167),
.B2(n_111),
.Y(n_1728)
);

BUFx12f_ASAP7_75t_L g1729 ( 
.A(n_1453),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1440),
.B(n_127),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1570),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1667),
.A2(n_1512),
.B1(n_1535),
.B2(n_1533),
.C(n_1532),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1544),
.Y(n_1733)
);

OAI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1568),
.A2(n_1462),
.B(n_1459),
.C(n_1449),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1544),
.Y(n_1735)
);

AOI222xp33_ASAP7_75t_L g1736 ( 
.A1(n_1568),
.A2(n_1512),
.B1(n_108),
.B2(n_1528),
.C1(n_1530),
.C2(n_1518),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1672),
.A2(n_1449),
.B1(n_1370),
.B2(n_1493),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1569),
.A2(n_1490),
.B1(n_1466),
.B2(n_1440),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1569),
.A2(n_1466),
.B1(n_1445),
.B2(n_1395),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1578),
.A2(n_1402),
.B(n_1422),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1585),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1559),
.B(n_1370),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1581),
.B(n_1577),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1653),
.A2(n_1370),
.B1(n_1493),
.B2(n_1518),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1673),
.A2(n_1478),
.B1(n_1453),
.B2(n_1525),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1574),
.A2(n_1503),
.B1(n_1462),
.B2(n_1445),
.C(n_1459),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1653),
.A2(n_1660),
.B1(n_1674),
.B2(n_1670),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1660),
.A2(n_1526),
.B1(n_1429),
.B2(n_1438),
.Y(n_1748)
);

AOI22x1_ASAP7_75t_L g1749 ( 
.A1(n_1560),
.A2(n_1525),
.B1(n_1445),
.B2(n_1478),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1668),
.B(n_1369),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1583),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1551),
.A2(n_1526),
.B(n_1525),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1576),
.B(n_1455),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1589),
.B(n_1369),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1729),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_SL g1756 ( 
.A1(n_1565),
.A2(n_1478),
.B1(n_1369),
.B2(n_1526),
.Y(n_1756)
);

CKINVDCx6p67_ASAP7_75t_R g1757 ( 
.A(n_1553),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_L g1758 ( 
.A(n_1651),
.B(n_1504),
.C(n_1468),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1611),
.B(n_1478),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_SL g1760 ( 
.A1(n_1565),
.A2(n_1478),
.B1(n_1438),
.B2(n_1488),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1729),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1595),
.A2(n_1546),
.B1(n_1575),
.B2(n_1582),
.Y(n_1762)
);

OAI211xp5_ASAP7_75t_L g1763 ( 
.A1(n_1715),
.A2(n_1540),
.B(n_1504),
.C(n_1534),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1616),
.B(n_1455),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1566),
.A2(n_1489),
.B1(n_1537),
.B2(n_1488),
.C(n_1507),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1674),
.A2(n_1415),
.B1(n_1419),
.B2(n_1399),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1595),
.A2(n_1458),
.B1(n_1481),
.B2(n_1472),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1711),
.A2(n_1504),
.B1(n_1468),
.B2(n_1489),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1705),
.A2(n_1540),
.B1(n_1458),
.B2(n_1472),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1679),
.A2(n_1415),
.B1(n_1419),
.B2(n_1475),
.Y(n_1770)
);

OAI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1694),
.A2(n_1468),
.B(n_1517),
.C(n_1507),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1593),
.B(n_1605),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1679),
.A2(n_1381),
.B1(n_1506),
.B2(n_1517),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1600),
.A2(n_1402),
.B(n_1471),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1603),
.B(n_1454),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1597),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1717),
.A2(n_1537),
.B1(n_1506),
.B2(n_1381),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1704),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1599),
.A2(n_1537),
.B1(n_1421),
.B2(n_1426),
.Y(n_1779)
);

INVx6_ASAP7_75t_L g1780 ( 
.A(n_1707),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1553),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1547),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1599),
.A2(n_1426),
.B1(n_1421),
.B2(n_1361),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1562),
.A2(n_1427),
.B(n_1454),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1708),
.Y(n_1785)
);

BUFx10_ASAP7_75t_L g1786 ( 
.A(n_1542),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1654),
.A2(n_1427),
.B1(n_1361),
.B2(n_1365),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1583),
.Y(n_1788)
);

BUFx8_ASAP7_75t_SL g1789 ( 
.A(n_1545),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1700),
.A2(n_1422),
.B1(n_1378),
.B2(n_1375),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1597),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1588),
.A2(n_1603),
.B1(n_1574),
.B2(n_1579),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1606),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1562),
.A2(n_1367),
.B(n_1378),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1588),
.A2(n_1375),
.B1(n_1371),
.B2(n_1368),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1541),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1694),
.A2(n_1631),
.B(n_1728),
.C(n_1725),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1609),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1654),
.A2(n_1368),
.B1(n_1365),
.B2(n_1371),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1628),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1633),
.B(n_1666),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1636),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1725),
.A2(n_110),
.B1(n_124),
.B2(n_134),
.C(n_148),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1675),
.A2(n_151),
.B1(n_152),
.B2(n_1631),
.C(n_1676),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1714),
.A2(n_1716),
.B1(n_1720),
.B2(n_1728),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1648),
.B(n_1668),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1720),
.A2(n_1634),
.B1(n_1680),
.B2(n_1703),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1693),
.B(n_1610),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1671),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1650),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1634),
.A2(n_1558),
.B1(n_1582),
.B2(n_1719),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1610),
.B(n_1613),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1548),
.A2(n_1644),
.B1(n_1639),
.B2(n_1621),
.C(n_1662),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1643),
.Y(n_1814)
);

AOI222xp33_ASAP7_75t_L g1815 ( 
.A1(n_1584),
.A2(n_1644),
.B1(n_1548),
.B2(n_1690),
.C1(n_1571),
.C2(n_1552),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1697),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1545),
.A2(n_1624),
.B1(n_1627),
.B2(n_1617),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1591),
.A2(n_1573),
.B(n_1615),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1555),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1645),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1681),
.A2(n_1584),
.B1(n_1556),
.B2(n_1730),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1572),
.A2(n_1621),
.B1(n_1606),
.B2(n_1640),
.Y(n_1822)
);

AOI21xp33_ASAP7_75t_L g1823 ( 
.A1(n_1617),
.A2(n_1626),
.B(n_1563),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1564),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1646),
.A2(n_1652),
.B1(n_1587),
.B2(n_1561),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1590),
.B(n_1596),
.Y(n_1826)
);

BUFx5_ASAP7_75t_L g1827 ( 
.A(n_1724),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1641),
.A2(n_1689),
.B1(n_1687),
.B2(n_1601),
.C(n_1626),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1556),
.A2(n_1730),
.B1(n_1713),
.B2(n_1685),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1625),
.B(n_1622),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1691),
.B(n_1695),
.Y(n_1831)
);

BUFx4f_ASAP7_75t_SL g1832 ( 
.A(n_1640),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1701),
.A2(n_1556),
.B1(n_1659),
.B2(n_1656),
.Y(n_1833)
);

OAI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1663),
.A2(n_1632),
.B1(n_1557),
.B2(n_1637),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1701),
.A2(n_1556),
.B1(n_1601),
.B2(n_1730),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1702),
.A2(n_1663),
.B1(n_1721),
.B2(n_1686),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1618),
.B(n_1586),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1618),
.B(n_1697),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1612),
.A2(n_1567),
.B(n_1664),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1618),
.B(n_1592),
.Y(n_1840)
);

INVx4_ASAP7_75t_L g1841 ( 
.A(n_1722),
.Y(n_1841)
);

OAI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1632),
.A2(n_1557),
.B1(n_1722),
.B2(n_1638),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1604),
.A2(n_1630),
.B(n_1623),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1550),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1686),
.Y(n_1845)
);

AO221x1_ASAP7_75t_L g1846 ( 
.A1(n_1623),
.A2(n_1604),
.B1(n_1657),
.B2(n_1638),
.C(n_1549),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1554),
.A2(n_1642),
.B(n_1677),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1696),
.B(n_1709),
.Y(n_1848)
);

INVxp33_ASAP7_75t_L g1849 ( 
.A(n_1594),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1685),
.B(n_1713),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1698),
.B(n_1699),
.Y(n_1851)
);

NAND2x1_ASAP7_75t_L g1852 ( 
.A(n_1557),
.B(n_1669),
.Y(n_1852)
);

BUFx12f_ASAP7_75t_L g1853 ( 
.A(n_1707),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1608),
.A2(n_1614),
.B(n_1713),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1692),
.B(n_1706),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1629),
.A2(n_1592),
.B1(n_1549),
.B2(n_1669),
.C(n_1620),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1556),
.A2(n_1685),
.B1(n_1678),
.B2(n_1620),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1580),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1598),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1594),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1707),
.A2(n_1607),
.B1(n_1721),
.B2(n_1619),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1598),
.A2(n_1655),
.B1(n_1665),
.B2(n_1602),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1602),
.A2(n_1665),
.B1(n_1655),
.B2(n_1683),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1594),
.Y(n_1864)
);

OAI211xp5_ASAP7_75t_L g1865 ( 
.A1(n_1710),
.A2(n_1718),
.B(n_1723),
.C(n_1635),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1619),
.B(n_1647),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1635),
.A2(n_1683),
.B1(n_1712),
.B2(n_1727),
.C(n_1658),
.Y(n_1867)
);

OAI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1607),
.A2(n_1649),
.B1(n_1647),
.B2(n_1629),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1661),
.B(n_1682),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1649),
.A2(n_1607),
.B1(n_1594),
.B2(n_1726),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1688),
.A2(n_1726),
.B1(n_1607),
.B2(n_1684),
.Y(n_1871)
);

AOI21xp33_ASAP7_75t_L g1872 ( 
.A1(n_1712),
.A2(n_1727),
.B(n_1688),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1726),
.A2(n_1688),
.B1(n_1661),
.B2(n_1682),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1688),
.A2(n_1726),
.B1(n_1661),
.B2(n_1682),
.C(n_1543),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1661),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1875)
);

INVx4_ASAP7_75t_L g1876 ( 
.A(n_1682),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1543),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1543),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1543),
.A2(n_825),
.B1(n_670),
.B2(n_1015),
.C(n_1667),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1673),
.A2(n_1015),
.B1(n_1002),
.B2(n_1117),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1589),
.B(n_1015),
.Y(n_1882)
);

OAI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1667),
.A2(n_1117),
.B1(n_1715),
.B2(n_1672),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1576),
.B(n_1616),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1570),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1886)
);

INVx4_ASAP7_75t_L g1887 ( 
.A(n_1722),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1589),
.B(n_1015),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1889)
);

INVx4_ASAP7_75t_L g1890 ( 
.A(n_1722),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1568),
.A2(n_1015),
.B1(n_1117),
.B2(n_1049),
.Y(n_1894)
);

INVx5_ASAP7_75t_L g1895 ( 
.A(n_1557),
.Y(n_1895)
);

AOI222xp33_ASAP7_75t_L g1896 ( 
.A1(n_1667),
.A2(n_587),
.B1(n_830),
.B2(n_1015),
.C1(n_976),
.C2(n_1043),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1570),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_R g1898 ( 
.A(n_1702),
.B(n_1292),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1667),
.A2(n_1015),
.B1(n_1260),
.B2(n_976),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1589),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1570),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1570),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1826),
.B(n_1798),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1895),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1742),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1743),
.B(n_1830),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1792),
.A2(n_1892),
.B1(n_1893),
.B2(n_1891),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1808),
.B(n_1812),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1895),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1753),
.B(n_1878),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1882),
.B(n_1888),
.Y(n_1911)
);

AND2x2_ASAP7_75t_SL g1912 ( 
.A(n_1747),
.B(n_1805),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1894),
.A2(n_1803),
.B1(n_1759),
.B2(n_1846),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1772),
.B(n_1884),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1751),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1785),
.Y(n_1916)
);

INVx2_ASAP7_75t_SL g1917 ( 
.A(n_1895),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1800),
.B(n_1876),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1800),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1825),
.B(n_1823),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1827),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1876),
.B(n_1731),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1877),
.B(n_1827),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1827),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1809),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1809),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1883),
.A2(n_1747),
.B1(n_1889),
.B2(n_1891),
.C(n_1899),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1827),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1869),
.B(n_1764),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1877),
.B(n_1827),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1827),
.B(n_1874),
.Y(n_1931)
);

AOI21xp33_ASAP7_75t_L g1932 ( 
.A1(n_1879),
.A2(n_1896),
.B(n_1815),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1831),
.B(n_1825),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1852),
.Y(n_1934)
);

NAND3xp33_ASAP7_75t_L g1935 ( 
.A(n_1880),
.B(n_1889),
.C(n_1886),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1741),
.Y(n_1936)
);

NAND2x1_ASAP7_75t_L g1937 ( 
.A(n_1780),
.B(n_1871),
.Y(n_1937)
);

INVx3_ASAP7_75t_L g1938 ( 
.A(n_1839),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1802),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1885),
.Y(n_1940)
);

INVx4_ASAP7_75t_L g1941 ( 
.A(n_1895),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1897),
.B(n_1901),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1859),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1902),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1782),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1840),
.B(n_1843),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1740),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1814),
.B(n_1820),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1824),
.B(n_1775),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1796),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1840),
.B(n_1819),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1740),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1854),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1880),
.A2(n_1899),
.B1(n_1893),
.B2(n_1892),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1775),
.B(n_1740),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1865),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1900),
.B(n_1778),
.Y(n_1957)
);

AND2x6_ASAP7_75t_L g1958 ( 
.A(n_1776),
.B(n_1791),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1856),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_L g1960 ( 
.A(n_1868),
.B(n_1834),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1873),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1873),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1851),
.Y(n_1963)
);

AO21x2_ASAP7_75t_L g1964 ( 
.A1(n_1818),
.A2(n_1794),
.B(n_1774),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1844),
.B(n_1789),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1886),
.A2(n_1807),
.B1(n_1883),
.B2(n_1811),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1857),
.B(n_1850),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1847),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1801),
.B(n_1756),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1858),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1848),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1857),
.B(n_1837),
.Y(n_1972)
);

NOR2x1_ASAP7_75t_SL g1973 ( 
.A(n_1850),
.B(n_1734),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1862),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1864),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1837),
.B(n_1855),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1862),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1807),
.A2(n_1811),
.B1(n_1881),
.B2(n_1805),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1860),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1787),
.B(n_1799),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1838),
.B(n_1744),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1822),
.B(n_1795),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1749),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1863),
.Y(n_1985)
);

OAI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1797),
.A2(n_1804),
.B1(n_1875),
.B2(n_1762),
.C(n_1813),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1783),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1752),
.B(n_1767),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1737),
.B(n_1833),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1744),
.B(n_1748),
.Y(n_1990)
);

CKINVDCx10_ASAP7_75t_R g1991 ( 
.A(n_1757),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1748),
.B(n_1863),
.Y(n_1992)
);

NAND2xp33_ASAP7_75t_R g1993 ( 
.A(n_1733),
.B(n_1735),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1746),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1784),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1787),
.B(n_1799),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1832),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1872),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1768),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1816),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1768),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1864),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1758),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1790),
.B(n_1760),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1771),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1875),
.B(n_1797),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1934),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1915),
.B(n_1793),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1912),
.A2(n_1736),
.B1(n_1834),
.B2(n_1759),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1912),
.A2(n_1828),
.B1(n_1745),
.B2(n_1835),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1939),
.Y(n_2011)
);

OAI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1979),
.A2(n_1817),
.B1(n_1833),
.B2(n_1821),
.C(n_1829),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1912),
.A2(n_1835),
.B1(n_1842),
.B2(n_1732),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1910),
.B(n_1806),
.Y(n_2014)
);

OAI21x1_ASAP7_75t_L g2015 ( 
.A1(n_1938),
.A2(n_1779),
.B(n_1773),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1939),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1953),
.B(n_1898),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1971),
.B(n_1842),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_R g2019 ( 
.A(n_1993),
.B(n_1781),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1943),
.Y(n_2020)
);

OAI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1935),
.A2(n_1832),
.B1(n_1738),
.B2(n_1739),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1939),
.Y(n_2022)
);

AOI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_1932),
.A2(n_1737),
.B1(n_1777),
.B2(n_1868),
.C(n_1763),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1986),
.A2(n_1791),
.B1(n_1776),
.B2(n_1816),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1940),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1986),
.A2(n_1791),
.B1(n_1776),
.B2(n_1750),
.Y(n_2026)
);

NAND2xp33_ASAP7_75t_R g2027 ( 
.A(n_1953),
.B(n_1898),
.Y(n_2027)
);

NOR5xp2_ASAP7_75t_SL g2028 ( 
.A(n_1932),
.B(n_1870),
.C(n_1765),
.D(n_1836),
.E(n_1867),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1971),
.B(n_1788),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1977),
.B(n_1866),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_1935),
.A2(n_1777),
.B1(n_1770),
.B2(n_1773),
.C(n_1766),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1910),
.B(n_1766),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_R g2033 ( 
.A1(n_1967),
.A2(n_1750),
.B(n_1853),
.Y(n_2033)
);

INVxp67_ASAP7_75t_SL g2034 ( 
.A(n_1956),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1943),
.Y(n_2035)
);

AOI33xp33_ASAP7_75t_L g2036 ( 
.A1(n_1907),
.A2(n_1769),
.A3(n_1770),
.B1(n_1861),
.B2(n_1786),
.B3(n_1849),
.Y(n_2036)
);

NAND2xp33_ASAP7_75t_R g2037 ( 
.A(n_1965),
.B(n_1755),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1905),
.B(n_1755),
.Y(n_2038)
);

OAI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_1966),
.A2(n_1890),
.B(n_1887),
.C(n_1841),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1959),
.B(n_1791),
.Y(n_2040)
);

INVxp67_ASAP7_75t_SL g2041 ( 
.A(n_1956),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1954),
.A2(n_1927),
.B1(n_1913),
.B2(n_2006),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_1915),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_SL g2044 ( 
.A1(n_1913),
.A2(n_1780),
.B1(n_1890),
.B2(n_1841),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1910),
.B(n_1761),
.Y(n_2045)
);

OAI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_1927),
.A2(n_1761),
.B1(n_1887),
.B2(n_1780),
.C(n_1776),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1940),
.Y(n_2047)
);

AOI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_2006),
.A2(n_1920),
.B1(n_1961),
.B2(n_2005),
.C(n_1911),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1960),
.A2(n_1786),
.B1(n_1845),
.B2(n_1959),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1940),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1919),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1960),
.A2(n_1845),
.B1(n_1959),
.B2(n_1920),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1949),
.B(n_1845),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1938),
.A2(n_1845),
.B(n_1947),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1997),
.Y(n_2055)
);

AO21x2_ASAP7_75t_L g2056 ( 
.A1(n_1964),
.A2(n_1995),
.B(n_2003),
.Y(n_2056)
);

OAI211xp5_ASAP7_75t_SL g2057 ( 
.A1(n_1945),
.A2(n_2005),
.B(n_1977),
.C(n_1983),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1947),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1936),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1964),
.A2(n_1988),
.B(n_1973),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_SL g2061 ( 
.A1(n_1997),
.A2(n_1937),
.B1(n_1961),
.B2(n_1983),
.Y(n_2061)
);

OAI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1989),
.A2(n_1994),
.B1(n_1937),
.B2(n_1933),
.Y(n_2062)
);

INVx5_ASAP7_75t_L g2063 ( 
.A(n_1938),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_1906),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1919),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2003),
.A2(n_1994),
.B(n_2001),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_SL g2067 ( 
.A1(n_2004),
.A2(n_1973),
.B1(n_1981),
.B2(n_1996),
.Y(n_2067)
);

OAI33xp33_ASAP7_75t_L g2068 ( 
.A1(n_1945),
.A2(n_1933),
.A3(n_1962),
.B1(n_1957),
.B2(n_1908),
.B3(n_2001),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_1905),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1947),
.Y(n_2070)
);

OAI31xp33_ASAP7_75t_L g2071 ( 
.A1(n_1994),
.A2(n_1981),
.A3(n_1996),
.B(n_1989),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1925),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1936),
.Y(n_2073)
);

AOI211xp5_ASAP7_75t_SL g2074 ( 
.A1(n_1981),
.A2(n_1996),
.B(n_2004),
.C(n_1962),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_L g2075 ( 
.A(n_2003),
.B(n_1999),
.C(n_1995),
.Y(n_2075)
);

OAI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1997),
.A2(n_1984),
.B1(n_1908),
.B2(n_1972),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_1915),
.B(n_1918),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_1949),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1903),
.B(n_1906),
.Y(n_2079)
);

NOR3xp33_ASAP7_75t_L g2080 ( 
.A(n_1999),
.B(n_1984),
.C(n_2004),
.Y(n_2080)
);

OAI31xp33_ASAP7_75t_L g2081 ( 
.A1(n_1990),
.A2(n_1988),
.A3(n_1972),
.B(n_1992),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_SL g2082 ( 
.A1(n_1967),
.A2(n_1990),
.B(n_1992),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_1929),
.B(n_1903),
.Y(n_2083)
);

AOI222xp33_ASAP7_75t_L g2084 ( 
.A1(n_1969),
.A2(n_1967),
.B1(n_1985),
.B2(n_1974),
.C1(n_1978),
.C2(n_1988),
.Y(n_2084)
);

OAI321xp33_ASAP7_75t_L g2085 ( 
.A1(n_1984),
.A2(n_1985),
.A3(n_1978),
.B1(n_1974),
.B2(n_1987),
.C(n_1998),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1925),
.Y(n_2086)
);

NOR2x1_ASAP7_75t_L g2087 ( 
.A(n_2002),
.B(n_1957),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1952),
.Y(n_2088)
);

AOI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_1969),
.A2(n_1949),
.B1(n_1931),
.B2(n_1987),
.C(n_1988),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1967),
.A2(n_1946),
.B1(n_1976),
.B2(n_1951),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1926),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2064),
.B(n_1931),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_2043),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2011),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2011),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2022),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2083),
.B(n_1929),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_2079),
.B(n_1991),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2078),
.B(n_1931),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2083),
.B(n_1998),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_2071),
.B(n_1934),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2069),
.B(n_1987),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2007),
.B(n_1904),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2022),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2077),
.B(n_1930),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2077),
.B(n_1930),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2025),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2077),
.B(n_1930),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2032),
.B(n_1923),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2020),
.B(n_1944),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2032),
.B(n_1923),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2043),
.B(n_1923),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2045),
.B(n_1955),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_2063),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2025),
.Y(n_2115)
);

BUFx2_ASAP7_75t_L g2116 ( 
.A(n_2087),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_2035),
.B(n_1955),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2047),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2047),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2034),
.B(n_1944),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2045),
.B(n_1955),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2016),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2016),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_2041),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2007),
.B(n_1904),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2050),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2050),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2014),
.B(n_1928),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2014),
.B(n_1928),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2051),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2051),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2065),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2075),
.B(n_1944),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2065),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2072),
.B(n_1948),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2072),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2086),
.B(n_1948),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_2038),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2086),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_2058),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_2063),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_2063),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_2030),
.B(n_1991),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2091),
.B(n_1948),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2070),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_2063),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2091),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2053),
.B(n_1924),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2038),
.B(n_1916),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2070),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2059),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_2007),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2088),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2053),
.B(n_1924),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2089),
.B(n_2073),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2090),
.B(n_1924),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2060),
.B(n_2082),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2054),
.B(n_1904),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2074),
.B(n_1921),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2088),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2018),
.B(n_1942),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2140),
.Y(n_2162)
);

OAI21xp33_ASAP7_75t_SL g2163 ( 
.A1(n_2101),
.A2(n_2036),
.B(n_2081),
.Y(n_2163)
);

AOI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_2157),
.A2(n_2048),
.B1(n_2042),
.B2(n_2080),
.C(n_2076),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2100),
.B(n_2029),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2130),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2140),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_SL g2168 ( 
.A(n_2157),
.B(n_2062),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2109),
.B(n_2008),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2109),
.B(n_2008),
.Y(n_2170)
);

O2A1O1Ixp33_ASAP7_75t_L g2171 ( 
.A1(n_2155),
.A2(n_2021),
.B(n_2057),
.C(n_2012),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2161),
.B(n_2084),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2100),
.B(n_2056),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_2133),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2140),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2117),
.B(n_2056),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2111),
.B(n_2008),
.Y(n_2177)
);

AOI22xp33_ASAP7_75t_L g2178 ( 
.A1(n_2159),
.A2(n_2044),
.B1(n_2067),
.B2(n_2009),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2140),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2161),
.B(n_2066),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2111),
.B(n_2055),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2093),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2130),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2098),
.B(n_2055),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2131),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2155),
.B(n_1976),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2099),
.B(n_2054),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2131),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2132),
.Y(n_2189)
);

NAND2x2_ASAP7_75t_L g2190 ( 
.A(n_2114),
.B(n_2033),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2117),
.B(n_2056),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2099),
.B(n_2063),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2097),
.B(n_1970),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2132),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2105),
.B(n_1982),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2092),
.B(n_1914),
.Y(n_2196)
);

AOI32xp33_ASAP7_75t_L g2197 ( 
.A1(n_2159),
.A2(n_2052),
.A3(n_2017),
.B1(n_2010),
.B2(n_2013),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2105),
.B(n_2106),
.Y(n_2198)
);

INVx2_ASAP7_75t_SL g2199 ( 
.A(n_2152),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2106),
.B(n_1982),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2134),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2092),
.B(n_1914),
.Y(n_2202)
);

NOR2x1p5_ASAP7_75t_L g2203 ( 
.A(n_2133),
.B(n_1934),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2124),
.B(n_2023),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2108),
.B(n_1951),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2114),
.B(n_1934),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_2114),
.B(n_1934),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2108),
.B(n_1951),
.Y(n_2208)
);

AOI222xp33_ASAP7_75t_L g2209 ( 
.A1(n_2143),
.A2(n_2031),
.B1(n_2068),
.B2(n_2061),
.C1(n_2039),
.C2(n_2085),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2112),
.B(n_1951),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2112),
.B(n_2015),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_2141),
.B(n_1934),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2134),
.Y(n_2213)
);

OR2x6_ASAP7_75t_L g2214 ( 
.A(n_2141),
.B(n_2015),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2097),
.B(n_1970),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2136),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2150),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2166),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2166),
.Y(n_2219)
);

NAND3xp33_ASAP7_75t_L g2220 ( 
.A(n_2163),
.B(n_2036),
.C(n_2049),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2198),
.B(n_2116),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2163),
.B(n_2019),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_2171),
.A2(n_2017),
.B(n_2040),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2183),
.Y(n_2224)
);

NAND2x1_ASAP7_75t_L g2225 ( 
.A(n_2206),
.B(n_2116),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2183),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2174),
.B(n_2102),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2198),
.B(n_2138),
.Y(n_2228)
);

NAND4xp25_ASAP7_75t_L g2229 ( 
.A(n_2209),
.B(n_2164),
.C(n_2178),
.D(n_2204),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2184),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2180),
.B(n_2186),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2209),
.B(n_2124),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2162),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2168),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2172),
.B(n_2138),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2165),
.B(n_2102),
.Y(n_2236)
);

OAI21xp33_ASAP7_75t_SL g2237 ( 
.A1(n_2203),
.A2(n_2146),
.B(n_2142),
.Y(n_2237)
);

AND2x2_ASAP7_75t_SL g2238 ( 
.A(n_2206),
.B(n_2207),
.Y(n_2238)
);

OR2x4_ASAP7_75t_L g2239 ( 
.A(n_2165),
.B(n_2120),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2162),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2196),
.B(n_2120),
.Y(n_2241)
);

NOR2xp67_ASAP7_75t_L g2242 ( 
.A(n_2199),
.B(n_2141),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2195),
.B(n_2128),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2202),
.B(n_2046),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2203),
.B(n_2142),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2192),
.B(n_2148),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2162),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2182),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2182),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2185),
.Y(n_2250)
);

AOI21xp33_ASAP7_75t_SL g2251 ( 
.A1(n_2197),
.A2(n_2037),
.B(n_2027),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2185),
.Y(n_2252)
);

OA21x2_ASAP7_75t_L g2253 ( 
.A1(n_2217),
.A2(n_2142),
.B(n_2146),
.Y(n_2253)
);

NOR2x1_ASAP7_75t_L g2254 ( 
.A(n_2206),
.B(n_2152),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2188),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2192),
.B(n_2148),
.Y(n_2256)
);

NAND2xp33_ASAP7_75t_R g2257 ( 
.A(n_2206),
.B(n_2028),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2188),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2189),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2195),
.B(n_2128),
.Y(n_2260)
);

INVxp67_ASAP7_75t_L g2261 ( 
.A(n_2181),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2189),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2194),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2200),
.B(n_2129),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2167),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2167),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2194),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2201),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2201),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2213),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2213),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2181),
.B(n_2110),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2238),
.Y(n_2273)
);

OAI211xp5_ASAP7_75t_SL g2274 ( 
.A1(n_2232),
.A2(n_2197),
.B(n_2173),
.C(n_2026),
.Y(n_2274)
);

O2A1O1Ixp33_ASAP7_75t_SL g2275 ( 
.A1(n_2222),
.A2(n_2093),
.B(n_2199),
.C(n_2146),
.Y(n_2275)
);

OAI31xp33_ASAP7_75t_L g2276 ( 
.A1(n_2229),
.A2(n_2207),
.A3(n_2212),
.B(n_2211),
.Y(n_2276)
);

OAI332xp33_ASAP7_75t_L g2277 ( 
.A1(n_2235),
.A2(n_2173),
.A3(n_2191),
.B1(n_2176),
.B2(n_2110),
.B3(n_2216),
.C1(n_2217),
.C2(n_2149),
.Y(n_2277)
);

AOI31xp33_ASAP7_75t_L g2278 ( 
.A1(n_2220),
.A2(n_2024),
.A3(n_2207),
.B(n_2212),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2238),
.B(n_2200),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2246),
.B(n_2169),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_L g2281 ( 
.A(n_2251),
.B(n_2214),
.C(n_2211),
.Y(n_2281)
);

OAI21xp33_ASAP7_75t_L g2282 ( 
.A1(n_2234),
.A2(n_2214),
.B(n_2187),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2225),
.Y(n_2283)
);

AOI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2257),
.A2(n_2190),
.B1(n_1946),
.B2(n_2212),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_2225),
.Y(n_2285)
);

OAI22xp5_ASAP7_75t_L g2286 ( 
.A1(n_2249),
.A2(n_2190),
.B1(n_2214),
.B2(n_1946),
.Y(n_2286)
);

NOR2x1_ASAP7_75t_L g2287 ( 
.A(n_2254),
.B(n_2207),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2244),
.A2(n_2190),
.B1(n_1946),
.B2(n_2212),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2231),
.B(n_2248),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2255),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2243),
.B(n_2193),
.Y(n_2291)
);

AOI222xp33_ASAP7_75t_L g2292 ( 
.A1(n_2249),
.A2(n_2028),
.B1(n_1963),
.B2(n_2216),
.C1(n_2187),
.C2(n_1950),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2218),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_L g2294 ( 
.A1(n_2230),
.A2(n_1963),
.B1(n_1950),
.B2(n_2151),
.C1(n_1970),
.C2(n_2156),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2218),
.Y(n_2295)
);

AOI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_2261),
.A2(n_2214),
.B1(n_2156),
.B2(n_1964),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2223),
.B(n_2241),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2219),
.B(n_2151),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2230),
.A2(n_2214),
.B(n_2158),
.Y(n_2299)
);

INVxp67_ASAP7_75t_L g2300 ( 
.A(n_2272),
.Y(n_2300)
);

OR2x6_ASAP7_75t_L g2301 ( 
.A(n_2242),
.B(n_1941),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2224),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2260),
.B(n_2193),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2228),
.B(n_2169),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2246),
.B(n_2170),
.Y(n_2305)
);

O2A1O1Ixp33_ASAP7_75t_L g2306 ( 
.A1(n_2237),
.A2(n_2176),
.B(n_2191),
.C(n_1964),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2271),
.Y(n_2307)
);

OR2x2_ASAP7_75t_L g2308 ( 
.A(n_2264),
.B(n_2215),
.Y(n_2308)
);

NOR2x1_ASAP7_75t_SL g2309 ( 
.A(n_2227),
.B(n_2170),
.Y(n_2309)
);

AOI211xp5_ASAP7_75t_L g2310 ( 
.A1(n_2245),
.A2(n_2158),
.B(n_2215),
.C(n_2103),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2256),
.B(n_2177),
.Y(n_2311)
);

AOI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_2245),
.A2(n_1958),
.B1(n_2177),
.B2(n_2158),
.Y(n_2312)
);

NAND2x1_ASAP7_75t_SL g2313 ( 
.A(n_2245),
.B(n_2158),
.Y(n_2313)
);

INVxp67_ASAP7_75t_L g2314 ( 
.A(n_2221),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2236),
.B(n_2149),
.Y(n_2315)
);

AOI221xp5_ASAP7_75t_L g2316 ( 
.A1(n_2277),
.A2(n_2267),
.B1(n_2250),
.B2(n_2269),
.C(n_2268),
.Y(n_2316)
);

OA22x2_ASAP7_75t_L g2317 ( 
.A1(n_2297),
.A2(n_2221),
.B1(n_2252),
.B2(n_2258),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2300),
.B(n_2228),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2314),
.B(n_2256),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2273),
.B(n_2239),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2293),
.Y(n_2321)
);

O2A1O1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2274),
.A2(n_2227),
.B(n_2270),
.C(n_2224),
.Y(n_2322)
);

NAND4xp25_ASAP7_75t_L g2323 ( 
.A(n_2276),
.B(n_2271),
.C(n_2270),
.D(n_2226),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2292),
.B(n_2239),
.Y(n_2324)
);

OAI21xp33_ASAP7_75t_L g2325 ( 
.A1(n_2289),
.A2(n_2236),
.B(n_2263),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2289),
.B(n_2239),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2292),
.B(n_2290),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2295),
.Y(n_2328)
);

O2A1O1Ixp5_ASAP7_75t_L g2329 ( 
.A1(n_2281),
.A2(n_2226),
.B(n_2259),
.C(n_2262),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2275),
.A2(n_2259),
.B(n_2253),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2302),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2307),
.Y(n_2332)
);

A2O1A1Ixp33_ASAP7_75t_L g2333 ( 
.A1(n_2278),
.A2(n_1917),
.B(n_1909),
.C(n_2103),
.Y(n_2333)
);

OAI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2284),
.A2(n_2288),
.B1(n_2278),
.B2(n_2287),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2279),
.B(n_2205),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2298),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_2285),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2309),
.B(n_2205),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2285),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2283),
.B(n_2208),
.Y(n_2340)
);

AOI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2282),
.A2(n_2296),
.B1(n_2294),
.B2(n_2286),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2312),
.A2(n_2208),
.B1(n_2210),
.B2(n_2103),
.Y(n_2342)
);

OAI322xp33_ASAP7_75t_L g2343 ( 
.A1(n_2306),
.A2(n_2299),
.A3(n_2286),
.B1(n_2315),
.B2(n_2308),
.C1(n_2291),
.C2(n_2303),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2313),
.Y(n_2344)
);

OAI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2301),
.A2(n_2253),
.B1(n_1917),
.B2(n_1909),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2337),
.Y(n_2346)
);

INVx1_ASAP7_75t_SL g2347 ( 
.A(n_2318),
.Y(n_2347)
);

NAND2xp33_ASAP7_75t_R g2348 ( 
.A(n_2324),
.B(n_2301),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2326),
.B(n_2325),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_R g2350 ( 
.A(n_2327),
.B(n_2304),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2326),
.B(n_2322),
.Y(n_2351)
);

NOR3xp33_ASAP7_75t_L g2352 ( 
.A(n_2334),
.B(n_2310),
.C(n_2298),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2337),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2319),
.B(n_2294),
.Y(n_2354)
);

OR2x2_ASAP7_75t_L g2355 ( 
.A(n_2323),
.B(n_2280),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2320),
.B(n_2301),
.Y(n_2356)
);

OAI21xp33_ASAP7_75t_SL g2357 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2305),
.Y(n_2357)
);

NAND2xp33_ASAP7_75t_SL g2358 ( 
.A(n_2341),
.B(n_2233),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2335),
.B(n_2210),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2339),
.Y(n_2360)
);

OAI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2329),
.A2(n_2253),
.B(n_2265),
.Y(n_2361)
);

INVxp67_ASAP7_75t_L g2362 ( 
.A(n_2317),
.Y(n_2362)
);

INVxp67_ASAP7_75t_L g2363 ( 
.A(n_2344),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2321),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2336),
.B(n_2233),
.Y(n_2365)
);

NOR2xp67_ASAP7_75t_SL g2366 ( 
.A(n_2330),
.B(n_1941),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2328),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2331),
.B(n_2240),
.Y(n_2368)
);

AOI211xp5_ASAP7_75t_L g2369 ( 
.A1(n_2343),
.A2(n_2266),
.B(n_2265),
.C(n_2247),
.Y(n_2369)
);

NOR3xp33_ASAP7_75t_L g2370 ( 
.A(n_2351),
.B(n_2358),
.C(n_2349),
.Y(n_2370)
);

AOI211xp5_ASAP7_75t_SL g2371 ( 
.A1(n_2362),
.A2(n_2333),
.B(n_2345),
.C(n_2338),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2363),
.B(n_2332),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2358),
.A2(n_2333),
.B(n_2316),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2360),
.B(n_2340),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2346),
.Y(n_2375)
);

NAND4xp75_ASAP7_75t_L g2376 ( 
.A(n_2357),
.B(n_2353),
.C(n_2356),
.D(n_2360),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2347),
.B(n_2340),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2355),
.B(n_2338),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2352),
.B(n_2341),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2368),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2364),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_2356),
.B(n_2342),
.Y(n_2382)
);

NAND4xp25_ASAP7_75t_L g2383 ( 
.A(n_2348),
.B(n_2266),
.C(n_2247),
.D(n_2240),
.Y(n_2383)
);

AOI211xp5_ASAP7_75t_L g2384 ( 
.A1(n_2354),
.A2(n_2350),
.B(n_2366),
.C(n_2361),
.Y(n_2384)
);

OAI211xp5_ASAP7_75t_SL g2385 ( 
.A1(n_2379),
.A2(n_2369),
.B(n_2367),
.C(n_2350),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2375),
.Y(n_2386)
);

OAI211xp5_ASAP7_75t_SL g2387 ( 
.A1(n_2384),
.A2(n_2365),
.B(n_2348),
.C(n_2345),
.Y(n_2387)
);

OAI221xp5_ASAP7_75t_SL g2388 ( 
.A1(n_2373),
.A2(n_2359),
.B1(n_2179),
.B2(n_2175),
.C(n_2167),
.Y(n_2388)
);

NOR4xp75_ASAP7_75t_L g2389 ( 
.A(n_2376),
.B(n_2144),
.C(n_2135),
.D(n_2137),
.Y(n_2389)
);

AOI221xp5_ASAP7_75t_L g2390 ( 
.A1(n_2370),
.A2(n_2217),
.B1(n_2179),
.B2(n_2175),
.C(n_2136),
.Y(n_2390)
);

OAI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2370),
.A2(n_2371),
.B1(n_2378),
.B2(n_2382),
.C(n_2377),
.Y(n_2391)
);

OAI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2374),
.A2(n_2179),
.B1(n_2175),
.B2(n_2125),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2372),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2383),
.A2(n_2125),
.B1(n_2103),
.B2(n_1958),
.Y(n_2394)
);

AOI21xp33_ASAP7_75t_SL g2395 ( 
.A1(n_2380),
.A2(n_2125),
.B(n_1909),
.Y(n_2395)
);

OAI211xp5_ASAP7_75t_L g2396 ( 
.A1(n_2381),
.A2(n_1941),
.B(n_2002),
.C(n_1917),
.Y(n_2396)
);

AOI322xp5_ASAP7_75t_L g2397 ( 
.A1(n_2379),
.A2(n_2129),
.A3(n_2113),
.B1(n_2121),
.B2(n_2125),
.C1(n_2154),
.C2(n_2145),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2385),
.A2(n_2391),
.B1(n_2387),
.B2(n_2394),
.Y(n_2398)
);

NOR3xp33_ASAP7_75t_L g2399 ( 
.A(n_2393),
.B(n_1941),
.C(n_2002),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2395),
.B(n_1975),
.Y(n_2400)
);

AOI211x1_ASAP7_75t_L g2401 ( 
.A1(n_2396),
.A2(n_2137),
.B(n_2135),
.C(n_2144),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2386),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2390),
.B(n_1975),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_R g2404 ( 
.A(n_2389),
.B(n_1958),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_2392),
.Y(n_2405)
);

AOI221xp5_ASAP7_75t_L g2406 ( 
.A1(n_2388),
.A2(n_2139),
.B1(n_2147),
.B2(n_2095),
.C(n_2096),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2397),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2386),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_2405),
.B(n_2154),
.Y(n_2409)
);

AOI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2407),
.A2(n_1958),
.B1(n_1975),
.B2(n_2139),
.Y(n_2410)
);

NOR3xp33_ASAP7_75t_L g2411 ( 
.A(n_2398),
.B(n_1980),
.C(n_2147),
.Y(n_2411)
);

XNOR2xp5_ASAP7_75t_L g2412 ( 
.A(n_2402),
.B(n_1922),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2408),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2399),
.B(n_2113),
.Y(n_2414)
);

AO22x2_ASAP7_75t_L g2415 ( 
.A1(n_2400),
.A2(n_2118),
.B1(n_2094),
.B2(n_2095),
.Y(n_2415)
);

AOI221x1_ASAP7_75t_L g2416 ( 
.A1(n_2404),
.A2(n_2096),
.B1(n_2094),
.B2(n_2104),
.C(n_2118),
.Y(n_2416)
);

OAI21xp33_ASAP7_75t_SL g2417 ( 
.A1(n_2403),
.A2(n_2121),
.B(n_2107),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2404),
.B(n_2123),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2409),
.Y(n_2419)
);

AND2x2_ASAP7_75t_SL g2420 ( 
.A(n_2411),
.B(n_2406),
.Y(n_2420)
);

INVx3_ASAP7_75t_SL g2421 ( 
.A(n_2413),
.Y(n_2421)
);

OAI21xp5_ASAP7_75t_SL g2422 ( 
.A1(n_2410),
.A2(n_2401),
.B(n_2000),
.Y(n_2422)
);

AO22x2_ASAP7_75t_L g2423 ( 
.A1(n_2418),
.A2(n_2416),
.B1(n_2414),
.B2(n_2412),
.Y(n_2423)
);

OAI221xp5_ASAP7_75t_L g2424 ( 
.A1(n_2417),
.A2(n_2415),
.B1(n_2115),
.B2(n_2107),
.C(n_2104),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2415),
.A2(n_2115),
.B1(n_2119),
.B2(n_2150),
.Y(n_2425)
);

OR2x2_ASAP7_75t_L g2426 ( 
.A(n_2419),
.B(n_2127),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_2421),
.Y(n_2427)
);

CKINVDCx20_ASAP7_75t_R g2428 ( 
.A(n_2423),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2420),
.B(n_2122),
.Y(n_2429)
);

OAI22x1_ASAP7_75t_L g2430 ( 
.A1(n_2427),
.A2(n_2422),
.B1(n_2424),
.B2(n_2425),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2429),
.B(n_2122),
.Y(n_2431)
);

AOI22x1_ASAP7_75t_L g2432 ( 
.A1(n_2430),
.A2(n_2426),
.B1(n_2428),
.B2(n_2431),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2432),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2432),
.Y(n_2434)
);

OAI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2433),
.A2(n_2428),
.B(n_2123),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2434),
.A2(n_1968),
.B(n_2119),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2435),
.Y(n_2437)
);

AOI22xp33_ASAP7_75t_L g2438 ( 
.A1(n_2436),
.A2(n_1975),
.B1(n_2153),
.B2(n_2150),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2437),
.A2(n_1975),
.B1(n_2153),
.B2(n_2160),
.Y(n_2439)
);

OAI221xp5_ASAP7_75t_L g2440 ( 
.A1(n_2439),
.A2(n_2438),
.B1(n_2127),
.B2(n_2126),
.C(n_2160),
.Y(n_2440)
);

AOI211xp5_ASAP7_75t_L g2441 ( 
.A1(n_2440),
.A2(n_2126),
.B(n_1975),
.C(n_2145),
.Y(n_2441)
);


endmodule