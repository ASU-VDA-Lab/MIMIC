module fake_netlist_6_986_n_2043 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2043);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2043;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_SL g200 ( 
.A(n_78),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_27),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_100),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_51),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_69),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_88),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_190),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_64),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_13),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_15),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_38),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_150),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_54),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_129),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_127),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_64),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_66),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_93),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_57),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_92),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_56),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_169),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_77),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_54),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_38),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_124),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_84),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_86),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_22),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_133),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_25),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_67),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_199),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_69),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_116),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_120),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_98),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_140),
.Y(n_261)
);

CKINVDCx11_ASAP7_75t_R g262 ( 
.A(n_89),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_188),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_144),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_61),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_23),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_99),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_30),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_115),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_82),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_118),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_51),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_48),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_162),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_106),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_134),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_18),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_148),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_52),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_95),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_122),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_67),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_71),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_117),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_10),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_76),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_10),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_156),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_175),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_173),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_114),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_149),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_105),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_63),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_136),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_152),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_167),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_91),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_198),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_131),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_110),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_174),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_103),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_154),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_85),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_16),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_2),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_158),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_171),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_96),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_182),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_4),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_25),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_191),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_5),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_70),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_181),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_28),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_125),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_147),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_68),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_170),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_111),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_63),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_28),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_23),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_41),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_196),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_163),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_101),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_19),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_130),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_30),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_36),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_58),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_0),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_195),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_172),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_79),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_65),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_13),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_141),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_46),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_132),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_160),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_151),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_73),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_12),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_83),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_104),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_49),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_102),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_161),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_0),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_44),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_113),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_26),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_20),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_74),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_59),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_194),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_166),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_185),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_52),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_16),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_45),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_70),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_59),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_68),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_27),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_60),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_12),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_9),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_65),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_19),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_48),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_3),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_1),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_39),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_50),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_3),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_159),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_15),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_29),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_33),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_41),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_192),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_8),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_119),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_121),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_213),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_262),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_285),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_298),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_304),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_256),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_267),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_257),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_261),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_264),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_313),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_201),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_350),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_265),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_273),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_230),
.B(n_6),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_274),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_278),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_283),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_370),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_326),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_399),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_286),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_225),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_226),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_281),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_289),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_338),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_245),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g439 ( 
.A(n_201),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_345),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_291),
.B(n_7),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_245),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_293),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_297),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_301),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_245),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_228),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_203),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_303),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_245),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_306),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_245),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_329),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_344),
.B(n_7),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_213),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_296),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_307),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_329),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_329),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_308),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_329),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_311),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_329),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_317),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_292),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_318),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_319),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_322),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_325),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_296),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_203),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_292),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_247),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_200),
.B(n_8),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_327),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_330),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_331),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_353),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_200),
.B(n_9),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_358),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_361),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_371),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_344),
.B(n_11),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_384),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_391),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_396),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_246),
.B(n_14),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_379),
.B(n_14),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_393),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_205),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_204),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_499),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_465),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_438),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_465),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_246),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_465),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_465),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_400),
.A2(n_227),
.B(n_217),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_465),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_442),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_448),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_476),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_217),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_227),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

AND3x2_ASAP7_75t_L g522 ( 
.A(n_478),
.B(n_335),
.C(n_295),
.Y(n_522)
);

BUFx8_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_400),
.B(n_269),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_450),
.Y(n_527)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_475),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_489),
.B(n_269),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_452),
.Y(n_532)
);

OA21x2_ASAP7_75t_L g533 ( 
.A1(n_408),
.A2(n_248),
.B(n_219),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_408),
.A2(n_276),
.B(n_271),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_500),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_476),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_476),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_453),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_494),
.B(n_224),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_416),
.B(n_271),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_458),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_405),
.A2(n_332),
.B1(n_387),
.B2(n_389),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_458),
.Y(n_546)
);

BUFx8_ASAP7_75t_L g547 ( 
.A(n_486),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_416),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_420),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_425),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_425),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_428),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_401),
.B(n_276),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_461),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g559 ( 
.A1(n_428),
.A2(n_437),
.B(n_463),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_401),
.B(n_379),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_463),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_467),
.B(n_202),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_455),
.B(n_388),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_402),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_469),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_469),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_471),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_471),
.B(n_209),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_490),
.B(n_214),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_443),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_495),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_495),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_421),
.B(n_250),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_580),
.B(n_434),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_508),
.B(n_410),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_533),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_R g586 ( 
.A(n_508),
.B(n_415),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_532),
.B(n_409),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_411),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_514),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_533),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_510),
.B(n_441),
.C(n_496),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_412),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_577),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_510),
.B(n_413),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_532),
.B(n_418),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_519),
.A2(n_477),
.B1(n_488),
.B2(n_454),
.Y(n_599)
);

BUFx6f_ASAP7_75t_SL g600 ( 
.A(n_530),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_542),
.B(n_419),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_545),
.A2(n_223),
.B1(n_508),
.B2(n_324),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_577),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_523),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_523),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_533),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_533),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_555),
.B(n_560),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_559),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_532),
.B(n_422),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_532),
.B(n_424),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_532),
.B(n_426),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

NOR2x1p5_ASAP7_75t_L g616 ( 
.A(n_560),
.B(n_388),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_542),
.B(n_431),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_532),
.B(n_435),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_514),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_519),
.B(n_444),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_517),
.B(n_410),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_560),
.B(n_204),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_519),
.B(n_451),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_555),
.B(n_456),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_560),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_517),
.B(n_434),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_519),
.B(n_460),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_542),
.B(n_462),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_503),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_503),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_562),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_542),
.B(n_440),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_520),
.B(n_464),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_559),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_520),
.B(n_466),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_529),
.B(n_470),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_529),
.B(n_472),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_520),
.B(n_480),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_509),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_559),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_559),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_520),
.B(n_473),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_545),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_559),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_562),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_555),
.B(n_455),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_530),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_555),
.B(n_486),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_481),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_514),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_514),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_536),
.B(n_482),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_536),
.B(n_485),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_509),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_501),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_561),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_565),
.B(n_496),
.Y(n_665)
);

NAND3xp33_ASAP7_75t_L g666 ( 
.A(n_525),
.B(n_488),
.C(n_454),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_561),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_565),
.B(n_491),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_530),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_565),
.B(n_447),
.Y(n_670)
);

OAI21xp33_ASAP7_75t_SL g671 ( 
.A1(n_513),
.A2(n_365),
.B(n_248),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_530),
.B(n_493),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_530),
.B(n_440),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_548),
.B(n_292),
.Y(n_676)
);

INVx4_ASAP7_75t_SL g677 ( 
.A(n_528),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_561),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_548),
.B(n_310),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_549),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_563),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_569),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_523),
.B(n_439),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_549),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_523),
.B(n_445),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_565),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_509),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_514),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_548),
.B(n_449),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_523),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_514),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_548),
.B(n_534),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_548),
.B(n_457),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_514),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_514),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_549),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_549),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_525),
.B(n_241),
.C(n_233),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_545),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_550),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_547),
.Y(n_701)
);

AND2x6_ASAP7_75t_L g702 ( 
.A(n_550),
.B(n_292),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_547),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_509),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_522),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_569),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_550),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_569),
.Y(n_708)
);

OAI21xp33_ASAP7_75t_SL g709 ( 
.A1(n_513),
.A2(n_365),
.B(n_219),
.Y(n_709)
);

AND2x2_ASAP7_75t_SL g710 ( 
.A(n_548),
.B(n_292),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_534),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_514),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_509),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_550),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_509),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_569),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_534),
.B(n_429),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_572),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_534),
.B(n_382),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_572),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_552),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_552),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_509),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_522),
.B(n_468),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_540),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_547),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_572),
.Y(n_728)
);

BUFx8_ASAP7_75t_SL g729 ( 
.A(n_501),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_552),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_540),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_541),
.B(n_242),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_576),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_676),
.B(n_547),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_SL g735 ( 
.A(n_606),
.B(n_566),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_621),
.A2(n_484),
.B1(n_487),
.B2(n_479),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_595),
.B(n_541),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_646),
.B(n_541),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_655),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_594),
.B(n_630),
.C(n_617),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_669),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_646),
.B(n_541),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_669),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_610),
.B(n_625),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_676),
.B(n_547),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_665),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_597),
.B(n_432),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_646),
.B(n_558),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_646),
.B(n_558),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_582),
.B(n_433),
.Y(n_751)
);

O2A1O1Ixp5_ASAP7_75t_L g752 ( 
.A1(n_581),
.A2(n_543),
.B(n_525),
.C(n_564),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_625),
.B(n_558),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_610),
.B(n_558),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_627),
.B(n_552),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_611),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_611),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_666),
.B(n_564),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_624),
.B(n_436),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_676),
.B(n_547),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_629),
.B(n_637),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_633),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_640),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_627),
.B(n_553),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_639),
.B(n_566),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_686),
.B(n_553),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_584),
.B(n_501),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_686),
.B(n_553),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_710),
.B(n_553),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_710),
.B(n_554),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_633),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_710),
.B(n_347),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_584),
.B(n_207),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_626),
.B(n_347),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_638),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_638),
.B(n_554),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_665),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_720),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_644),
.B(n_554),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_644),
.B(n_645),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_645),
.B(n_554),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_670),
.B(n_564),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_670),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_581),
.B(n_316),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_626),
.B(n_347),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_642),
.B(n_403),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_711),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_606),
.B(n_404),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_720),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_649),
.B(n_543),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_651),
.B(n_244),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_656),
.B(n_406),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_626),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_649),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_651),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_656),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_711),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_585),
.B(n_316),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_641),
.B(n_414),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_718),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_666),
.B(n_543),
.Y(n_801)
);

NOR3xp33_ASAP7_75t_L g802 ( 
.A(n_647),
.B(n_376),
.C(n_339),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_626),
.B(n_347),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_585),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_657),
.B(n_568),
.Y(n_805)
);

BUFx6f_ASAP7_75t_SL g806 ( 
.A(n_603),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_589),
.A2(n_535),
.B1(n_513),
.B2(n_252),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_589),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_672),
.B(n_568),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_587),
.B(n_568),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_660),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_598),
.B(n_612),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_613),
.B(n_568),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_614),
.B(n_347),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_619),
.B(n_505),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_591),
.A2(n_574),
.B(n_570),
.C(n_394),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_591),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_604),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_689),
.B(n_372),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_662),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_652),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_692),
.A2(n_574),
.B(n_570),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_663),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_662),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_693),
.B(n_675),
.Y(n_826)
);

OAI22x1_ASAP7_75t_R g827 ( 
.A1(n_647),
.A2(n_427),
.B1(n_430),
.B2(n_417),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_718),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_616),
.B(n_258),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_616),
.B(n_260),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_668),
.B(n_205),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_679),
.B(n_372),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_L g833 ( 
.A(n_594),
.B(n_599),
.C(n_588),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_604),
.B(n_372),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_608),
.B(n_609),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_586),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_608),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_623),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_664),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_623),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_609),
.B(n_664),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_727),
.B(n_316),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_601),
.A2(n_208),
.B1(n_210),
.B2(n_346),
.Y(n_843)
);

AND2x6_ASAP7_75t_SL g844 ( 
.A(n_725),
.B(n_249),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_622),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_667),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_673),
.B(n_505),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_673),
.B(n_505),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_600),
.A2(n_636),
.B1(n_727),
.B2(n_705),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_674),
.B(n_506),
.Y(n_850)
);

BUFx6f_ASAP7_75t_SL g851 ( 
.A(n_603),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_628),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_674),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_622),
.B(n_206),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_L g855 ( 
.A(n_678),
.B(n_316),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_678),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_705),
.B(n_208),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_703),
.B(n_570),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_628),
.B(n_210),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_583),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_583),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_732),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_671),
.B(n_372),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_L g864 ( 
.A(n_602),
.B(n_251),
.C(n_243),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_590),
.B(n_506),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_699),
.B(n_211),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_635),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_662),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_671),
.B(n_709),
.Y(n_869)
);

NOR2x1p5_ASAP7_75t_L g870 ( 
.A(n_607),
.B(n_206),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_590),
.B(n_506),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_590),
.B(n_507),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_600),
.A2(n_235),
.B1(n_352),
.B2(n_346),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_683),
.B(n_211),
.Y(n_874)
);

AND2x6_ASAP7_75t_SL g875 ( 
.A(n_729),
.B(n_253),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_602),
.B(n_212),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_596),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_590),
.B(n_507),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_620),
.B(n_507),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_685),
.B(n_596),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_709),
.B(n_372),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_635),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_600),
.B(n_218),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_662),
.B(n_316),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_620),
.B(n_516),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_662),
.B(n_316),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_687),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_698),
.B(n_255),
.C(n_254),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_687),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_620),
.B(n_516),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_620),
.B(n_516),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_592),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_687),
.B(n_713),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_607),
.B(n_574),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_712),
.B(n_218),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_658),
.B(n_521),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_687),
.B(n_316),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_618),
.B(n_382),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_687),
.B(n_316),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_658),
.B(n_521),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_698),
.A2(n_684),
.B1(n_696),
.B2(n_680),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_618),
.A2(n_272),
.B1(n_279),
.B2(n_299),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_658),
.B(n_521),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_737),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_737),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_800),
.B(n_828),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_761),
.B(n_680),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_763),
.B(n_690),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_774),
.A2(n_696),
.B(n_684),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_782),
.B(n_697),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_SL g911 ( 
.A1(n_772),
.A2(n_300),
.B(n_309),
.C(n_305),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_782),
.B(n_697),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_741),
.A2(n_701),
.B1(n_328),
.B2(n_336),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_745),
.A2(n_513),
.B(n_535),
.C(n_394),
.Y(n_914)
);

OAI21xp33_ASAP7_75t_L g915 ( 
.A1(n_866),
.A2(n_215),
.B(n_212),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_745),
.B(n_700),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_790),
.A2(n_681),
.B(n_712),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_835),
.A2(n_681),
.B(n_712),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_804),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_812),
.B(n_713),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_744),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_787),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_744),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_801),
.A2(n_681),
.B(n_712),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_820),
.A2(n_337),
.B(n_312),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_780),
.A2(n_715),
.B(n_713),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_793),
.B(n_713),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_738),
.B(n_783),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_776),
.A2(n_715),
.B(n_713),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_779),
.A2(n_715),
.B(n_653),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_806),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_833),
.A2(n_360),
.B1(n_357),
.B2(n_700),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_793),
.B(n_715),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_793),
.B(n_715),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_827),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_822),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_811),
.B(n_603),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_814),
.B(n_603),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_783),
.B(n_707),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_774),
.A2(n_714),
.B(n_707),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_862),
.B(n_714),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_785),
.A2(n_723),
.B(n_722),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_821),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_785),
.A2(n_723),
.B(n_722),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_781),
.A2(n_653),
.B(n_643),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_758),
.B(n_643),
.Y(n_946)
);

OR2x6_ASAP7_75t_L g947 ( 
.A(n_852),
.B(n_290),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_787),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_739),
.A2(n_653),
.B(n_643),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_862),
.B(n_730),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_808),
.B(n_704),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_831),
.B(n_730),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_818),
.B(n_819),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_778),
.B(n_704),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_803),
.A2(n_535),
.B(n_593),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_860),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_826),
.A2(n_334),
.B(n_397),
.C(n_381),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_874),
.A2(n_535),
.B(n_320),
.C(n_359),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_736),
.B(n_222),
.C(n_221),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_756),
.A2(n_704),
.B1(n_724),
.B2(n_231),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_800),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_743),
.A2(n_653),
.B(n_724),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_749),
.A2(n_750),
.B(n_754),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_803),
.A2(n_653),
.B(n_724),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_789),
.B(n_658),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_893),
.A2(n_653),
.B(n_659),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_753),
.B(n_659),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_893),
.A2(n_688),
.B(n_659),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_816),
.B(n_818),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_805),
.A2(n_688),
.B(n_659),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_809),
.A2(n_691),
.B(n_688),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_824),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_752),
.A2(n_605),
.B(n_593),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_819),
.B(n_688),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_828),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_837),
.B(n_691),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_845),
.B(n_215),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_826),
.A2(n_302),
.B(n_366),
.C(n_733),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_837),
.B(n_691),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_810),
.A2(n_694),
.B(n_691),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_834),
.A2(n_615),
.B(n_605),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_813),
.A2(n_695),
.B(n_694),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_755),
.A2(n_695),
.B(n_694),
.Y(n_983)
);

AND2x2_ASAP7_75t_SL g984 ( 
.A(n_842),
.B(n_524),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_756),
.B(n_694),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_839),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_764),
.A2(n_726),
.B(n_695),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_757),
.B(n_762),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_786),
.A2(n_695),
.B1(n_731),
.B2(n_726),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_766),
.A2(n_768),
.B(n_823),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_759),
.A2(n_726),
.B1(n_731),
.B2(n_222),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_834),
.A2(n_731),
.B(n_726),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_769),
.A2(n_731),
.B(n_504),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_757),
.B(n_615),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_841),
.A2(n_632),
.B(n_631),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_821),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_762),
.A2(n_221),
.B1(n_231),
.B2(n_235),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_771),
.B(n_631),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_770),
.A2(n_504),
.B(n_632),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_796),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_792),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_765),
.B(n_859),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_852),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_771),
.A2(n_216),
.B(n_220),
.C(n_229),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_773),
.B(n_326),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_775),
.B(n_634),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_775),
.B(n_634),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_784),
.A2(n_504),
.B(n_509),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_794),
.B(n_677),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_794),
.B(n_648),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_784),
.A2(n_504),
.B(n_509),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_767),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_841),
.A2(n_650),
.B(n_648),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_740),
.B(n_650),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_894),
.B(n_858),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_SL g1016 ( 
.A(n_877),
.B(n_354),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_836),
.B(n_259),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_747),
.B(n_654),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_849),
.B(n_677),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_734),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_798),
.A2(n_504),
.B(n_515),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_829),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_777),
.B(n_654),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_821),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_798),
.A2(n_504),
.B(n_515),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_795),
.A2(n_772),
.B(n_820),
.C(n_869),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_825),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_869),
.A2(n_807),
.B(n_817),
.Y(n_1028)
);

AOI33xp33_ASAP7_75t_L g1029 ( 
.A1(n_838),
.A2(n_840),
.A3(n_830),
.B1(n_829),
.B2(n_791),
.B3(n_843),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_842),
.A2(n_815),
.B(n_825),
.Y(n_1030)
);

AOI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_748),
.A2(n_266),
.B(n_263),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_799),
.B(n_326),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_742),
.B(n_682),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_751),
.B(n_268),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_861),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_791),
.B(n_682),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_892),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_825),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_791),
.B(n_706),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_797),
.B(n_706),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_880),
.B(n_239),
.C(n_236),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_876),
.B(n_270),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_815),
.A2(n_504),
.B(n_515),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_892),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_895),
.B(n_708),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_846),
.A2(n_856),
.B(n_853),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_865),
.A2(n_716),
.B(n_708),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_838),
.B(n_677),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_840),
.B(n_677),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_857),
.B(n_716),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_868),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_806),
.B(n_354),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_898),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_863),
.A2(n_733),
.B(n_728),
.C(n_721),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_854),
.B(n_275),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_867),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_870),
.B(n_524),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_868),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_868),
.A2(n_504),
.B(n_515),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_864),
.B(n_735),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_734),
.A2(n_398),
.B1(n_340),
.B2(n_352),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_887),
.A2(n_504),
.B(n_515),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_887),
.A2(n_504),
.B(n_515),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_887),
.A2(n_531),
.B(n_515),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_788),
.B(n_280),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_871),
.A2(n_719),
.B(n_717),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_802),
.B(n_829),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_746),
.B(n_240),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_746),
.A2(n_349),
.B1(n_220),
.B2(n_229),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_832),
.A2(n_728),
.B(n_721),
.C(n_719),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_882),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_830),
.B(n_717),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_889),
.A2(n_515),
.B(n_531),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_889),
.A2(n_515),
.B(n_531),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_830),
.B(n_524),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_883),
.B(n_526),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_889),
.A2(n_531),
.B(n_540),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_847),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_832),
.A2(n_511),
.B(n_537),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_872),
.A2(n_531),
.B(n_540),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_898),
.B(n_340),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_898),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_878),
.A2(n_531),
.B(n_540),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_760),
.A2(n_398),
.B1(n_373),
.B2(n_321),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_848),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_850),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_901),
.B(n_879),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_760),
.B(n_540),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_888),
.A2(n_556),
.B1(n_579),
.B2(n_578),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_969),
.A2(n_898),
.B1(n_873),
.B2(n_881),
.Y(n_1090)
);

OAI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_1034),
.A2(n_232),
.B(n_216),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1012),
.B(n_902),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1034),
.A2(n_1002),
.B(n_1042),
.C(n_1026),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1060),
.A2(n_1067),
.B1(n_906),
.B2(n_1001),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_1031),
.B(n_284),
.C(n_282),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_SL g1096 ( 
.A(n_972),
.B(n_806),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1032),
.B(n_287),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1069),
.A2(n_907),
.B1(n_984),
.B2(n_1028),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_1003),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_1000),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_963),
.A2(n_890),
.B(n_885),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1069),
.A2(n_863),
.B1(n_881),
.B2(n_851),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_919),
.Y(n_1103)
);

INVx3_ASAP7_75t_SL g1104 ( 
.A(n_931),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1086),
.B(n_891),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_SL g1106 ( 
.A1(n_958),
.A2(n_899),
.B(n_897),
.C(n_886),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_990),
.A2(n_903),
.B(n_900),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1042),
.A2(n_855),
.B(n_899),
.C(n_886),
.Y(n_1108)
);

AOI22x1_ASAP7_75t_L g1109 ( 
.A1(n_1030),
.A2(n_855),
.B1(n_526),
.B2(n_579),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_906),
.B(n_884),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1045),
.A2(n_896),
.B(n_897),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_L g1112 ( 
.A(n_1041),
.B(n_288),
.C(n_395),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1078),
.B(n_884),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1060),
.A2(n_959),
.B1(n_1022),
.B2(n_1017),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_922),
.B(n_851),
.Y(n_1115)
);

AND2x6_ASAP7_75t_SL g1116 ( 
.A(n_908),
.B(n_1065),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1029),
.A2(n_294),
.B(n_314),
.C(n_315),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_924),
.A2(n_917),
.B(n_920),
.Y(n_1118)
);

BUFx4f_ASAP7_75t_SL g1119 ( 
.A(n_922),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1016),
.A2(n_354),
.B1(n_364),
.B2(n_234),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_927),
.A2(n_531),
.B(n_540),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_937),
.B(n_844),
.Y(n_1122)
);

O2A1O1Ixp5_ASAP7_75t_L g1123 ( 
.A1(n_1015),
.A2(n_551),
.B(n_526),
.C(n_579),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_913),
.A2(n_557),
.B(n_571),
.C(n_567),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1005),
.B(n_323),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_927),
.A2(n_531),
.B(n_540),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_1000),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_961),
.B(n_75),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_977),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1078),
.B(n_527),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_933),
.A2(n_531),
.B(n_540),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_R g1132 ( 
.A(n_935),
.B(n_875),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1085),
.B(n_527),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_364),
.B1(n_578),
.B2(n_527),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_947),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1085),
.B(n_538),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_975),
.B(n_538),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_933),
.A2(n_540),
.B(n_539),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_936),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1084),
.A2(n_567),
.B(n_571),
.C(n_557),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_908),
.B(n_364),
.Y(n_1141)
);

INVx11_ASAP7_75t_L g1142 ( 
.A(n_1057),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1055),
.B(n_938),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_910),
.B(n_538),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1004),
.A2(n_571),
.B(n_567),
.C(n_557),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_934),
.A2(n_539),
.B(n_512),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1004),
.A2(n_544),
.B(n_556),
.C(n_551),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_934),
.A2(n_539),
.B(n_512),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_956),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_926),
.A2(n_539),
.B(n_512),
.Y(n_1151)
);

AOI22x1_ASAP7_75t_L g1152 ( 
.A1(n_970),
.A2(n_980),
.B1(n_982),
.B2(n_971),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1029),
.A2(n_392),
.B(n_390),
.C(n_369),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_920),
.A2(n_918),
.B(n_967),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_937),
.A2(n_556),
.B1(n_578),
.B2(n_544),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_915),
.A2(n_551),
.B(n_546),
.C(n_544),
.Y(n_1156)
);

AO32x2_ASAP7_75t_L g1157 ( 
.A1(n_932),
.A2(n_17),
.A3(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_1157)
);

CKINVDCx16_ASAP7_75t_R g1158 ( 
.A(n_1052),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_975),
.B(n_546),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_912),
.A2(n_539),
.B(n_511),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_947),
.Y(n_1161)
);

AND2x2_ASAP7_75t_SL g1162 ( 
.A(n_1065),
.B(n_17),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_948),
.B(n_961),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_995),
.A2(n_573),
.B(n_546),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_948),
.B(n_333),
.Y(n_1165)
);

OAI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_947),
.A2(n_234),
.B1(n_355),
.B2(n_351),
.Y(n_1166)
);

AOI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1035),
.A2(n_576),
.B1(n_573),
.B2(n_356),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1037),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1055),
.A2(n_368),
.B(n_367),
.C(n_363),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1088),
.A2(n_537),
.B(n_512),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1053),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1082),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1088),
.A2(n_539),
.B(n_511),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_928),
.B(n_362),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1081),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1081),
.B(n_232),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_1020),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1082),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1049),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_1068),
.A2(n_957),
.B(n_973),
.C(n_978),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_916),
.B(n_573),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1087),
.A2(n_341),
.B1(n_277),
.B2(n_238),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_986),
.B(n_80),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1076),
.B(n_237),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1049),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_923),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_929),
.A2(n_511),
.B(n_518),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1075),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_952),
.B(n_342),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_941),
.B(n_573),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_939),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_904),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_905),
.B(n_342),
.Y(n_1194)
);

OAI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_997),
.A2(n_343),
.B(n_348),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_921),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1015),
.B(n_343),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_950),
.B(n_1050),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1061),
.Y(n_1199)
);

OR2x6_ASAP7_75t_SL g1200 ( 
.A(n_1056),
.B(n_348),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1018),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1071),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1023),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1024),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_953),
.B(n_573),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1024),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_953),
.B(n_573),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1072),
.B(n_349),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1072),
.B(n_351),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_988),
.A2(n_385),
.B1(n_375),
.B2(n_377),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1046),
.B(n_355),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1024),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_994),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_988),
.B(n_576),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1040),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_998),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1033),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1036),
.A2(n_1039),
.B(n_946),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_958),
.A2(n_576),
.B(n_537),
.C(n_518),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1024),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_946),
.A2(n_537),
.B(n_518),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_965),
.B(n_518),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1027),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_914),
.A2(n_380),
.B1(n_378),
.B2(n_377),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1027),
.B(n_139),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_996),
.B(n_575),
.Y(n_1226)
);

AOI33xp33_ASAP7_75t_L g1227 ( 
.A1(n_911),
.A2(n_380),
.A3(n_378),
.B1(n_375),
.B2(n_29),
.B3(n_31),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1027),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1006),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_954),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_996),
.B(n_21),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_991),
.A2(n_575),
.B(n_563),
.C(n_31),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_989),
.A2(n_575),
.B(n_563),
.C(n_32),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_943),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_914),
.A2(n_702),
.B(n_528),
.Y(n_1235)
);

AND2x6_ASAP7_75t_L g1236 ( 
.A(n_1058),
.B(n_563),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1010),
.A2(n_528),
.B1(n_575),
.B2(n_563),
.Y(n_1237)
);

INVx6_ASAP7_75t_L g1238 ( 
.A(n_1027),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1058),
.B(n_24),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1014),
.B(n_26),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1038),
.B(n_32),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1093),
.A2(n_1185),
.B(n_1190),
.C(n_1098),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1169),
.A2(n_911),
.B(n_1019),
.C(n_960),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1119),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1098),
.A2(n_999),
.B(n_983),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1108),
.A2(n_987),
.B(n_940),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1107),
.A2(n_944),
.B(n_1019),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1143),
.B(n_1007),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1139),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1101),
.A2(n_955),
.B(n_930),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1090),
.A2(n_993),
.B(n_1070),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_1115),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1164),
.A2(n_1118),
.B(n_1152),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1154),
.A2(n_985),
.B(n_974),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1103),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1149),
.Y(n_1256)
);

OAI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1120),
.A2(n_1089),
.B1(n_1013),
.B2(n_1047),
.C(n_1066),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1192),
.B(n_979),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1118),
.A2(n_1079),
.B(n_909),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1090),
.A2(n_1051),
.B(n_1054),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1218),
.A2(n_962),
.B(n_949),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1198),
.A2(n_943),
.B(n_945),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1201),
.B(n_976),
.Y(n_1263)
);

AOI221x1_ASAP7_75t_L g1264 ( 
.A1(n_1102),
.A2(n_992),
.B1(n_981),
.B2(n_964),
.C(n_968),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1117),
.A2(n_1048),
.B(n_1009),
.C(n_951),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1097),
.B(n_1038),
.Y(n_1266)
);

OA22x2_ASAP7_75t_L g1267 ( 
.A1(n_1129),
.A2(n_1048),
.B1(n_1009),
.B2(n_951),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1170),
.A2(n_942),
.B(n_1083),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1182),
.A2(n_925),
.B1(n_976),
.B2(n_1080),
.C(n_1043),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1127),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1149),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1114),
.B(n_943),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1102),
.A2(n_1051),
.A3(n_1008),
.B(n_1011),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1198),
.A2(n_943),
.B(n_966),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1197),
.A2(n_1021),
.B(n_1025),
.C(n_1073),
.Y(n_1275)
);

BUFx2_ASAP7_75t_R g1276 ( 
.A(n_1104),
.Y(n_1276)
);

AO32x2_ASAP7_75t_L g1277 ( 
.A1(n_1224),
.A2(n_1038),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_1277)
);

AO21x1_ASAP7_75t_L g1278 ( 
.A1(n_1240),
.A2(n_1074),
.B(n_1064),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1203),
.B(n_1038),
.Y(n_1279)
);

AO32x2_ASAP7_75t_L g1280 ( 
.A1(n_1224),
.A2(n_33),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1115),
.B(n_1077),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1179),
.Y(n_1282)
);

OAI22x1_ASAP7_75t_L g1283 ( 
.A1(n_1094),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1199),
.A2(n_1062),
.B1(n_1059),
.B2(n_1063),
.Y(n_1284)
);

AOI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1111),
.A2(n_702),
.B(n_575),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1125),
.B(n_40),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1105),
.A2(n_528),
.B1(n_563),
.B2(n_575),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1158),
.B(n_563),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1193),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1122),
.B(n_42),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1174),
.B(n_43),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1099),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1111),
.A2(n_702),
.B(n_575),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_L g1294 ( 
.A(n_1141),
.B(n_563),
.C(n_575),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1232),
.A2(n_702),
.A3(n_44),
.B(n_45),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1180),
.A2(n_575),
.B(n_563),
.Y(n_1296)
);

AOI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1144),
.A2(n_1170),
.B(n_1222),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1105),
.A2(n_575),
.B(n_563),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1091),
.A2(n_43),
.B(n_46),
.C(n_47),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1100),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1092),
.B(n_47),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1208),
.B(n_49),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1153),
.A2(n_107),
.B(n_197),
.C(n_193),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1116),
.B(n_53),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1149),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1162),
.A2(n_702),
.B1(n_528),
.B2(n_57),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_SL g1307 ( 
.A(n_1095),
.B(n_1134),
.C(n_1195),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1233),
.A2(n_94),
.B(n_184),
.C(n_180),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1113),
.A2(n_702),
.B(n_90),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1196),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1113),
.A2(n_702),
.B(n_87),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1215),
.A2(n_135),
.B(n_177),
.Y(n_1312)
);

NAND3xp33_ASAP7_75t_L g1313 ( 
.A(n_1182),
.B(n_1112),
.C(n_1209),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1106),
.A2(n_108),
.B(n_176),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1231),
.A2(n_60),
.A3(n_61),
.B(n_62),
.Y(n_1315)
);

NOR2xp67_ASAP7_75t_L g1316 ( 
.A(n_1189),
.B(n_1179),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1144),
.A2(n_123),
.B(n_155),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1234),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1171),
.Y(n_1319)
);

AO21x2_ASAP7_75t_L g1320 ( 
.A1(n_1235),
.A2(n_109),
.B(n_143),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1220),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1123),
.A2(n_528),
.B(n_128),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1177),
.A2(n_528),
.B1(n_72),
.B2(n_73),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1234),
.A2(n_528),
.B(n_1128),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1217),
.A2(n_1202),
.B1(n_1186),
.B2(n_1230),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1161),
.B(n_1135),
.Y(n_1326)
);

NAND2x1_ASAP7_75t_L g1327 ( 
.A(n_1238),
.B(n_1137),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1186),
.B(n_1223),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1175),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1211),
.A2(n_1110),
.B1(n_1183),
.B2(n_1176),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1213),
.B(n_1216),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1187),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1150),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1142),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1181),
.A2(n_1133),
.B(n_1130),
.Y(n_1335)
);

AO32x2_ASAP7_75t_L g1336 ( 
.A1(n_1210),
.A2(n_1157),
.A3(n_1237),
.B1(n_1227),
.B2(n_1147),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1172),
.B(n_1110),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1181),
.A2(n_1133),
.B(n_1136),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1229),
.B(n_1194),
.Y(n_1339)
);

BUFx10_ASAP7_75t_L g1340 ( 
.A(n_1128),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1200),
.Y(n_1341)
);

BUFx10_ASAP7_75t_L g1342 ( 
.A(n_1239),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1130),
.B(n_1136),
.Y(n_1343)
);

AOI31xp67_ASAP7_75t_L g1344 ( 
.A1(n_1155),
.A2(n_1222),
.A3(n_1214),
.B(n_1191),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1178),
.A2(n_1165),
.B1(n_1241),
.B2(n_1163),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1210),
.B(n_1168),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1184),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1214),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1205),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1220),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1188),
.A2(n_1151),
.B(n_1221),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1166),
.B(n_1191),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1205),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1212),
.B(n_1228),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1096),
.Y(n_1356)
);

AO22x2_ASAP7_75t_L g1357 ( 
.A1(n_1157),
.A2(n_1225),
.B1(n_1235),
.B2(n_1207),
.Y(n_1357)
);

AO32x2_ASAP7_75t_L g1358 ( 
.A1(n_1157),
.A2(n_1237),
.A3(n_1145),
.B1(n_1219),
.B2(n_1167),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1156),
.A2(n_1140),
.B(n_1160),
.C(n_1124),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1109),
.A2(n_1173),
.B(n_1207),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1226),
.A2(n_1148),
.B(n_1146),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1138),
.A2(n_1226),
.B(n_1126),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1137),
.A2(n_1159),
.B(n_1121),
.Y(n_1363)
);

BUFx2_ASAP7_75t_R g1364 ( 
.A(n_1132),
.Y(n_1364)
);

O2A1O1Ixp5_ASAP7_75t_L g1365 ( 
.A1(n_1131),
.A2(n_1225),
.B(n_1159),
.C(n_1137),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1163),
.A2(n_1236),
.B(n_1159),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1236),
.A2(n_1238),
.B(n_1220),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1236),
.A2(n_990),
.B(n_1107),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1236),
.A2(n_990),
.B(n_1107),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1236),
.A2(n_990),
.B(n_1107),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1238),
.A2(n_1093),
.B(n_1002),
.C(n_1034),
.Y(n_1371)
);

AOI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1118),
.A2(n_1088),
.B(n_1154),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1149),
.Y(n_1373)
);

AO31x2_ASAP7_75t_L g1374 ( 
.A1(n_1118),
.A2(n_1098),
.A3(n_958),
.B(n_1154),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1093),
.A2(n_1002),
.B(n_1034),
.C(n_1031),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1093),
.A2(n_1098),
.B(n_963),
.Y(n_1376)
);

AOI31xp67_ASAP7_75t_L g1377 ( 
.A1(n_1114),
.A2(n_820),
.A3(n_1088),
.B(n_826),
.Y(n_1377)
);

BUFx4_ASAP7_75t_SL g1378 ( 
.A(n_1099),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_1115),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1093),
.A2(n_1098),
.B(n_963),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1107),
.A2(n_990),
.B(n_1101),
.Y(n_1381)
);

CKINVDCx11_ASAP7_75t_R g1382 ( 
.A(n_1104),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1162),
.A2(n_1002),
.B1(n_1199),
.B2(n_1034),
.Y(n_1383)
);

AOI221x1_ASAP7_75t_L g1384 ( 
.A1(n_1093),
.A2(n_1098),
.B1(n_741),
.B2(n_1102),
.C(n_1118),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1114),
.B(n_741),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1104),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1093),
.A2(n_1002),
.B(n_1034),
.C(n_741),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1107),
.A2(n_990),
.B(n_1101),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1141),
.A2(n_1016),
.B1(n_788),
.B2(n_1199),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1162),
.A2(n_1002),
.B1(n_1034),
.B2(n_595),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1107),
.A2(n_990),
.B(n_1101),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1143),
.B(n_792),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1093),
.A2(n_1002),
.B(n_1034),
.C(n_741),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1093),
.A2(n_746),
.B(n_734),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1118),
.A2(n_1088),
.B(n_1154),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_SL g1396 ( 
.A1(n_1143),
.A2(n_1002),
.B(n_1067),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1141),
.A2(n_1016),
.B1(n_788),
.B2(n_1199),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1115),
.B(n_906),
.Y(n_1398)
);

CKINVDCx11_ASAP7_75t_R g1399 ( 
.A(n_1382),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1374),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1256),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1249),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1290),
.A2(n_1357),
.B1(n_1313),
.B2(n_1304),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1357),
.A2(n_1313),
.B1(n_1291),
.B2(n_1302),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1300),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1343),
.B(n_1385),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1390),
.A2(n_1383),
.B1(n_1307),
.B2(n_1385),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1340),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1378),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1349),
.B(n_1387),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1398),
.B(n_1347),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1386),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1340),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1350),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1244),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1318),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1289),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1383),
.A2(n_1323),
.B1(n_1306),
.B2(n_1397),
.Y(n_1418)
);

INVx5_ASAP7_75t_L g1419 ( 
.A(n_1271),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1330),
.A2(n_1242),
.B1(n_1389),
.B2(n_1306),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_1326),
.Y(n_1421)
);

BUFx8_ASAP7_75t_L g1422 ( 
.A(n_1329),
.Y(n_1422)
);

BUFx2_ASAP7_75t_SL g1423 ( 
.A(n_1292),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1392),
.A2(n_1323),
.B1(n_1283),
.B2(n_1286),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1341),
.A2(n_1266),
.B1(n_1356),
.B2(n_1339),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1354),
.Y(n_1426)
);

AOI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1375),
.A2(n_1393),
.B(n_1371),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1353),
.A2(n_1272),
.B1(n_1345),
.B2(n_1281),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1319),
.Y(n_1429)
);

BUFx8_ASAP7_75t_SL g1430 ( 
.A(n_1398),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1281),
.A2(n_1301),
.B1(n_1346),
.B2(n_1380),
.Y(n_1431)
);

BUFx8_ASAP7_75t_L g1432 ( 
.A(n_1334),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1305),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1294),
.A2(n_1257),
.B1(n_1312),
.B2(n_1376),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1347),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1374),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1252),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1294),
.A2(n_1380),
.B1(n_1376),
.B2(n_1311),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1325),
.A2(n_1248),
.B1(n_1342),
.B2(n_1337),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1252),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1276),
.Y(n_1441)
);

CKINVDCx6p67_ASAP7_75t_R g1442 ( 
.A(n_1379),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1364),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1310),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1335),
.B(n_1338),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1332),
.A2(n_1270),
.B1(n_1316),
.B2(n_1337),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1374),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1288),
.A2(n_1327),
.B1(n_1314),
.B2(n_1263),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1255),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1379),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1305),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_SL g1452 ( 
.A(n_1305),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1373),
.Y(n_1453)
);

CKINVDCx6p67_ASAP7_75t_R g1454 ( 
.A(n_1373),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1373),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1355),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1321),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1267),
.A2(n_1342),
.B1(n_1320),
.B2(n_1348),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1331),
.A2(n_1394),
.B1(n_1258),
.B2(n_1279),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1320),
.A2(n_1284),
.B1(n_1317),
.B2(n_1282),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1384),
.A2(n_1277),
.B1(n_1280),
.B2(n_1246),
.Y(n_1461)
);

CKINVDCx6p67_ASAP7_75t_R g1462 ( 
.A(n_1321),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1351),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1278),
.A2(n_1269),
.B1(n_1363),
.B2(n_1245),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1262),
.B(n_1274),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1318),
.Y(n_1466)
);

CKINVDCx11_ASAP7_75t_R g1467 ( 
.A(n_1321),
.Y(n_1467)
);

BUFx2_ASAP7_75t_SL g1468 ( 
.A(n_1351),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1328),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1367),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1359),
.A2(n_1260),
.B1(n_1275),
.B2(n_1299),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1277),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1277),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1315),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1324),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1308),
.A2(n_1303),
.B1(n_1265),
.B2(n_1309),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1361),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1297),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1251),
.A2(n_1247),
.B1(n_1370),
.B2(n_1369),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1287),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1315),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1298),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1315),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1366),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1295),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1295),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1295),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1396),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1368),
.A2(n_1362),
.B1(n_1250),
.B2(n_1360),
.Y(n_1489)
);

INVx11_ASAP7_75t_L g1490 ( 
.A(n_1365),
.Y(n_1490)
);

BUFx12f_ASAP7_75t_L g1491 ( 
.A(n_1280),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1243),
.A2(n_1391),
.B1(n_1381),
.B2(n_1388),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1336),
.Y(n_1493)
);

BUFx4f_ASAP7_75t_SL g1494 ( 
.A(n_1377),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1360),
.Y(n_1495)
);

BUFx8_ASAP7_75t_SL g1496 ( 
.A(n_1372),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1322),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1336),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1336),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1395),
.A2(n_1261),
.B1(n_1254),
.B2(n_1322),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1293),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1358),
.A2(n_1293),
.B1(n_1253),
.B2(n_1344),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1264),
.A2(n_1296),
.B1(n_1285),
.B2(n_1358),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1268),
.A2(n_1259),
.B1(n_1352),
.B2(n_1358),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1273),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1273),
.A2(n_1002),
.B(n_1390),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1273),
.A2(n_1162),
.B1(n_1383),
.B2(n_1390),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1378),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1382),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1340),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1002),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1382),
.Y(n_1512)
);

BUFx10_ASAP7_75t_L g1513 ( 
.A(n_1326),
.Y(n_1513)
);

NAND2x1p5_ASAP7_75t_L g1514 ( 
.A(n_1327),
.B(n_1366),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1002),
.Y(n_1515)
);

CKINVDCx6p67_ASAP7_75t_R g1516 ( 
.A(n_1382),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1270),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1383),
.A2(n_1323),
.B1(n_1306),
.B2(n_1141),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1333),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1313),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1340),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1340),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1340),
.Y(n_1523)
);

BUFx2_ASAP7_75t_SL g1524 ( 
.A(n_1244),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1383),
.A2(n_1323),
.B1(n_1306),
.B2(n_1141),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1340),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1256),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1290),
.A2(n_1162),
.B1(n_1141),
.B2(n_1002),
.Y(n_1528)
);

OAI21xp33_ASAP7_75t_L g1529 ( 
.A1(n_1390),
.A2(n_1034),
.B(n_1002),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1256),
.Y(n_1530)
);

INVx8_ASAP7_75t_L g1531 ( 
.A(n_1256),
.Y(n_1531)
);

CKINVDCx11_ASAP7_75t_R g1532 ( 
.A(n_1382),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1313),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1313),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1390),
.A2(n_1383),
.B1(n_1199),
.B2(n_799),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1313),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1327),
.B(n_1366),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1256),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1313),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1382),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1382),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1313),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1382),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1290),
.A2(n_1162),
.B1(n_1141),
.B2(n_1002),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1300),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1383),
.A2(n_1323),
.B1(n_1306),
.B2(n_1141),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1390),
.A2(n_1162),
.B1(n_1383),
.B2(n_1002),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1382),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1249),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1474),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1481),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1400),
.B(n_1436),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1483),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1486),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_SL g1555 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1478),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1449),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1517),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1406),
.B(n_1407),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1419),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1485),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1500),
.A2(n_1465),
.B(n_1492),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1402),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1400),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1491),
.B(n_1445),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1404),
.B(n_1403),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1518),
.A2(n_1546),
.B1(n_1525),
.B2(n_1535),
.Y(n_1567)
);

BUFx4f_ASAP7_75t_L g1568 ( 
.A(n_1442),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1404),
.B(n_1403),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1503),
.A2(n_1465),
.B(n_1461),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1436),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1406),
.B(n_1529),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1447),
.B(n_1472),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1447),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1518),
.A2(n_1525),
.B1(n_1546),
.B2(n_1544),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1528),
.B(n_1544),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1473),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1487),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1487),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1493),
.B(n_1498),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1505),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1499),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1414),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1484),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1470),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1417),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1414),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1444),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1426),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1479),
.A2(n_1504),
.B(n_1489),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1426),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1495),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1446),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1418),
.A2(n_1420),
.B1(n_1425),
.B2(n_1439),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1506),
.B(n_1431),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1549),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1410),
.B(n_1461),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1495),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1504),
.A2(n_1477),
.B(n_1464),
.Y(n_1599)
);

OA21x2_ASAP7_75t_L g1600 ( 
.A1(n_1427),
.A2(n_1476),
.B(n_1471),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1514),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1430),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1427),
.A2(n_1460),
.B(n_1458),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1514),
.A2(n_1537),
.B(n_1459),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1528),
.A2(n_1418),
.B1(n_1520),
.B2(n_1542),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1496),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1537),
.A2(n_1428),
.B(n_1466),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1501),
.B(n_1416),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1488),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1435),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1501),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1494),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1416),
.B(n_1466),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1494),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1519),
.B(n_1522),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1522),
.B(n_1523),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1434),
.A2(n_1536),
.B(n_1533),
.Y(n_1617)
);

AOI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1469),
.A2(n_1490),
.B(n_1434),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1523),
.A2(n_1526),
.B(n_1539),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1419),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1497),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1507),
.B(n_1534),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1482),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1438),
.B(n_1515),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1422),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1405),
.Y(n_1626)
);

OAI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1511),
.A2(n_1515),
.B1(n_1547),
.B2(n_1424),
.C(n_1438),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1545),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1502),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1502),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1456),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1422),
.Y(n_1632)
);

INVx4_ASAP7_75t_L g1633 ( 
.A(n_1408),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1503),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1480),
.A2(n_1547),
.B1(n_1511),
.B2(n_1448),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1423),
.A2(n_1440),
.B1(n_1437),
.B2(n_1415),
.C(n_1524),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1475),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1408),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1411),
.B(n_1429),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1408),
.Y(n_1640)
);

OR2x6_ASAP7_75t_L g1641 ( 
.A(n_1413),
.B(n_1510),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1454),
.A2(n_1462),
.B(n_1457),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1433),
.Y(n_1643)
);

BUFx2_ASAP7_75t_SL g1644 ( 
.A(n_1421),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1413),
.A2(n_1521),
.B(n_1510),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1530),
.Y(n_1646)
);

OA21x2_ASAP7_75t_L g1647 ( 
.A1(n_1457),
.A2(n_1468),
.B(n_1455),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1538),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1521),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1538),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1450),
.A2(n_1531),
.B(n_1452),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1401),
.B(n_1453),
.Y(n_1652)
);

AOI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1451),
.A2(n_1455),
.B(n_1450),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1463),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1463),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1463),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_SL g1657 ( 
.A1(n_1421),
.A2(n_1513),
.B1(n_1543),
.B2(n_1541),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1531),
.A2(n_1508),
.B(n_1409),
.C(n_1452),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1527),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1467),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1432),
.A2(n_1516),
.B(n_1412),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1432),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1617),
.A2(n_1509),
.B(n_1512),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1583),
.B(n_1548),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1575),
.A2(n_1399),
.B(n_1532),
.C(n_1540),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1605),
.A2(n_1627),
.B(n_1622),
.C(n_1576),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1564),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1565),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1621),
.B(n_1565),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1623),
.B(n_1631),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1622),
.A2(n_1624),
.B(n_1635),
.C(n_1569),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1567),
.A2(n_1594),
.B1(n_1569),
.B2(n_1566),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1604),
.B(n_1565),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1565),
.B(n_1557),
.Y(n_1674)
);

AO21x2_ASAP7_75t_L g1675 ( 
.A1(n_1562),
.A2(n_1614),
.B(n_1612),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1566),
.A2(n_1624),
.B1(n_1595),
.B2(n_1559),
.C(n_1634),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1644),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1593),
.B(n_1610),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1660),
.Y(n_1679)
);

AO21x1_ASAP7_75t_L g1680 ( 
.A1(n_1572),
.A2(n_1597),
.B(n_1587),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1583),
.B(n_1587),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1555),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1595),
.A2(n_1636),
.B(n_1604),
.C(n_1568),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1600),
.A2(n_1606),
.B1(n_1609),
.B2(n_1637),
.Y(n_1684)
);

AO32x2_ASAP7_75t_L g1685 ( 
.A1(n_1633),
.A2(n_1570),
.A3(n_1629),
.B1(n_1630),
.B2(n_1573),
.Y(n_1685)
);

NOR2x1_ASAP7_75t_SL g1686 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1647),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1600),
.A2(n_1562),
.B(n_1570),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1599),
.A2(n_1590),
.B(n_1634),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1607),
.B(n_1645),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1586),
.B(n_1588),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1600),
.A2(n_1603),
.B(n_1618),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1600),
.A2(n_1603),
.B(n_1618),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1603),
.A2(n_1590),
.B(n_1619),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1639),
.B(n_1637),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1596),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1573),
.B(n_1552),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_SL g1698 ( 
.A(n_1641),
.B(n_1653),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1603),
.A2(n_1619),
.B(n_1599),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1657),
.A2(n_1660),
.B1(n_1662),
.B2(n_1625),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1552),
.B(n_1563),
.Y(n_1701)
);

AO32x2_ASAP7_75t_L g1702 ( 
.A1(n_1633),
.A2(n_1629),
.A3(n_1630),
.B1(n_1580),
.B2(n_1560),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1607),
.A2(n_1554),
.B(n_1551),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1584),
.B(n_1601),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_SL g1705 ( 
.A1(n_1658),
.A2(n_1662),
.B(n_1609),
.C(n_1614),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1615),
.B(n_1626),
.Y(n_1706)
);

AOI211xp5_ASAP7_75t_L g1707 ( 
.A1(n_1609),
.A2(n_1612),
.B(n_1558),
.C(n_1628),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1644),
.A2(n_1616),
.B1(n_1640),
.B2(n_1638),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1592),
.B(n_1598),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1592),
.B(n_1598),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1647),
.A2(n_1611),
.B(n_1608),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1554),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1660),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1615),
.A2(n_1653),
.B(n_1651),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1577),
.B(n_1556),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1568),
.A2(n_1651),
.B(n_1601),
.C(n_1649),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_R g1717 ( 
.A(n_1660),
.B(n_1602),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1550),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1660),
.B2(n_1574),
.C(n_1571),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1602),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1625),
.A2(n_1632),
.B1(n_1568),
.B2(n_1641),
.Y(n_1721)
);

AO22x2_ASAP7_75t_L g1722 ( 
.A1(n_1553),
.A2(n_1579),
.B1(n_1578),
.B2(n_1581),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1638),
.B(n_1649),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1696),
.B(n_1581),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1663),
.A2(n_1649),
.B(n_1640),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1686),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1667),
.Y(n_1727)
);

OAI22x1_ASAP7_75t_SL g1728 ( 
.A1(n_1720),
.A2(n_1661),
.B1(n_1632),
.B2(n_1640),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1697),
.B(n_1582),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1683),
.B(n_1647),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1702),
.B(n_1580),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1667),
.Y(n_1732)
);

NOR2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1713),
.B(n_1638),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1702),
.B(n_1561),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1722),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1722),
.Y(n_1737)
);

BUFx12f_ASAP7_75t_L g1738 ( 
.A(n_1677),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1722),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1685),
.B(n_1561),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1685),
.B(n_1611),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1712),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_SL g1743 ( 
.A1(n_1672),
.A2(n_1620),
.B1(n_1661),
.B2(n_1560),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1685),
.B(n_1585),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1666),
.A2(n_1620),
.B1(n_1560),
.B2(n_1654),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1672),
.A2(n_1654),
.B1(n_1656),
.B2(n_1613),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1690),
.Y(n_1747)
);

OAI222xp33_ASAP7_75t_L g1748 ( 
.A1(n_1721),
.A2(n_1656),
.B1(n_1643),
.B2(n_1650),
.C1(n_1648),
.C2(n_1646),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1664),
.B(n_1655),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1690),
.B(n_1613),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1703),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1673),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1663),
.A2(n_1655),
.B1(n_1613),
.B2(n_1659),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1690),
.B(n_1643),
.Y(n_1755)
);

BUFx8_ASAP7_75t_SL g1756 ( 
.A(n_1679),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1718),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1718),
.Y(n_1758)
);

INVxp67_ASAP7_75t_SL g1759 ( 
.A(n_1710),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1664),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1681),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1701),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1681),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1704),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1709),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1736),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1727),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1727),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1749),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1751),
.B(n_1698),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1731),
.B(n_1734),
.Y(n_1771)
);

NOR3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1745),
.B(n_1700),
.C(n_1721),
.Y(n_1772)
);

OAI33xp33_ASAP7_75t_L g1773 ( 
.A1(n_1736),
.A2(n_1691),
.A3(n_1715),
.B1(n_1668),
.B2(n_1669),
.B3(n_1674),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.B(n_1687),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1732),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1751),
.B(n_1755),
.Y(n_1776)
);

OAI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1752),
.A2(n_1688),
.B(n_1749),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1732),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1743),
.A2(n_1676),
.B1(n_1665),
.B2(n_1684),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1745),
.B(n_1707),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1751),
.B(n_1714),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1762),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1734),
.B(n_1687),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1756),
.Y(n_1785)
);

AND2x6_ASAP7_75t_L g1786 ( 
.A(n_1730),
.B(n_1751),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1730),
.B(n_1676),
.C(n_1694),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1738),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1725),
.A2(n_1671),
.B1(n_1746),
.B2(n_1754),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1738),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_L g1791 ( 
.A(n_1725),
.B(n_1694),
.C(n_1699),
.Y(n_1791)
);

OAI33xp33_ASAP7_75t_L g1792 ( 
.A1(n_1737),
.A2(n_1739),
.A3(n_1760),
.B1(n_1758),
.B2(n_1757),
.B3(n_1724),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_L g1793 ( 
.A(n_1746),
.B(n_1699),
.C(n_1688),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1678),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1739),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1729),
.B(n_1689),
.Y(n_1796)
);

NOR2xp67_ASAP7_75t_L g1797 ( 
.A(n_1738),
.B(n_1711),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1757),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1728),
.A2(n_1693),
.B1(n_1692),
.B2(n_1680),
.C(n_1705),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1758),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1747),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1765),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1761),
.B(n_1706),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1755),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1764),
.B(n_1689),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1750),
.A2(n_1665),
.B1(n_1716),
.B2(n_1708),
.C(n_1682),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1742),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1764),
.B(n_1675),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1765),
.Y(n_1809)
);

OR2x6_ASAP7_75t_L g1810 ( 
.A(n_1753),
.B(n_1747),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1733),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1764),
.B(n_1675),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1774),
.B(n_1744),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1796),
.B(n_1749),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1774),
.B(n_1805),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1805),
.B(n_1744),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1801),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1795),
.B(n_1761),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1801),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1769),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1771),
.B(n_1741),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1785),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1766),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1741),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1796),
.B(n_1769),
.Y(n_1825)
);

NOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1787),
.B(n_1728),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1795),
.B(n_1763),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1804),
.B(n_1783),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1777),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1786),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1784),
.B(n_1752),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1777),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1770),
.B(n_1753),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1786),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1804),
.B(n_1740),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1808),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1770),
.B(n_1753),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1740),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1812),
.B(n_1776),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1812),
.B(n_1735),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1789),
.A2(n_1692),
.B1(n_1693),
.B2(n_1670),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1770),
.B(n_1753),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1767),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1776),
.B(n_1735),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1767),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1780),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1768),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1776),
.B(n_1752),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1768),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1775),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1775),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1778),
.Y(n_1852)
);

NOR2xp67_ASAP7_75t_L g1853 ( 
.A(n_1822),
.B(n_1811),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1823),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1822),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1823),
.Y(n_1856)
);

OAI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1826),
.A2(n_1799),
.B(n_1779),
.C(n_1793),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1835),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1826),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1817),
.B(n_1802),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1844),
.B(n_1833),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1846),
.B(n_1782),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1845),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1845),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1845),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1847),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1847),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1817),
.B(n_1809),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1822),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1846),
.B(n_1794),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1841),
.B(n_1800),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1847),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1849),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1822),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1835),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1822),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1833),
.B(n_1810),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1849),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1822),
.B(n_1788),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1849),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1826),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1817),
.B(n_1778),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1841),
.B(n_1800),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1819),
.B(n_1798),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1835),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1843),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1819),
.B(n_1791),
.Y(n_1891)
);

AND2x4_ASAP7_75t_SL g1892 ( 
.A(n_1822),
.B(n_1772),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1843),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1818),
.B(n_1807),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1831),
.B(n_1806),
.C(n_1797),
.Y(n_1896)
);

NAND4xp25_ASAP7_75t_L g1897 ( 
.A(n_1830),
.B(n_1790),
.C(n_1695),
.D(n_1719),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1818),
.B(n_1811),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1862),
.B(n_1833),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1865),
.Y(n_1900)
);

AND3x2_ASAP7_75t_L g1901 ( 
.A(n_1860),
.B(n_1834),
.C(n_1830),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1865),
.Y(n_1902)
);

AND2x4_ASAP7_75t_SL g1903 ( 
.A(n_1881),
.B(n_1679),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1874),
.B(n_1821),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1885),
.B(n_1717),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1868),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1887),
.B(n_1821),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1862),
.B(n_1833),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1873),
.B(n_1821),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1868),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1870),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1857),
.B(n_1839),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1863),
.B(n_1821),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1892),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1870),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1872),
.B(n_1733),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1858),
.B(n_1833),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1859),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1876),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1858),
.B(n_1869),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1861),
.B(n_1818),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1869),
.B(n_1833),
.Y(n_1922)
);

AND2x4_ASAP7_75t_SL g1923 ( 
.A(n_1881),
.B(n_1679),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1892),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1883),
.B(n_1839),
.Y(n_1925)
);

NAND2xp33_ASAP7_75t_R g1926 ( 
.A(n_1891),
.B(n_1830),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1897),
.B(n_1839),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1854),
.B(n_1839),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1853),
.B(n_1833),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1876),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1884),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1856),
.B(n_1815),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1861),
.B(n_1827),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1891),
.B(n_1815),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1898),
.B(n_1815),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1912),
.B(n_1855),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1927),
.A2(n_1896),
.B(n_1877),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1914),
.Y(n_1938)
);

OAI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1905),
.A2(n_1834),
.B1(n_1877),
.B2(n_1872),
.C(n_1880),
.Y(n_1939)
);

AOI221x1_ASAP7_75t_L g1940 ( 
.A1(n_1934),
.A2(n_1872),
.B1(n_1880),
.B2(n_1888),
.C(n_1894),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1899),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1929),
.B(n_1880),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1900),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1902),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1924),
.A2(n_1773),
.B1(n_1879),
.B2(n_1792),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1929),
.B(n_1785),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1920),
.B(n_1917),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1929),
.A2(n_1790),
.B1(n_1834),
.B2(n_1786),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1920),
.A2(n_1879),
.B1(n_1786),
.B2(n_1842),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1906),
.Y(n_1950)
);

AOI21xp33_ASAP7_75t_L g1951 ( 
.A1(n_1926),
.A2(n_1871),
.B(n_1886),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1910),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1917),
.B(n_1871),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1926),
.A2(n_1786),
.B1(n_1837),
.B2(n_1842),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1903),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1899),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1922),
.B(n_1837),
.Y(n_1957)
);

NAND2x1_ASAP7_75t_L g1958 ( 
.A(n_1908),
.B(n_1786),
.Y(n_1958)
);

OAI211xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1925),
.A2(n_1928),
.B(n_1907),
.C(n_1904),
.Y(n_1959)
);

OAI322xp33_ASAP7_75t_L g1960 ( 
.A1(n_1932),
.A2(n_1878),
.A3(n_1867),
.B1(n_1859),
.B2(n_1889),
.C1(n_1886),
.C2(n_1884),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1922),
.B(n_1824),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1935),
.A2(n_1867),
.B1(n_1878),
.B2(n_1889),
.C(n_1875),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1943),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1944),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1937),
.A2(n_1901),
.B1(n_1913),
.B2(n_1909),
.Y(n_1965)
);

OAI21xp33_ASAP7_75t_SL g1966 ( 
.A1(n_1951),
.A2(n_1908),
.B(n_1921),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1938),
.B(n_1947),
.Y(n_1967)
);

NAND4xp25_ASAP7_75t_SL g1968 ( 
.A(n_1945),
.B(n_1933),
.C(n_1921),
.D(n_1901),
.Y(n_1968)
);

NOR2x1_ASAP7_75t_R g1969 ( 
.A(n_1946),
.B(n_1726),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1945),
.A2(n_1931),
.B1(n_1930),
.B2(n_1911),
.C(n_1919),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1950),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1952),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1955),
.B(n_1903),
.Y(n_1973)
);

O2A1O1Ixp33_ASAP7_75t_SL g1974 ( 
.A1(n_1946),
.A2(n_1933),
.B(n_1915),
.C(n_1918),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1936),
.B(n_1923),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1954),
.A2(n_1916),
.B1(n_1923),
.B2(n_1842),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1953),
.Y(n_1977)
);

OAI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1959),
.A2(n_1916),
.B(n_1918),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1939),
.A2(n_1866),
.B1(n_1864),
.B2(n_1882),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1949),
.A2(n_1837),
.B1(n_1842),
.B2(n_1781),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1941),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1941),
.B(n_1828),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1942),
.A2(n_1837),
.B(n_1842),
.Y(n_1983)
);

NAND4xp25_ASAP7_75t_L g1984 ( 
.A(n_1965),
.B(n_1967),
.C(n_1970),
.D(n_1977),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1968),
.A2(n_1940),
.B(n_1942),
.Y(n_1985)
);

AND2x2_ASAP7_75t_SL g1986 ( 
.A(n_1965),
.B(n_1956),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1981),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1963),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1974),
.A2(n_1948),
.B(n_1960),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1973),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1964),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1971),
.B(n_1956),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1982),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1972),
.B(n_1962),
.Y(n_1994)
);

NAND4xp25_ASAP7_75t_L g1995 ( 
.A(n_1975),
.B(n_1957),
.C(n_1961),
.D(n_1837),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1978),
.B(n_1957),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1966),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1984),
.B(n_1979),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_L g1999 ( 
.A(n_1985),
.B(n_1989),
.C(n_1997),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1996),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1990),
.B(n_1969),
.Y(n_2001)
);

AND3x2_ASAP7_75t_L g2002 ( 
.A(n_1985),
.B(n_1837),
.C(n_1842),
.Y(n_2002)
);

OAI21xp33_ASAP7_75t_SL g2003 ( 
.A1(n_1986),
.A2(n_1979),
.B(n_1983),
.Y(n_2003)
);

NOR3xp33_ASAP7_75t_L g2004 ( 
.A(n_1994),
.B(n_1995),
.C(n_1992),
.Y(n_2004)
);

OA211x2_ASAP7_75t_L g2005 ( 
.A1(n_1994),
.A2(n_1958),
.B(n_1976),
.C(n_1827),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1992),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1987),
.Y(n_2007)
);

NAND4xp75_ASAP7_75t_L g2008 ( 
.A(n_1988),
.B(n_1642),
.C(n_1980),
.D(n_1848),
.Y(n_2008)
);

NOR2xp67_ASAP7_75t_L g2009 ( 
.A(n_2006),
.B(n_1991),
.Y(n_2009)
);

OAI211xp5_ASAP7_75t_SL g2010 ( 
.A1(n_1998),
.A2(n_1993),
.B(n_1893),
.C(n_1890),
.Y(n_2010)
);

OAI32xp33_ASAP7_75t_L g2011 ( 
.A1(n_2003),
.A2(n_1836),
.A3(n_1831),
.B1(n_1829),
.B2(n_1895),
.Y(n_2011)
);

AOI211xp5_ASAP7_75t_L g2012 ( 
.A1(n_1999),
.A2(n_1837),
.B(n_1842),
.C(n_1748),
.Y(n_2012)
);

AOI322xp5_ASAP7_75t_L g2013 ( 
.A1(n_2004),
.A2(n_1824),
.A3(n_1816),
.B1(n_1838),
.B2(n_1840),
.C1(n_1813),
.C2(n_1815),
.Y(n_2013)
);

AOI21xp33_ASAP7_75t_SL g2014 ( 
.A1(n_2001),
.A2(n_1642),
.B(n_1831),
.Y(n_2014)
);

OAI221xp5_ASAP7_75t_SL g2015 ( 
.A1(n_2013),
.A2(n_2000),
.B1(n_2007),
.B2(n_2005),
.C(n_2002),
.Y(n_2015)
);

O2A1O1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_2011),
.A2(n_2008),
.B(n_1829),
.C(n_1831),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_2009),
.A2(n_1895),
.B(n_1814),
.Y(n_2017)
);

NOR3xp33_ASAP7_75t_SL g2018 ( 
.A(n_2010),
.B(n_1748),
.C(n_1723),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_2014),
.A2(n_1829),
.B1(n_1832),
.B2(n_1836),
.C(n_1848),
.Y(n_2019)
);

AOI21xp33_ASAP7_75t_L g2020 ( 
.A1(n_2012),
.A2(n_1829),
.B(n_1832),
.Y(n_2020)
);

AOI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_2011),
.A2(n_1829),
.B1(n_1832),
.B2(n_1836),
.C(n_1848),
.Y(n_2021)
);

XNOR2xp5_ASAP7_75t_L g2022 ( 
.A(n_2018),
.B(n_2017),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2015),
.Y(n_2023)
);

XNOR2xp5_ASAP7_75t_L g2024 ( 
.A(n_2019),
.B(n_1642),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_2021),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2016),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_2020),
.B(n_1836),
.Y(n_2027)
);

OAI211xp5_ASAP7_75t_SL g2028 ( 
.A1(n_2023),
.A2(n_1836),
.B(n_1832),
.C(n_1814),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_2026),
.B(n_1848),
.Y(n_2029)
);

NOR2x1_ASAP7_75t_L g2030 ( 
.A(n_2022),
.B(n_1850),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_SL g2031 ( 
.A1(n_2029),
.A2(n_2025),
.B1(n_2024),
.B2(n_2027),
.Y(n_2031)
);

AOI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_2031),
.A2(n_2025),
.B1(n_2028),
.B2(n_2030),
.Y(n_2032)
);

INVxp67_ASAP7_75t_SL g2033 ( 
.A(n_2032),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_2032),
.A2(n_1825),
.B1(n_1814),
.B2(n_1850),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_2033),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2034),
.B(n_1850),
.Y(n_2036)
);

AOI221xp5_ASAP7_75t_L g2037 ( 
.A1(n_2035),
.A2(n_1851),
.B1(n_1850),
.B2(n_1852),
.C(n_1843),
.Y(n_2037)
);

NAND2x1p5_ASAP7_75t_L g2038 ( 
.A(n_2036),
.B(n_1642),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_2038),
.A2(n_1814),
.B(n_1825),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2039),
.B(n_2037),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2040),
.A2(n_1851),
.B1(n_1850),
.B2(n_1852),
.C(n_1843),
.Y(n_2041)
);

OAI221xp5_ASAP7_75t_L g2042 ( 
.A1(n_2041),
.A2(n_1851),
.B1(n_1825),
.B2(n_1852),
.C(n_1820),
.Y(n_2042)
);

AOI211xp5_ASAP7_75t_L g2043 ( 
.A1(n_2042),
.A2(n_1620),
.B(n_1825),
.C(n_1652),
.Y(n_2043)
);


endmodule