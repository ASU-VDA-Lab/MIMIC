module fake_jpeg_24938_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_25),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_14),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_36),
.C(n_23),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_12),
.C(n_19),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_11),
.B(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_11),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_23),
.B1(n_19),
.B2(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_22),
.B1(n_20),
.B2(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_40),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_29),
.B(n_21),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_17),
.B1(n_3),
.B2(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_50),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_55),
.B1(n_41),
.B2(n_7),
.Y(n_59)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_30),
.B1(n_31),
.B2(n_45),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_6),
.B1(n_8),
.B2(n_51),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_57),
.B(n_35),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_53),
.C(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_57),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_41),
.B(n_7),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_61),
.B(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_65),
.B1(n_62),
.B2(n_56),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_62),
.C(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_68),
.B1(n_69),
.B2(n_55),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_55),
.Y(n_72)
);


endmodule