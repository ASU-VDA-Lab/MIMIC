module fake_netlist_6_402_n_2277 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2277);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2277;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_1207;
wire n_811;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_1159;
wire n_276;
wire n_995;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_181),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_215),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_109),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_71),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_93),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_19),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_114),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_144),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_178),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_0),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_69),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_192),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_38),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_84),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_4),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_199),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_161),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_43),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_54),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_79),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_171),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_131),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_182),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_190),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_72),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_43),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_75),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_166),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_65),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_217),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_222),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_83),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_67),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_113),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_216),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_158),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_65),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_103),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_142),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_194),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_116),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_115),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_90),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_100),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_107),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_80),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_25),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_17),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_221),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_59),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_48),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_177),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_207),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_126),
.Y(n_302)
);

BUFx8_ASAP7_75t_SL g303 ( 
.A(n_140),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_130),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_136),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_108),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

INVxp33_ASAP7_75t_SL g310 ( 
.A(n_42),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_0),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_77),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_48),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_118),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_204),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_111),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_165),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_155),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_185),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_72),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_176),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_97),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_153),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_83),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_87),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_68),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_25),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_4),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_99),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_39),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_187),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_120),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_170),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_75),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_157),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_41),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_30),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_122),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_213),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_89),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_163),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_196),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_51),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_180),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_52),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_22),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_223),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_127),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_134),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_63),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_9),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_101),
.Y(n_354)
);

BUFx2_ASAP7_75t_SL g355 ( 
.A(n_86),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_156),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_74),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_102),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_132),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_68),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_34),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_208),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_14),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_145),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_179),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_138),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_174),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_149),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_31),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_104),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_148),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_191),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_86),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_82),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_21),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_141),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_96),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_52),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_92),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_91),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_64),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_64),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_188),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_226),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_44),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_123),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_201),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_11),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_77),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_14),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_76),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_112),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_6),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_49),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_95),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_15),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_79),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_27),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_2),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_98),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_227),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_13),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_186),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_26),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_119),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_81),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_71),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_33),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_88),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_42),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_76),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_169),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_128),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_220),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_80),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_35),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_41),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_159),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_73),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_147),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_164),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_69),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_11),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_45),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_27),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_198),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_51),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_10),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_1),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_32),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_124),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_110),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_209),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_167),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_151),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_57),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_58),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_50),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_150),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_211),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_62),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_78),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_212),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_50),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_129),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_18),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_15),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_399),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_394),
.B(n_1),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_394),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_394),
.B(n_3),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_233),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g456 ( 
.A(n_233),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_394),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_295),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_295),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_384),
.B(n_3),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_311),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_311),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_303),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_228),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_229),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_230),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_245),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_231),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_236),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_251),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_251),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_237),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_R g480 ( 
.A(n_384),
.B(n_5),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_239),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_364),
.B(n_6),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_323),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_244),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_261),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_312),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_261),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_240),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_246),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_242),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_288),
.B(n_7),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_269),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_249),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_245),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_288),
.B(n_7),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_255),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_263),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_252),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_256),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_250),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_262),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_265),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_263),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_269),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_267),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_271),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_268),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_287),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_370),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_306),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_276),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_280),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_281),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_322),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_282),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_291),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_292),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_297),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_305),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_307),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_250),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_346),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_271),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_309),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_279),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_279),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_331),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_285),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_331),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_314),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_361),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_285),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_304),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_354),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_361),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_316),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_318),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_304),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_327),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_393),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_320),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_324),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_326),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_406),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_419),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_428),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_293),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_327),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_434),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_335),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_253),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_253),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_277),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_332),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_335),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_352),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_277),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_352),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_334),
.Y(n_559)
);

INVx4_ASAP7_75t_R g560 ( 
.A(n_293),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_337),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_342),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_357),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_349),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_357),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_374),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_350),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_374),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_364),
.B(n_8),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_482),
.B(n_234),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_490),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_463),
.A2(n_428),
.B1(n_437),
.B2(n_397),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_482),
.B(n_340),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_470),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_490),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_477),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_490),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_319),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_477),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_490),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_478),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_491),
.B(n_319),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_478),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_569),
.B(n_340),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_259),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_494),
.B(n_294),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_497),
.B(n_503),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_495),
.B(n_351),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_449),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_497),
.B(n_264),
.Y(n_594)
);

CKINVDCx14_ASAP7_75t_R g595 ( 
.A(n_551),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_485),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_552),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_310),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_452),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_452),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_503),
.B(n_454),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_487),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_557),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_457),
.B(n_264),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_487),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_458),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_459),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_460),
.B(n_254),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_461),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_461),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_492),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_462),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_451),
.B(n_254),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_504),
.B(n_360),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_462),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_504),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_506),
.B(n_363),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_506),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_523),
.B(n_366),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_523),
.B(n_367),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_526),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_526),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_528),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_560),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_465),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_465),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_532),
.B(n_259),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_469),
.Y(n_640)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_488),
.B(n_232),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_533),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_533),
.B(n_301),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_469),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_494),
.A2(n_235),
.B1(n_258),
.B2(n_407),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_521),
.B(n_286),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_538),
.B(n_301),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_471),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_538),
.B(n_369),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_539),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_471),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_539),
.B(n_343),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_467),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_474),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_548),
.B(n_371),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_548),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_500),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_474),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_550),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_550),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_555),
.B(n_266),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_466),
.B(n_372),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_521),
.B(n_294),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_570),
.B(n_468),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_602),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_593),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_646),
.B(n_355),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_570),
.B(n_472),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_573),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_635),
.B(n_475),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_570),
.B(n_592),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_622),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_598),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_598),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_593),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_602),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_602),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_635),
.B(n_476),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_592),
.B(n_479),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_635),
.B(n_481),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_598),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_607),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_585),
.B(n_484),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_604),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_604),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_620),
.A2(n_483),
.B1(n_299),
.B2(n_450),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_635),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_585),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_657),
.Y(n_691)
);

INVx8_ASAP7_75t_L g692 ( 
.A(n_635),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_572),
.B(n_480),
.C(n_489),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_604),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_635),
.B(n_493),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_611),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_622),
.B(n_498),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_598),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_607),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_573),
.B(n_555),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_600),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_573),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_622),
.B(n_499),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_657),
.B(n_527),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_598),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_611),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_587),
.B(n_556),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_598),
.Y(n_708)
);

NOR2x1p5_ASAP7_75t_L g709 ( 
.A(n_653),
.B(n_389),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_635),
.B(n_501),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_598),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_611),
.Y(n_712)
);

XNOR2xp5_ASAP7_75t_L g713 ( 
.A(n_572),
.B(n_496),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_635),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_605),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_605),
.Y(n_716)
);

AOI21x1_ASAP7_75t_L g717 ( 
.A1(n_614),
.A2(n_274),
.B(n_266),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_587),
.B(n_556),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_598),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_622),
.B(n_502),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_587),
.B(n_558),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_664),
.A2(n_529),
.B1(n_546),
.B2(n_527),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_580),
.B(n_505),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_605),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_601),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_605),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_590),
.B(n_507),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_605),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_591),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_595),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_589),
.B(n_512),
.C(n_511),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_658),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_646),
.A2(n_515),
.B1(n_516),
.B2(n_513),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_591),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_663),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_622),
.B(n_517),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_600),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_622),
.B(n_518),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_608),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_662),
.B(n_558),
.Y(n_741)
);

INVx5_ASAP7_75t_L g742 ( 
.A(n_601),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_590),
.B(n_519),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_601),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_608),
.Y(n_745)
);

BUFx8_ASAP7_75t_SL g746 ( 
.A(n_597),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_664),
.B(n_520),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_608),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_620),
.B(n_524),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_608),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_601),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_607),
.B(n_242),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_610),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_645),
.B(n_355),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_610),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_620),
.A2(n_299),
.B1(n_535),
.B2(n_531),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_620),
.B(n_530),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_663),
.B(n_536),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_580),
.B(n_537),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_662),
.B(n_594),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_589),
.B(n_542),
.C(n_541),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_621),
.B(n_543),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_591),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_614),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_641),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_601),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_620),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_641),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_621),
.B(n_554),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_610),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_610),
.Y(n_771)
);

INVx6_ASAP7_75t_L g772 ( 
.A(n_601),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_601),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_658),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_613),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_613),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_643),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_613),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_613),
.Y(n_779)
);

AND2x6_ASAP7_75t_L g780 ( 
.A(n_614),
.B(n_343),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_625),
.B(n_559),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_614),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_641),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_614),
.Y(n_784)
);

BUFx10_ASAP7_75t_L g785 ( 
.A(n_643),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_595),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_601),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_643),
.A2(n_389),
.B1(n_391),
.B2(n_390),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_616),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_612),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_612),
.Y(n_791)
);

AND2x2_ASAP7_75t_SL g792 ( 
.A(n_639),
.B(n_344),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_625),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_612),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_629),
.B(n_561),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_662),
.B(n_274),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_612),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_597),
.Y(n_798)
);

NOR2x1p5_ASAP7_75t_L g799 ( 
.A(n_629),
.B(n_390),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_594),
.B(n_563),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_616),
.Y(n_801)
);

AND2x2_ASAP7_75t_SL g802 ( 
.A(n_639),
.B(n_344),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_643),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_597),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_630),
.B(n_562),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_612),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_645),
.A2(n_567),
.B1(n_564),
.B2(n_546),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_612),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_612),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_594),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_612),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_643),
.B(n_283),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_577),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_630),
.B(n_391),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_577),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_SL g816 ( 
.A(n_649),
.B(n_238),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_649),
.B(n_655),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_616),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_655),
.B(n_529),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_582),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_616),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_617),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_730),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_810),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_793),
.A2(n_510),
.B1(n_514),
.B2(n_508),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_666),
.A2(n_398),
.B1(n_408),
.B2(n_392),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_793),
.A2(n_534),
.B1(n_540),
.B2(n_522),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_798),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_685),
.B(n_684),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_762),
.A2(n_545),
.B1(n_549),
.B2(n_544),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_672),
.B(n_486),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_690),
.B(n_767),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_798),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_667),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_684),
.B(n_623),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_723),
.B(n_509),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_699),
.B(n_623),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_749),
.B(n_247),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_730),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_699),
.B(n_623),
.Y(n_840)
);

AO221x1_ASAP7_75t_L g841 ( 
.A1(n_668),
.A2(n_257),
.B1(n_444),
.B2(n_242),
.C(n_392),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_673),
.B(n_623),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_795),
.B(n_623),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_767),
.B(n_242),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_704),
.B(n_606),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_670),
.B(n_455),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_760),
.B(n_627),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_757),
.B(n_336),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_681),
.B(n_456),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_736),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_735),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_817),
.A2(n_702),
.B1(n_670),
.B2(n_816),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_767),
.B(n_242),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_760),
.B(n_627),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_666),
.A2(n_408),
.B1(n_412),
.B2(n_398),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_810),
.B(n_627),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_702),
.B(n_525),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_735),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_691),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_678),
.B(n_627),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_678),
.B(n_679),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_679),
.B(n_627),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_698),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_763),
.B(n_640),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_763),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_697),
.B(n_444),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_817),
.B(n_640),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_764),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_703),
.B(n_444),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_674),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_720),
.B(n_444),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_817),
.A2(n_377),
.B1(n_378),
.B2(n_373),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_817),
.B(n_640),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_693),
.B(n_756),
.C(n_688),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_733),
.B(n_606),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_769),
.B(n_241),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_737),
.B(n_640),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_781),
.B(n_243),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_739),
.B(n_640),
.Y(n_879)
);

NOR2x1p5_ASAP7_75t_L g880 ( 
.A(n_736),
.B(n_248),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_792),
.B(n_647),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_805),
.B(n_659),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_792),
.B(n_659),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_764),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_733),
.Y(n_885)
);

OAI221xp5_ASAP7_75t_L g886 ( 
.A1(n_788),
.A2(n_412),
.B1(n_420),
.B2(n_425),
.C(n_426),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_813),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_799),
.Y(n_888)
);

NAND3xp33_ASAP7_75t_L g889 ( 
.A(n_734),
.B(n_599),
.C(n_270),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_802),
.B(n_647),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_813),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_802),
.B(n_659),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_665),
.B(n_260),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_780),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_815),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_700),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_669),
.B(n_759),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_741),
.B(n_659),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_668),
.A2(n_606),
.B1(n_413),
.B2(n_286),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_741),
.B(n_815),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_820),
.B(n_659),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_820),
.B(n_647),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_782),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_777),
.B(n_647),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_774),
.B(n_420),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_800),
.B(n_647),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_777),
.B(n_652),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_704),
.B(n_599),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_819),
.B(n_272),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_800),
.B(n_784),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_784),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_777),
.B(n_652),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_700),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_796),
.B(n_652),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_677),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_796),
.B(n_652),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_785),
.B(n_652),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_814),
.B(n_273),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_668),
.A2(n_381),
.B1(n_385),
.B2(n_380),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_701),
.Y(n_920)
);

BUFx6f_ASAP7_75t_SL g921 ( 
.A(n_754),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_796),
.A2(n_426),
.B1(n_429),
.B2(n_425),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_814),
.B(n_275),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_707),
.B(n_637),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_774),
.B(n_599),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_707),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_807),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_668),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_814),
.B(n_582),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_701),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_814),
.A2(n_283),
.B1(n_284),
.B2(n_289),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_799),
.A2(n_387),
.B1(n_388),
.B2(n_401),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_718),
.B(n_637),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_718),
.B(n_637),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_721),
.A2(n_447),
.B(n_429),
.C(n_290),
.Y(n_935)
);

NOR2x1p5_ASAP7_75t_L g936 ( 
.A(n_732),
.B(n_278),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_721),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_812),
.B(n_284),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_715),
.B(n_716),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_716),
.B(n_637),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_724),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_709),
.A2(n_446),
.B1(n_436),
.B2(n_433),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_724),
.B(n_637),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_L g944 ( 
.A(n_780),
.B(n_402),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_722),
.B(n_584),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_785),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_709),
.B(n_584),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_726),
.B(n_637),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_803),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_803),
.B(n_404),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_726),
.B(n_410),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_729),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_728),
.B(n_637),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_728),
.B(n_637),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_812),
.B(n_415),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_761),
.B(n_296),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_812),
.B(n_790),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_772),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_772),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_754),
.B(n_447),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_686),
.Y(n_961)
);

AO22x2_ASAP7_75t_L g962 ( 
.A1(n_727),
.A2(n_289),
.B1(n_290),
.B2(n_300),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_698),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_743),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_686),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_687),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_738),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_752),
.A2(n_661),
.B(n_660),
.C(n_656),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_L g969 ( 
.A(n_747),
.B(n_308),
.C(n_298),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_780),
.A2(n_341),
.B1(n_441),
.B2(n_440),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_790),
.B(n_644),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_797),
.B(n_421),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_797),
.B(n_422),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_806),
.B(n_644),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_687),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_806),
.B(n_427),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_738),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_808),
.B(n_644),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_L g979 ( 
.A(n_780),
.B(n_300),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_754),
.B(n_586),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_808),
.B(n_644),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_740),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_754),
.B(n_586),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_809),
.B(n_302),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_809),
.B(n_644),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_698),
.B(n_644),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_832),
.A2(n_692),
.B(n_689),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_829),
.B(n_894),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_824),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_946),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_849),
.B(n_694),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_824),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_849),
.B(n_838),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_884),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_832),
.A2(n_692),
.B(n_689),
.Y(n_995)
);

NAND2x1_ASAP7_75t_L g996 ( 
.A(n_946),
.B(n_772),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_904),
.A2(n_692),
.B(n_689),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_884),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_836),
.A2(n_713),
.B(n_758),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_850),
.B(n_786),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_903),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_838),
.B(n_694),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_894),
.B(n_675),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_904),
.A2(n_692),
.B(n_714),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_884),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_848),
.B(n_876),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_884),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_836),
.B(n_713),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_883),
.A2(n_771),
.B(n_770),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_958),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_896),
.B(n_588),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_907),
.A2(n_714),
.B(n_725),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_848),
.B(n_696),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_876),
.B(n_696),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_907),
.A2(n_714),
.B(n_725),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_878),
.B(n_706),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_958),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_878),
.B(n_712),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_843),
.A2(n_680),
.B1(n_682),
.B2(n_671),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_831),
.B(n_675),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_861),
.A2(n_752),
.B(n_771),
.C(n_770),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_831),
.B(n_783),
.C(n_317),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_823),
.B(n_675),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_897),
.B(n_786),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_839),
.B(n_676),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_851),
.B(n_858),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_912),
.A2(n_787),
.B(n_725),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_912),
.A2(n_791),
.B(n_787),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_897),
.B(n_695),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_917),
.A2(n_879),
.B(n_877),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_917),
.A2(n_791),
.B(n_787),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_893),
.A2(n_780),
.B1(n_710),
.B2(n_705),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_842),
.A2(n_916),
.B(n_914),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_865),
.B(n_676),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_911),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_845),
.B(n_765),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_924),
.A2(n_791),
.B(n_708),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_875),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_933),
.A2(n_708),
.B(n_698),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_900),
.A2(n_776),
.B(n_775),
.C(n_745),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_852),
.A2(n_302),
.B1(n_330),
.B2(n_315),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_934),
.A2(n_882),
.B(n_906),
.Y(n_1042)
);

NOR2xp67_ASAP7_75t_L g1043 ( 
.A(n_825),
.B(n_717),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_867),
.A2(n_717),
.B(n_775),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_887),
.B(n_676),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_891),
.B(n_705),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_881),
.A2(n_708),
.B(n_698),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_846),
.A2(n_321),
.B(n_313),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_857),
.B(n_768),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_941),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_892),
.A2(n_854),
.B(n_847),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_874),
.A2(n_315),
.B1(n_330),
.B2(n_333),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_937),
.B(n_804),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_895),
.B(n_705),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_935),
.A2(n_776),
.B(n_745),
.C(n_748),
.Y(n_1055)
);

BUFx4f_ASAP7_75t_L g1056 ( 
.A(n_875),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_866),
.A2(n_748),
.B(n_740),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_881),
.A2(n_744),
.B(n_708),
.Y(n_1058)
);

AOI33xp33_ASAP7_75t_L g1059 ( 
.A1(n_826),
.A2(n_568),
.A3(n_566),
.B1(n_565),
.B2(n_563),
.B3(n_656),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_711),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_828),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_880),
.B(n_731),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_893),
.B(n_711),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_885),
.B(n_913),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_898),
.B(n_711),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_946),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_890),
.A2(n_963),
.B(n_863),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_961),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_830),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_926),
.B(n_719),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_965),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_890),
.A2(n_744),
.B(n_708),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_927),
.B(n_719),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_947),
.B(n_719),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_928),
.B(n_751),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_833),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_859),
.B(n_751),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_875),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_966),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_856),
.A2(n_957),
.B(n_837),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_935),
.A2(n_750),
.B(n_753),
.C(n_755),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_864),
.A2(n_753),
.B(n_750),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_894),
.B(n_751),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_894),
.B(n_766),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_835),
.A2(n_811),
.B(n_744),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_975),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_840),
.B(n_766),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_868),
.B(n_766),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_945),
.B(n_773),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_860),
.B(n_773),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_909),
.B(n_328),
.C(n_325),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_873),
.A2(n_811),
.B(n_744),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_902),
.A2(n_811),
.B(n_744),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_862),
.B(n_773),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_826),
.A2(n_368),
.B(n_341),
.C(n_356),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_964),
.B(n_794),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_946),
.B(n_794),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_889),
.B(n_356),
.C(n_333),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_949),
.B(n_794),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_949),
.B(n_755),
.Y(n_1100)
);

CKINVDCx10_ASAP7_75t_R g1101 ( 
.A(n_921),
.Y(n_1101)
);

AND2x6_ASAP7_75t_L g1102 ( 
.A(n_949),
.B(n_980),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_929),
.B(n_731),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_905),
.B(n_804),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_949),
.B(n_778),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_909),
.B(n_939),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_901),
.B(n_778),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_956),
.B(n_779),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_905),
.B(n_588),
.Y(n_1109)
);

OAI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_886),
.A2(n_358),
.B1(n_359),
.B2(n_440),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_931),
.A2(n_779),
.B(n_642),
.C(n_638),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_844),
.A2(n_742),
.B(n_683),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_956),
.B(n_780),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_834),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_905),
.B(n_596),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_888),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_869),
.A2(n_871),
.B(n_853),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_844),
.A2(n_742),
.B(n_683),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_951),
.B(n_780),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_951),
.A2(n_772),
.B1(n_359),
.B2(n_441),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_853),
.A2(n_742),
.B(n_683),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_936),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_870),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_918),
.B(n_329),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_962),
.B(n_789),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_959),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_962),
.B(n_938),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_871),
.A2(n_683),
.B(n_789),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_962),
.B(n_938),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_855),
.A2(n_358),
.B(n_365),
.C(n_368),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_940),
.A2(n_818),
.B(n_801),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_968),
.A2(n_609),
.B(n_618),
.C(n_615),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_855),
.A2(n_365),
.B(n_396),
.C(n_414),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_925),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_922),
.B(n_801),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_960),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_983),
.Y(n_1137)
);

BUFx4f_ASAP7_75t_L g1138 ( 
.A(n_960),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_979),
.A2(n_683),
.B(n_818),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_944),
.A2(n_973),
.B(n_972),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_972),
.A2(n_822),
.B(n_821),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_959),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_960),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_973),
.A2(n_822),
.B(n_821),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_918),
.B(n_338),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_915),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_976),
.A2(n_575),
.B(n_571),
.Y(n_1147)
);

AOI21x1_ASAP7_75t_L g1148 ( 
.A1(n_986),
.A2(n_578),
.B(n_575),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_922),
.B(n_396),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_923),
.B(n_414),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_894),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_976),
.A2(n_575),
.B(n_571),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_923),
.A2(n_345),
.B(n_339),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_970),
.A2(n_435),
.B(n_432),
.C(n_660),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_920),
.B(n_432),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_930),
.B(n_435),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_971),
.A2(n_575),
.B(n_571),
.Y(n_1157)
);

INVx6_ASAP7_75t_L g1158 ( 
.A(n_984),
.Y(n_1158)
);

NOR2x1_ASAP7_75t_L g1159 ( 
.A(n_950),
.B(n_596),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_908),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_974),
.A2(n_579),
.B(n_571),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_978),
.A2(n_581),
.B(n_579),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_894),
.B(n_644),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_827),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_984),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_952),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_981),
.A2(n_581),
.B(n_579),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1151),
.A2(n_950),
.B(n_970),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1006),
.B(n_899),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1001),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1068),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_993),
.B(n_967),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_1061),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1008),
.A2(n_955),
.B(n_969),
.C(n_943),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1049),
.B(n_919),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1148),
.A2(n_985),
.B(n_953),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1008),
.B(n_746),
.Y(n_1177)
);

AOI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1150),
.A2(n_872),
.B(n_955),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1106),
.B(n_977),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_991),
.B(n_982),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_999),
.A2(n_942),
.B1(n_932),
.B2(n_921),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1029),
.A2(n_948),
.B1(n_954),
.B2(n_986),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1024),
.B(n_347),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1071),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_SL g1185 ( 
.A(n_990),
.B(n_565),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_990),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1061),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1151),
.A2(n_581),
.B(n_579),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_990),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1036),
.B(n_603),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_1038),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_SL g1192 ( 
.A(n_1124),
.B(n_445),
.C(n_403),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1042),
.A2(n_581),
.B(n_583),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_SL g1194 ( 
.A(n_990),
.B(n_566),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1029),
.A2(n_353),
.B1(n_379),
.B2(n_382),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_1076),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1053),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1113),
.A2(n_583),
.B(n_578),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1019),
.A2(n_841),
.B(n_631),
.C(n_661),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_1069),
.B(n_984),
.Y(n_1200)
);

BUFx12f_ASAP7_75t_L g1201 ( 
.A(n_1122),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1079),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1126),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1026),
.B(n_1002),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1013),
.B(n_984),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1066),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1033),
.A2(n_583),
.B(n_578),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1086),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1050),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1124),
.B(n_984),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1160),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1137),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1145),
.A2(n_632),
.B(n_650),
.C(n_618),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1145),
.B(n_609),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1073),
.B(n_615),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1073),
.A2(n_624),
.B(n_628),
.C(n_650),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1030),
.A2(n_583),
.B(n_631),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1089),
.B(n_624),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1140),
.A2(n_633),
.B(n_628),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1035),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1064),
.B(n_294),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_1136),
.B(n_632),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_988),
.A2(n_634),
.B(n_633),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_988),
.A2(n_634),
.B(n_642),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1164),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1014),
.B(n_638),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1080),
.A2(n_654),
.B(n_617),
.Y(n_1227)
);

INVx3_ASAP7_75t_SL g1228 ( 
.A(n_1134),
.Y(n_1228)
);

AOI22x1_ASAP7_75t_SL g1229 ( 
.A1(n_1078),
.A2(n_423),
.B1(n_395),
.B2(n_348),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1051),
.B(n_617),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1024),
.A2(n_568),
.B(n_648),
.C(n_636),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1070),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1043),
.A2(n_430),
.B(n_362),
.C(n_411),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1022),
.B(n_375),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1052),
.A2(n_574),
.B(n_576),
.C(n_648),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1109),
.B(n_294),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1011),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1063),
.A2(n_626),
.B(n_617),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1116),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1011),
.B(n_286),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1067),
.A2(n_654),
.B(n_619),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1091),
.A2(n_438),
.B(n_376),
.C(n_424),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1056),
.B(n_286),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1000),
.B(n_413),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_SL g1245 ( 
.A1(n_1041),
.A2(n_576),
.B(n_574),
.C(n_413),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1153),
.B(n_383),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1016),
.B(n_619),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1115),
.B(n_386),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_SL g1249 ( 
.A(n_1165),
.B(n_400),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1103),
.A2(n_443),
.B1(n_442),
.B2(n_439),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1103),
.B(n_386),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1108),
.A2(n_636),
.B(n_626),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1104),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1166),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1062),
.B(n_994),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1143),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1166),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1098),
.A2(n_431),
.B(n_405),
.C(n_409),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1077),
.B(n_417),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1149),
.A2(n_418),
.B1(n_386),
.B2(n_413),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_994),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1098),
.A2(n_648),
.B(n_636),
.C(n_654),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1018),
.A2(n_654),
.B(n_636),
.C(n_626),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1125),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1077),
.B(n_1048),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1126),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1114),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1020),
.B(n_619),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1009),
.A2(n_626),
.B(n_619),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1074),
.B(n_644),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1065),
.A2(n_651),
.B(n_168),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1127),
.A2(n_651),
.B(n_386),
.C(n_12),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1126),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1027),
.A2(n_651),
.B(n_224),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_989),
.B(n_651),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1028),
.A2(n_651),
.B(n_214),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1123),
.Y(n_1277)
);

BUFx2_ASAP7_75t_SL g1278 ( 
.A(n_1102),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_992),
.B(n_1075),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1095),
.A2(n_8),
.B(n_9),
.C(n_12),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1056),
.B(n_651),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1075),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1138),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_SL g1284 ( 
.A(n_1165),
.B(n_651),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1138),
.B(n_651),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1095),
.A2(n_13),
.B(n_16),
.C(n_18),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1135),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1129),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_998),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1130),
.A2(n_23),
.B(n_24),
.C(n_26),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_998),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1146),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1060),
.B(n_24),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1130),
.A2(n_1133),
.B1(n_1154),
.B2(n_1158),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1031),
.A2(n_205),
.B(n_202),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1096),
.B(n_28),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1159),
.A2(n_200),
.B1(n_197),
.B2(n_189),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1101),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1059),
.B(n_28),
.Y(n_1299)
);

OAI22x1_ASAP7_75t_L g1300 ( 
.A1(n_1120),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1102),
.A2(n_173),
.B1(n_172),
.B2(n_162),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1102),
.B(n_29),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_997),
.A2(n_154),
.B(n_139),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1005),
.B(n_133),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1133),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1102),
.B(n_125),
.Y(n_1306)
);

INVx5_ASAP7_75t_L g1307 ( 
.A(n_1165),
.Y(n_1307)
);

AO32x2_ASAP7_75t_L g1308 ( 
.A1(n_1005),
.A2(n_36),
.A3(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1007),
.B(n_37),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_R g1310 ( 
.A(n_1102),
.B(n_117),
.Y(n_1310)
);

BUFx2_ASAP7_75t_SL g1311 ( 
.A(n_1007),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1165),
.B(n_106),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1032),
.A2(n_40),
.B(n_44),
.Y(n_1313)
);

AO21x1_ASAP7_75t_L g1314 ( 
.A1(n_1117),
.A2(n_1040),
.B(n_1021),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1119),
.A2(n_1021),
.B(n_1132),
.C(n_1055),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1110),
.A2(n_40),
.B(n_46),
.C(n_47),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1154),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1126),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1010),
.B(n_105),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1010),
.A2(n_1017),
.B1(n_1158),
.B2(n_1142),
.Y(n_1320)
);

NOR3xp33_ASAP7_75t_L g1321 ( 
.A(n_1110),
.B(n_1059),
.C(n_1132),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1142),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1087),
.B(n_94),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1142),
.B(n_53),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1228),
.Y(n_1325)
);

NAND2x1_ASAP7_75t_L g1326 ( 
.A(n_1206),
.B(n_1142),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1170),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1239),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1217),
.A2(n_1057),
.B(n_1092),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1176),
.A2(n_1141),
.B(n_1144),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1183),
.A2(n_1111),
.B(n_1023),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1168),
.A2(n_1204),
.B(n_1210),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1171),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1178),
.A2(n_1111),
.B(n_1040),
.C(n_1055),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1314),
.A2(n_1093),
.A3(n_1047),
.B(n_1058),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1197),
.B(n_1155),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1169),
.A2(n_1158),
.B1(n_1025),
.B2(n_1034),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1214),
.A2(n_1004),
.B(n_995),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1315),
.A2(n_1072),
.A3(n_1039),
.B(n_1085),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_L g1340 ( 
.A(n_1200),
.B(n_1097),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1226),
.B(n_1090),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1173),
.B(n_1156),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1184),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1187),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1236),
.B(n_1044),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1246),
.B(n_1152),
.C(n_1147),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1202),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1172),
.B(n_1094),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1247),
.A2(n_987),
.B(n_1012),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1208),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1172),
.B(n_1107),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1264),
.A2(n_1100),
.B1(n_1105),
.B2(n_1054),
.Y(n_1352)
);

OAI22x1_ASAP7_75t_L g1353 ( 
.A1(n_1181),
.A2(n_1003),
.B1(n_1084),
.B2(n_1083),
.Y(n_1353)
);

AO32x2_ASAP7_75t_L g1354 ( 
.A1(n_1287),
.A2(n_1044),
.A3(n_1081),
.B1(n_1082),
.B2(n_1131),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1271),
.A2(n_1081),
.B(n_1037),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1195),
.A2(n_1287),
.B1(n_1317),
.B2(n_1305),
.C(n_1178),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1209),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_1298),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1244),
.B(n_1099),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1207),
.A2(n_1167),
.B(n_1162),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1248),
.B(n_1088),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1234),
.B(n_1046),
.C(n_1045),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1307),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1255),
.B(n_1283),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1271),
.A2(n_1163),
.B(n_1015),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1174),
.A2(n_1161),
.B(n_1157),
.C(n_1128),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1218),
.B(n_1264),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1225),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1211),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1247),
.A2(n_1163),
.B(n_1003),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1196),
.Y(n_1371)
);

OAI22x1_ASAP7_75t_L g1372 ( 
.A1(n_1243),
.A2(n_1084),
.B1(n_1083),
.B2(n_56),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1230),
.A2(n_996),
.B(n_1139),
.Y(n_1373)
);

CKINVDCx6p67_ASAP7_75t_R g1374 ( 
.A(n_1201),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1255),
.B(n_1121),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1265),
.A2(n_1118),
.B(n_1112),
.C(n_56),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1190),
.B(n_53),
.Y(n_1377)
);

AO32x2_ASAP7_75t_L g1378 ( 
.A1(n_1317),
.A2(n_55),
.A3(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1302),
.A2(n_85),
.B(n_60),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1218),
.B(n_55),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1277),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1307),
.B(n_60),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1182),
.A2(n_61),
.B(n_62),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1193),
.A2(n_61),
.B(n_63),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1205),
.A2(n_66),
.B(n_67),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1321),
.A2(n_66),
.B1(n_70),
.B2(n_73),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1199),
.A2(n_1182),
.B(n_1219),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1198),
.A2(n_70),
.B(n_74),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1263),
.A2(n_1313),
.B(n_1238),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1179),
.B(n_78),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1191),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1179),
.B(n_81),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1203),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1192),
.A2(n_82),
.B(n_84),
.C(n_85),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1268),
.A2(n_1180),
.B(n_1270),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1215),
.A2(n_1293),
.B(n_1270),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1252),
.A2(n_1223),
.B(n_1224),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1180),
.A2(n_1269),
.B(n_1276),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1269),
.A2(n_1241),
.B(n_1245),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1274),
.A2(n_1303),
.B(n_1295),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1249),
.A2(n_1279),
.B(n_1284),
.Y(n_1401)
);

AO21x1_ASAP7_75t_L g1402 ( 
.A1(n_1294),
.A2(n_1305),
.B(n_1296),
.Y(n_1402)
);

CKINVDCx16_ASAP7_75t_R g1403 ( 
.A(n_1244),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1281),
.A2(n_1259),
.B(n_1233),
.C(n_1231),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1232),
.B(n_1282),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1294),
.A2(n_1216),
.A3(n_1272),
.B(n_1262),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1306),
.A2(n_1213),
.B(n_1307),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1306),
.A2(n_1307),
.B(n_1188),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1222),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1237),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1251),
.A2(n_1258),
.B(n_1175),
.C(n_1316),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1189),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1312),
.A2(n_1206),
.B(n_1275),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1288),
.A2(n_1300),
.A3(n_1309),
.B(n_1242),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1221),
.B(n_1253),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1235),
.A2(n_1320),
.B(n_1286),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1212),
.B(n_1256),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1318),
.A2(n_1289),
.B(n_1291),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1280),
.A2(n_1290),
.B(n_1220),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1177),
.B(n_1250),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1289),
.A2(n_1291),
.B(n_1186),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1203),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1222),
.B(n_1322),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1186),
.A2(n_1285),
.B(n_1292),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1195),
.A2(n_1257),
.A3(n_1254),
.B(n_1267),
.Y(n_1425)
);

CKINVDCx9p33_ASAP7_75t_R g1426 ( 
.A(n_1229),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1203),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1222),
.B(n_1240),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1299),
.A2(n_1297),
.B(n_1323),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1301),
.A2(n_1319),
.B(n_1324),
.C(n_1278),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1319),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1266),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1260),
.A2(n_1304),
.B1(n_1323),
.B2(n_1194),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1266),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1185),
.A2(n_1323),
.B(n_1310),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1323),
.A2(n_1304),
.B(n_1189),
.Y(n_1436)
);

OAI211xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1308),
.A2(n_1304),
.B(n_1311),
.C(n_1273),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1266),
.A2(n_1273),
.B(n_1261),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1273),
.A2(n_1261),
.B(n_1308),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1308),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_SL g1441 ( 
.A1(n_1306),
.A2(n_1302),
.B(n_1129),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_SL g1442 ( 
.A1(n_1169),
.A2(n_1006),
.B(n_993),
.C(n_1178),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1168),
.A2(n_1151),
.B(n_673),
.Y(n_1443)
);

AOI221x1_ASAP7_75t_L g1444 ( 
.A1(n_1178),
.A2(n_1006),
.B1(n_1008),
.B2(n_993),
.C(n_1271),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1228),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1168),
.A2(n_1151),
.B(n_673),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1204),
.A2(n_1006),
.B1(n_993),
.B2(n_1008),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1315),
.A2(n_1006),
.B(n_1042),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1314),
.A2(n_1315),
.A3(n_1182),
.B(n_1294),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1168),
.A2(n_1006),
.B(n_673),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1315),
.A2(n_1006),
.B(n_1042),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1178),
.A2(n_1006),
.B(n_1008),
.C(n_993),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1168),
.A2(n_1151),
.B(n_673),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1315),
.A2(n_1006),
.B(n_1042),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1168),
.A2(n_1151),
.B(n_673),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1168),
.A2(n_1151),
.B(n_673),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1230),
.A2(n_1140),
.B(n_1182),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1183),
.B(n_1008),
.C(n_836),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1170),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1170),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1244),
.B(n_1008),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1183),
.A2(n_1008),
.B1(n_836),
.B2(n_999),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1204),
.B(n_1006),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1170),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1168),
.A2(n_1151),
.B(n_673),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1314),
.A2(n_1315),
.A3(n_1182),
.B(n_1294),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1244),
.B(n_1008),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_SL g1474 ( 
.A(n_1183),
.B(n_1008),
.C(n_1006),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1190),
.B(n_1036),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1187),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1183),
.B(n_1008),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1204),
.B(n_1006),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1187),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1204),
.B(n_1006),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1239),
.Y(n_1483)
);

AND2x4_ASAP7_75t_SL g1484 ( 
.A(n_1225),
.B(n_1061),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1255),
.B(n_1283),
.Y(n_1485)
);

INVx5_ASAP7_75t_L g1486 ( 
.A(n_1304),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1236),
.B(n_846),
.Y(n_1487)
);

INVxp67_ASAP7_75t_SL g1488 ( 
.A(n_1187),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_SL g1489 ( 
.A1(n_1169),
.A2(n_1006),
.B(n_993),
.C(n_1178),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1228),
.Y(n_1490)
);

AOI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1230),
.A2(n_1140),
.B(n_1182),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1227),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1357),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1368),
.Y(n_1495)
);

BUFx10_ASAP7_75t_L g1496 ( 
.A(n_1484),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1328),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1477),
.A2(n_1462),
.B(n_1467),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1422),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1327),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1333),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1468),
.A2(n_1478),
.B1(n_1482),
.B2(n_1466),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1483),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1343),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1474),
.A2(n_1356),
.B1(n_1472),
.B2(n_1447),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1363),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1356),
.A2(n_1472),
.B1(n_1447),
.B2(n_1402),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1490),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1347),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1403),
.A2(n_1386),
.B1(n_1420),
.B2(n_1486),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1386),
.A2(n_1482),
.B1(n_1478),
.B2(n_1468),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1350),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1374),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1452),
.A2(n_1444),
.B(n_1362),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1412),
.Y(n_1515)
);

INVx6_ASAP7_75t_L g1516 ( 
.A(n_1412),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1422),
.Y(n_1517)
);

BUFx8_ASAP7_75t_L g1518 ( 
.A(n_1445),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1363),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1358),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1464),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1423),
.Y(n_1522)
);

CKINVDCx11_ASAP7_75t_R g1523 ( 
.A(n_1358),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1439),
.Y(n_1524)
);

BUFx8_ASAP7_75t_L g1525 ( 
.A(n_1409),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1364),
.A2(n_1485),
.B1(n_1325),
.B2(n_1423),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1465),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1475),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1469),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1486),
.A2(n_1367),
.B1(n_1433),
.B2(n_1405),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1448),
.A2(n_1455),
.B1(n_1451),
.B2(n_1429),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1486),
.A2(n_1440),
.B1(n_1455),
.B2(n_1448),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1426),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1451),
.A2(n_1429),
.B1(n_1380),
.B2(n_1437),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1486),
.A2(n_1440),
.B1(n_1380),
.B2(n_1378),
.Y(n_1535)
);

INVx6_ASAP7_75t_L g1536 ( 
.A(n_1364),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1367),
.B(n_1487),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1485),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1391),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_L g1540 ( 
.A(n_1427),
.Y(n_1540)
);

CKINVDCx11_ASAP7_75t_R g1541 ( 
.A(n_1325),
.Y(n_1541)
);

BUFx12f_ASAP7_75t_L g1542 ( 
.A(n_1377),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1369),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1476),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1394),
.A2(n_1411),
.B(n_1428),
.Y(n_1545)
);

CKINVDCx6p67_ASAP7_75t_R g1546 ( 
.A(n_1427),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1371),
.Y(n_1547)
);

INVx6_ASAP7_75t_L g1548 ( 
.A(n_1427),
.Y(n_1548)
);

INVx6_ASAP7_75t_L g1549 ( 
.A(n_1415),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1410),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1410),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1418),
.B(n_1421),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1419),
.A2(n_1361),
.B1(n_1390),
.B2(n_1392),
.Y(n_1553)
);

CKINVDCx6p67_ASAP7_75t_R g1554 ( 
.A(n_1405),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1381),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1336),
.A2(n_1431),
.B1(n_1342),
.B2(n_1372),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1488),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1390),
.A2(n_1392),
.B1(n_1341),
.B2(n_1351),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1344),
.Y(n_1559)
);

BUFx8_ASAP7_75t_SL g1560 ( 
.A(n_1434),
.Y(n_1560)
);

INVx6_ASAP7_75t_L g1561 ( 
.A(n_1375),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1419),
.A2(n_1385),
.B1(n_1387),
.B2(n_1416),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1378),
.A2(n_1382),
.B1(n_1387),
.B2(n_1416),
.Y(n_1563)
);

BUFx8_ASAP7_75t_SL g1564 ( 
.A(n_1393),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1341),
.A2(n_1345),
.B1(n_1351),
.B2(n_1355),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1481),
.B(n_1425),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1442),
.A2(n_1489),
.B(n_1331),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1355),
.A2(n_1348),
.B1(n_1441),
.B2(n_1359),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1348),
.A2(n_1382),
.B1(n_1389),
.B2(n_1450),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1389),
.A2(n_1450),
.B1(n_1332),
.B2(n_1352),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1393),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1352),
.A2(n_1353),
.B1(n_1337),
.B2(n_1398),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1425),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1430),
.A2(n_1417),
.B1(n_1331),
.B2(n_1407),
.Y(n_1574)
);

CKINVDCx11_ASAP7_75t_R g1575 ( 
.A(n_1375),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1436),
.A2(n_1376),
.B(n_1383),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1414),
.B(n_1471),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1432),
.Y(n_1578)
);

BUFx10_ASAP7_75t_L g1579 ( 
.A(n_1379),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1432),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1334),
.A2(n_1436),
.B1(n_1337),
.B2(n_1413),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1425),
.B(n_1414),
.Y(n_1582)
);

BUFx8_ASAP7_75t_SL g1583 ( 
.A(n_1401),
.Y(n_1583)
);

CKINVDCx14_ASAP7_75t_R g1584 ( 
.A(n_1340),
.Y(n_1584)
);

CKINVDCx6p67_ASAP7_75t_R g1585 ( 
.A(n_1378),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1414),
.B(n_1471),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1438),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1435),
.A2(n_1346),
.B1(n_1365),
.B2(n_1400),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1449),
.B(n_1471),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1384),
.Y(n_1590)
);

BUFx12f_ASAP7_75t_L g1591 ( 
.A(n_1326),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1424),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1408),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1395),
.A2(n_1365),
.B1(n_1399),
.B2(n_1388),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1449),
.Y(n_1595)
);

CKINVDCx14_ASAP7_75t_R g1596 ( 
.A(n_1404),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1399),
.A2(n_1397),
.B1(n_1370),
.B2(n_1338),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1397),
.A2(n_1453),
.B1(n_1470),
.B2(n_1460),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1406),
.Y(n_1599)
);

BUFx12f_ASAP7_75t_L g1600 ( 
.A(n_1396),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1406),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1406),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1449),
.A2(n_1443),
.B1(n_1459),
.B2(n_1446),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1461),
.A2(n_1491),
.B(n_1366),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1373),
.A2(n_1349),
.B1(n_1493),
.B2(n_1457),
.Y(n_1605)
);

BUFx10_ASAP7_75t_L g1606 ( 
.A(n_1339),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1335),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1335),
.Y(n_1608)
);

BUFx12f_ASAP7_75t_L g1609 ( 
.A(n_1335),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1454),
.A2(n_1458),
.B1(n_1480),
.B2(n_1479),
.Y(n_1610)
);

CKINVDCx11_ASAP7_75t_R g1611 ( 
.A(n_1354),
.Y(n_1611)
);

BUFx10_ASAP7_75t_L g1612 ( 
.A(n_1354),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1456),
.A2(n_1492),
.B1(n_1473),
.B2(n_1463),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1354),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1360),
.Y(n_1615)
);

BUFx12f_ASAP7_75t_L g1616 ( 
.A(n_1329),
.Y(n_1616)
);

BUFx12f_ASAP7_75t_L g1617 ( 
.A(n_1330),
.Y(n_1617)
);

OAI22x1_ASAP7_75t_L g1618 ( 
.A1(n_1467),
.A2(n_1462),
.B1(n_1477),
.B2(n_1466),
.Y(n_1618)
);

INVx6_ASAP7_75t_L g1619 ( 
.A(n_1328),
.Y(n_1619)
);

CKINVDCx6p67_ASAP7_75t_R g1620 ( 
.A(n_1374),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1621)
);

BUFx2_ASAP7_75t_SL g1622 ( 
.A(n_1328),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1462),
.A2(n_1008),
.B1(n_1477),
.B2(n_1467),
.Y(n_1623)
);

CKINVDCx11_ASAP7_75t_R g1624 ( 
.A(n_1358),
.Y(n_1624)
);

NAND2x1p5_ASAP7_75t_L g1625 ( 
.A(n_1486),
.B(n_990),
.Y(n_1625)
);

CKINVDCx11_ASAP7_75t_R g1626 ( 
.A(n_1358),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1357),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1484),
.Y(n_1629)
);

CKINVDCx11_ASAP7_75t_R g1630 ( 
.A(n_1358),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1477),
.A2(n_1008),
.B1(n_1462),
.B2(n_1474),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1472),
.A2(n_1008),
.B1(n_1477),
.B2(n_1462),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1472),
.A2(n_1008),
.B1(n_1477),
.B2(n_1462),
.Y(n_1635)
);

CKINVDCx10_ASAP7_75t_R g1636 ( 
.A(n_1403),
.Y(n_1636)
);

BUFx8_ASAP7_75t_L g1637 ( 
.A(n_1445),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1447),
.B(n_1477),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1472),
.A2(n_1462),
.B1(n_1467),
.B2(n_1403),
.Y(n_1640)
);

CKINVDCx11_ASAP7_75t_R g1641 ( 
.A(n_1358),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1472),
.A2(n_1008),
.B1(n_1477),
.B2(n_1462),
.Y(n_1643)
);

BUFx12f_ASAP7_75t_L g1644 ( 
.A(n_1490),
.Y(n_1644)
);

INVx6_ASAP7_75t_L g1645 ( 
.A(n_1328),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1328),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1447),
.B(n_1477),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1447),
.B(n_1477),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1357),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1368),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1462),
.A2(n_1008),
.B1(n_1477),
.B2(n_1467),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1008),
.B2(n_1474),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1484),
.Y(n_1654)
);

BUFx8_ASAP7_75t_L g1655 ( 
.A(n_1445),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1357),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1462),
.A2(n_1008),
.B1(n_1477),
.B2(n_1467),
.Y(n_1657)
);

INVx6_ASAP7_75t_L g1658 ( 
.A(n_1328),
.Y(n_1658)
);

INVx4_ASAP7_75t_L g1659 ( 
.A(n_1490),
.Y(n_1659)
);

BUFx8_ASAP7_75t_L g1660 ( 
.A(n_1445),
.Y(n_1660)
);

OAI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1472),
.A2(n_1462),
.B1(n_1467),
.B2(n_1403),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1368),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1368),
.Y(n_1663)
);

BUFx8_ASAP7_75t_SL g1664 ( 
.A(n_1490),
.Y(n_1664)
);

OAI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1472),
.A2(n_1462),
.B1(n_1467),
.B2(n_1403),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1609),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1573),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1549),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1595),
.Y(n_1669)
);

OA21x2_ASAP7_75t_L g1670 ( 
.A1(n_1604),
.A2(n_1514),
.B(n_1594),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1608),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1594),
.A2(n_1597),
.B(n_1570),
.Y(n_1672)
);

INVx5_ASAP7_75t_SL g1673 ( 
.A(n_1554),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1577),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1601),
.B(n_1602),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1502),
.B(n_1639),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1549),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1582),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1600),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1593),
.A2(n_1625),
.B(n_1574),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1589),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1586),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1557),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1610),
.A2(n_1613),
.B(n_1605),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1610),
.A2(n_1613),
.B(n_1605),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1524),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1566),
.B(n_1585),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1597),
.A2(n_1570),
.B(n_1576),
.Y(n_1688)
);

OAI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1647),
.A2(n_1648),
.B1(n_1498),
.B2(n_1652),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1607),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1607),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1563),
.B(n_1507),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1606),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1495),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1575),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1563),
.B(n_1507),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1599),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1617),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1590),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1592),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1598),
.A2(n_1552),
.B(n_1588),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1500),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1552),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1598),
.A2(n_1581),
.B(n_1567),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1543),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1625),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1537),
.B(n_1623),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1501),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1549),
.Y(n_1709)
);

AO21x1_ASAP7_75t_SL g1710 ( 
.A1(n_1534),
.A2(n_1531),
.B(n_1562),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1612),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1558),
.A2(n_1530),
.B(n_1545),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1504),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1547),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1509),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1562),
.A2(n_1572),
.B(n_1531),
.Y(n_1716)
);

CKINVDCx16_ASAP7_75t_R g1717 ( 
.A(n_1571),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1572),
.A2(n_1569),
.B(n_1568),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1512),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1621),
.B(n_1628),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1612),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1521),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1534),
.A2(n_1569),
.B(n_1568),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1527),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1529),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1616),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1565),
.B(n_1532),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1565),
.B(n_1532),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1587),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1535),
.B(n_1505),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1555),
.Y(n_1731)
);

OA21x2_ASAP7_75t_L g1732 ( 
.A1(n_1614),
.A2(n_1553),
.B(n_1505),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1615),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1561),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1561),
.B(n_1618),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1561),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1526),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1535),
.B(n_1553),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1494),
.Y(n_1739)
);

AOI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1640),
.A2(n_1665),
.B(n_1661),
.C(n_1530),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1640),
.B(n_1661),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1579),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1665),
.B(n_1559),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1621),
.B(n_1628),
.Y(n_1744)
);

AO21x2_ASAP7_75t_L g1745 ( 
.A1(n_1558),
.A2(n_1556),
.B(n_1603),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1627),
.Y(n_1746)
);

AOI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1578),
.A2(n_1656),
.B(n_1649),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1596),
.A2(n_1584),
.B1(n_1634),
.B2(n_1643),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1579),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1506),
.A2(n_1519),
.B(n_1511),
.Y(n_1750)
);

BUFx2_ASAP7_75t_SL g1751 ( 
.A(n_1551),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1634),
.B(n_1635),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1611),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1603),
.Y(n_1754)
);

OAI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1511),
.A2(n_1632),
.B(n_1653),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1583),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1632),
.A2(n_1633),
.B(n_1653),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1496),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1499),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1635),
.B(n_1643),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1499),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1550),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1544),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1517),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1528),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1510),
.B(n_1650),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1525),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1633),
.B(n_1638),
.Y(n_1768)
);

AO21x2_ASAP7_75t_L g1769 ( 
.A1(n_1510),
.A2(n_1650),
.B(n_1638),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1642),
.A2(n_1631),
.B(n_1591),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1580),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1642),
.A2(n_1546),
.B(n_1516),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1522),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1536),
.Y(n_1774)
);

AND2x6_ASAP7_75t_L g1775 ( 
.A(n_1654),
.B(n_1497),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1536),
.A2(n_1538),
.B(n_1548),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1538),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1538),
.B(n_1528),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1525),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1515),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1515),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1629),
.B(n_1542),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1516),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1540),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1663),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1540),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1548),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1564),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1651),
.B(n_1662),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1496),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1560),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1541),
.B(n_1622),
.Y(n_1792)
);

OA21x2_ASAP7_75t_L g1793 ( 
.A1(n_1539),
.A2(n_1637),
.B(n_1660),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1659),
.B(n_1503),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1619),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1619),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1518),
.A2(n_1655),
.B(n_1660),
.Y(n_1798)
);

AO21x1_ASAP7_75t_L g1799 ( 
.A1(n_1518),
.A2(n_1655),
.B(n_1636),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1619),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1646),
.B(n_1513),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1680),
.A2(n_1508),
.B(n_1533),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1717),
.B(n_1664),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1717),
.B(n_1644),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1689),
.B(n_1658),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1748),
.A2(n_1645),
.B1(n_1658),
.B2(n_1620),
.Y(n_1806)
);

AO21x2_ASAP7_75t_L g1807 ( 
.A1(n_1684),
.A2(n_1685),
.B(n_1701),
.Y(n_1807)
);

O2A1O1Ixp33_ASAP7_75t_SL g1808 ( 
.A1(n_1740),
.A2(n_1520),
.B(n_1523),
.C(n_1624),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1741),
.A2(n_1645),
.B1(n_1658),
.B2(n_1641),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1705),
.B(n_1645),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1702),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1676),
.B(n_1626),
.Y(n_1812)
);

NOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1680),
.B(n_1630),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1757),
.A2(n_1755),
.B(n_1704),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1733),
.B(n_1683),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1757),
.A2(n_1755),
.B(n_1704),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1733),
.B(n_1678),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_SL g1818 ( 
.A1(n_1752),
.A2(n_1760),
.B(n_1743),
.Y(n_1818)
);

AO32x2_ASAP7_75t_L g1819 ( 
.A1(n_1737),
.A2(n_1706),
.A3(n_1681),
.B1(n_1682),
.B2(n_1678),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1702),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1775),
.Y(n_1821)
);

OR2x2_ASAP7_75t_SL g1822 ( 
.A(n_1798),
.B(n_1793),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1760),
.A2(n_1766),
.B(n_1718),
.C(n_1770),
.Y(n_1823)
);

BUFx12f_ASAP7_75t_L g1824 ( 
.A(n_1767),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1687),
.B(n_1753),
.Y(n_1825)
);

O2A1O1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1720),
.A2(n_1744),
.B(n_1768),
.C(n_1766),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1682),
.B(n_1681),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1753),
.B(n_1709),
.Y(n_1828)
);

NAND4xp25_ASAP7_75t_L g1829 ( 
.A(n_1707),
.B(n_1692),
.C(n_1696),
.D(n_1738),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1668),
.B(n_1677),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1756),
.A2(n_1730),
.B1(n_1692),
.B2(n_1696),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1737),
.B(n_1727),
.Y(n_1832)
);

AND2x2_ASAP7_75t_SL g1833 ( 
.A(n_1730),
.B(n_1738),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1735),
.B(n_1718),
.Y(n_1834)
);

A2O1A1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1770),
.A2(n_1727),
.B(n_1728),
.C(n_1754),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1728),
.A2(n_1754),
.B(n_1756),
.C(n_1772),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1789),
.B(n_1694),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1666),
.B(n_1773),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1666),
.B(n_1735),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1735),
.B(n_1772),
.Y(n_1840)
);

O2A1O1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1769),
.A2(n_1756),
.B(n_1712),
.C(n_1745),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1735),
.B(n_1715),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1735),
.B(n_1715),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1763),
.B(n_1722),
.Y(n_1844)
);

NAND2xp33_ASAP7_75t_L g1845 ( 
.A(n_1775),
.B(n_1756),
.Y(n_1845)
);

NAND4xp25_ASAP7_75t_L g1846 ( 
.A(n_1695),
.B(n_1679),
.C(n_1765),
.D(n_1792),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1769),
.A2(n_1712),
.B1(n_1716),
.B2(n_1688),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1675),
.B(n_1776),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1679),
.A2(n_1673),
.B1(n_1695),
.B2(n_1779),
.Y(n_1849)
);

AO32x1_ASAP7_75t_L g1850 ( 
.A1(n_1669),
.A2(n_1671),
.A3(n_1690),
.B1(n_1674),
.B2(n_1691),
.Y(n_1850)
);

AO32x2_ASAP7_75t_L g1851 ( 
.A1(n_1706),
.A2(n_1758),
.A3(n_1790),
.B1(n_1732),
.B2(n_1710),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1708),
.Y(n_1852)
);

NAND4xp25_ASAP7_75t_L g1853 ( 
.A(n_1695),
.B(n_1765),
.C(n_1792),
.D(n_1779),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1701),
.A2(n_1742),
.B(n_1749),
.C(n_1758),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1722),
.B(n_1725),
.Y(n_1855)
);

A2O1A1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1742),
.A2(n_1749),
.B(n_1790),
.C(n_1710),
.Y(n_1856)
);

OA21x2_ASAP7_75t_L g1857 ( 
.A1(n_1684),
.A2(n_1685),
.B(n_1750),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1712),
.B(n_1698),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1725),
.B(n_1708),
.Y(n_1859)
);

AO21x2_ASAP7_75t_L g1860 ( 
.A1(n_1747),
.A2(n_1699),
.B(n_1693),
.Y(n_1860)
);

A2O1A1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1742),
.A2(n_1749),
.B(n_1750),
.C(n_1698),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_SL g1862 ( 
.A(n_1765),
.B(n_1767),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1747),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1785),
.B(n_1782),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1751),
.B(n_1714),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1686),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1713),
.Y(n_1867)
);

O2A1O1Ixp33_ASAP7_75t_SL g1868 ( 
.A1(n_1794),
.A2(n_1791),
.B(n_1788),
.C(n_1778),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1713),
.B(n_1719),
.Y(n_1869)
);

OR2x6_ASAP7_75t_L g1870 ( 
.A(n_1726),
.B(n_1688),
.Y(n_1870)
);

AND2x6_ASAP7_75t_L g1871 ( 
.A(n_1673),
.B(n_1726),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1800),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1719),
.Y(n_1873)
);

A2O1A1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1742),
.A2(n_1749),
.B(n_1698),
.C(n_1796),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1762),
.B(n_1801),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1726),
.B(n_1688),
.Y(n_1876)
);

OR2x6_ASAP7_75t_L g1877 ( 
.A(n_1726),
.B(n_1688),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1697),
.A2(n_1699),
.B(n_1669),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1675),
.B(n_1776),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1775),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1716),
.A2(n_1723),
.B(n_1672),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1769),
.A2(n_1745),
.B(n_1797),
.C(n_1796),
.Y(n_1882)
);

OA21x2_ASAP7_75t_L g1883 ( 
.A1(n_1697),
.A2(n_1667),
.B(n_1700),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1675),
.B(n_1776),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1759),
.B(n_1761),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_SL g1886 ( 
.A(n_1745),
.B(n_1726),
.Y(n_1886)
);

AO21x1_ASAP7_75t_L g1887 ( 
.A1(n_1739),
.A2(n_1746),
.B(n_1724),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1673),
.A2(n_1716),
.B1(n_1797),
.B2(n_1791),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1761),
.B(n_1764),
.Y(n_1889)
);

OR2x6_ASAP7_75t_L g1890 ( 
.A(n_1726),
.B(n_1675),
.Y(n_1890)
);

NOR3xp33_ASAP7_75t_SL g1891 ( 
.A(n_1780),
.B(n_1781),
.C(n_1783),
.Y(n_1891)
);

AO32x2_ASAP7_75t_L g1892 ( 
.A1(n_1706),
.A2(n_1732),
.A3(n_1674),
.B1(n_1716),
.B2(n_1670),
.Y(n_1892)
);

O2A1O1Ixp33_ASAP7_75t_SL g1893 ( 
.A1(n_1788),
.A2(n_1783),
.B(n_1780),
.C(n_1781),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1788),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1799),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1801),
.Y(n_1896)
);

A2O1A1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1698),
.A2(n_1734),
.B(n_1777),
.C(n_1774),
.Y(n_1897)
);

INVxp67_ASAP7_75t_SL g1898 ( 
.A(n_1863),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1881),
.B(n_1672),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1871),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1887),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1878),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1817),
.B(n_1815),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1878),
.Y(n_1904)
);

CKINVDCx16_ASAP7_75t_R g1905 ( 
.A(n_1862),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1811),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1855),
.B(n_1732),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1819),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1822),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1820),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1866),
.B(n_1732),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1883),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1852),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1848),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1819),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1883),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1867),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1881),
.B(n_1672),
.Y(n_1918)
);

AND2x2_ASAP7_75t_SL g1919 ( 
.A(n_1833),
.B(n_1672),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1892),
.B(n_1711),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1892),
.B(n_1711),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1873),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1844),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1814),
.B(n_1721),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1819),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1806),
.A2(n_1723),
.B1(n_1775),
.B2(n_1736),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1816),
.B(n_1670),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1816),
.B(n_1670),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1857),
.B(n_1670),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1827),
.B(n_1729),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1834),
.B(n_1671),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1869),
.Y(n_1932)
);

AND2x4_ASAP7_75t_SL g1933 ( 
.A(n_1821),
.B(n_1880),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1859),
.Y(n_1934)
);

INVx4_ASAP7_75t_L g1935 ( 
.A(n_1871),
.Y(n_1935)
);

BUFx5_ASAP7_75t_L g1936 ( 
.A(n_1871),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1860),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1851),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1871),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1870),
.B(n_1876),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1812),
.B(n_1795),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1860),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1848),
.B(n_1703),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1823),
.B(n_1731),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_SL g1945 ( 
.A1(n_1895),
.A2(n_1723),
.B1(n_1673),
.B2(n_1798),
.Y(n_1945)
);

NOR2x1_ASAP7_75t_SL g1946 ( 
.A(n_1877),
.B(n_1703),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1850),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1850),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1890),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1850),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1912),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1902),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1939),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1912),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1940),
.B(n_1879),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1902),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1940),
.B(n_1879),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1940),
.B(n_1884),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1904),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1923),
.Y(n_1960)
);

OAI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1945),
.A2(n_1818),
.B1(n_1826),
.B2(n_1841),
.C(n_1835),
.Y(n_1961)
);

BUFx3_ASAP7_75t_L g1962 ( 
.A(n_1939),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1912),
.Y(n_1963)
);

OAI33xp33_ASAP7_75t_L g1964 ( 
.A1(n_1901),
.A2(n_1831),
.A3(n_1829),
.B1(n_1853),
.B2(n_1846),
.B3(n_1849),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1904),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1906),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1916),
.Y(n_1967)
);

AO21x2_ASAP7_75t_L g1968 ( 
.A1(n_1937),
.A2(n_1854),
.B(n_1861),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1914),
.B(n_1840),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1909),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1914),
.B(n_1840),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1898),
.B(n_1847),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1898),
.B(n_1882),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1909),
.B(n_1840),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1907),
.B(n_1807),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1919),
.A2(n_1813),
.B1(n_1829),
.B2(n_1723),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_1916),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1910),
.Y(n_1978)
);

AOI331xp33_ASAP7_75t_L g1979 ( 
.A1(n_1901),
.A2(n_1818),
.A3(n_1802),
.B1(n_1875),
.B2(n_1804),
.B3(n_1803),
.C1(n_1799),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1907),
.B(n_1842),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1909),
.B(n_1851),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_SL g1982 ( 
.A1(n_1905),
.A2(n_1809),
.B1(n_1798),
.B2(n_1793),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1934),
.B(n_1858),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1943),
.B(n_1851),
.Y(n_1984)
);

AO21x2_ASAP7_75t_L g1985 ( 
.A1(n_1937),
.A2(n_1886),
.B(n_1888),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1913),
.Y(n_1986)
);

NOR4xp25_ASAP7_75t_SL g1987 ( 
.A(n_1908),
.B(n_1893),
.C(n_1868),
.D(n_1874),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1943),
.B(n_1839),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1903),
.B(n_1843),
.Y(n_1989)
);

AOI31xp33_ASAP7_75t_L g1990 ( 
.A1(n_1945),
.A2(n_1813),
.A3(n_1808),
.B(n_1809),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1917),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1903),
.B(n_1885),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1944),
.A2(n_1805),
.B1(n_1836),
.B2(n_1828),
.C(n_1832),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1934),
.B(n_1858),
.Y(n_1994)
);

OAI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1926),
.A2(n_1853),
.B1(n_1846),
.B2(n_1862),
.C(n_1856),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1919),
.A2(n_1897),
.B(n_1891),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1911),
.B(n_1889),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1933),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1911),
.B(n_1729),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1943),
.B(n_1838),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1917),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1920),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1922),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1922),
.Y(n_2004)
);

INVx5_ASAP7_75t_SL g2005 ( 
.A(n_1919),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1966),
.B(n_1932),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1952),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1966),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1974),
.B(n_1946),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_2005),
.B(n_1946),
.Y(n_2010)
);

AND2x4_ASAP7_75t_SL g2011 ( 
.A(n_1960),
.B(n_1900),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_2005),
.B(n_1970),
.Y(n_2012)
);

INVxp67_ASAP7_75t_L g2013 ( 
.A(n_1973),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1978),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1951),
.Y(n_2015)
);

BUFx12f_ASAP7_75t_L g2016 ( 
.A(n_1953),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1999),
.B(n_1975),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1951),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_2005),
.B(n_1938),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1951),
.Y(n_2020)
);

BUFx12f_ASAP7_75t_L g2021 ( 
.A(n_1953),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1978),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1951),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_2002),
.B(n_1938),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_1970),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2005),
.B(n_1974),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1986),
.B(n_1908),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1963),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2005),
.B(n_1938),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1986),
.B(n_1915),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1981),
.B(n_1938),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1979),
.B(n_1905),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1991),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1991),
.Y(n_2034)
);

NOR4xp25_ASAP7_75t_SL g2035 ( 
.A(n_1961),
.B(n_1915),
.C(n_1925),
.D(n_1894),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2001),
.B(n_1925),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1963),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2001),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1999),
.B(n_1944),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1975),
.B(n_1930),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2002),
.B(n_1938),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2002),
.B(n_1938),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2003),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1981),
.B(n_1938),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2003),
.B(n_1920),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1955),
.B(n_1949),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2004),
.B(n_1921),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2004),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_1961),
.B(n_1993),
.C(n_1973),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1952),
.B(n_1921),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1963),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1955),
.B(n_1949),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1956),
.Y(n_2053)
);

AND2x4_ASAP7_75t_L g2054 ( 
.A(n_1998),
.B(n_1931),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1998),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1954),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1957),
.B(n_1924),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1953),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1956),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1959),
.B(n_1921),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1959),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2007),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_2026),
.B(n_1962),
.Y(n_2063)
);

BUFx3_ASAP7_75t_L g2064 ( 
.A(n_2016),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2039),
.B(n_1980),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2013),
.B(n_1993),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2008),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2028),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2026),
.B(n_1957),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2008),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2049),
.A2(n_1982),
.B1(n_1964),
.B2(n_1995),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2039),
.B(n_1980),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2014),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2014),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_SL g2075 ( 
.A1(n_2049),
.A2(n_1982),
.B1(n_1996),
.B2(n_1995),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2046),
.B(n_1958),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_2012),
.B(n_1962),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2040),
.B(n_1989),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2046),
.B(n_1958),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2052),
.B(n_1988),
.Y(n_2080)
);

NOR5xp2_ASAP7_75t_L g2081 ( 
.A(n_2013),
.B(n_1990),
.C(n_1996),
.D(n_1967),
.E(n_1979),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2022),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_2012),
.B(n_2009),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2009),
.B(n_1962),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2032),
.A2(n_1990),
.B1(n_1976),
.B2(n_1987),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2025),
.B(n_1972),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2040),
.B(n_1989),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_2016),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_SL g2089 ( 
.A(n_2016),
.B(n_1964),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_L g2090 ( 
.A(n_2025),
.B(n_1788),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2052),
.B(n_1988),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2022),
.Y(n_2092)
);

NAND3xp33_ASAP7_75t_L g2093 ( 
.A(n_2035),
.B(n_1987),
.C(n_1972),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_2021),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2057),
.B(n_2058),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_2021),
.Y(n_2096)
);

INVx1_ASAP7_75t_SL g2097 ( 
.A(n_2021),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2017),
.B(n_1992),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2033),
.Y(n_2099)
);

INVxp67_ASAP7_75t_L g2100 ( 
.A(n_2055),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2017),
.B(n_1992),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2033),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2034),
.Y(n_2103)
);

OAI33xp33_ASAP7_75t_L g2104 ( 
.A1(n_2027),
.A2(n_1965),
.A3(n_1983),
.B1(n_1994),
.B2(n_1950),
.B3(n_1948),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2057),
.B(n_2011),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_2010),
.B(n_1998),
.Y(n_2106)
);

AOI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2035),
.A2(n_1968),
.B(n_1845),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2011),
.B(n_1997),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_2011),
.B(n_1824),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2034),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2038),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2038),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_2055),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2028),
.Y(n_2114)
);

OAI31xp33_ASAP7_75t_L g2115 ( 
.A1(n_2019),
.A2(n_1927),
.A3(n_1928),
.B(n_1971),
.Y(n_2115)
);

NAND2x1p5_ASAP7_75t_L g2116 ( 
.A(n_2010),
.B(n_1900),
.Y(n_2116)
);

NOR3xp33_ASAP7_75t_L g2117 ( 
.A(n_2019),
.B(n_1928),
.C(n_1927),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_2009),
.Y(n_2118)
);

INVxp67_ASAP7_75t_SL g2119 ( 
.A(n_2090),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_2083),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2068),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2062),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2083),
.B(n_2009),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2071),
.B(n_2031),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2062),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2067),
.Y(n_2126)
);

INVxp67_ASAP7_75t_SL g2127 ( 
.A(n_2081),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2089),
.B(n_2031),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2083),
.B(n_2044),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2070),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2065),
.B(n_2027),
.Y(n_2131)
);

OAI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2085),
.A2(n_1939),
.B1(n_1935),
.B2(n_1900),
.Y(n_2132)
);

NAND2x1p5_ASAP7_75t_L g2133 ( 
.A(n_2094),
.B(n_1798),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2073),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2072),
.B(n_2030),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2068),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2074),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_2086),
.B(n_2030),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2066),
.B(n_2044),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2082),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2098),
.B(n_2036),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2105),
.B(n_2029),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2092),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_2100),
.Y(n_2144)
);

O2A1O1Ixp33_ASAP7_75t_L g2145 ( 
.A1(n_2093),
.A2(n_2029),
.B(n_2007),
.C(n_2059),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2101),
.B(n_2036),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2075),
.B(n_2088),
.Y(n_2147)
);

NOR2x1_ASAP7_75t_L g2148 ( 
.A(n_2064),
.B(n_1793),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2075),
.A2(n_1793),
.B(n_1968),
.Y(n_2149)
);

AND2x4_ASAP7_75t_SL g2150 ( 
.A(n_2063),
.B(n_2054),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2097),
.B(n_2006),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2077),
.B(n_2054),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2077),
.B(n_2054),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2078),
.B(n_2061),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2099),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_L g2156 ( 
.A(n_2081),
.B(n_1936),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2087),
.B(n_2061),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2116),
.B(n_2054),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2102),
.Y(n_2159)
);

AOI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_2127),
.A2(n_2104),
.B(n_2107),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2129),
.Y(n_2161)
);

INVxp67_ASAP7_75t_L g2162 ( 
.A(n_2144),
.Y(n_2162)
);

O2A1O1Ixp33_ASAP7_75t_SL g2163 ( 
.A1(n_2149),
.A2(n_2100),
.B(n_2106),
.C(n_2113),
.Y(n_2163)
);

NAND4xp25_ASAP7_75t_L g2164 ( 
.A(n_2147),
.B(n_2064),
.C(n_2107),
.D(n_2117),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_2145),
.A2(n_2104),
.B(n_2106),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_2124),
.A2(n_2117),
.B1(n_2084),
.B2(n_2118),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2139),
.B(n_2094),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_SL g2168 ( 
.A(n_2132),
.B(n_2109),
.C(n_2115),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2122),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_2156),
.A2(n_2063),
.B1(n_2096),
.B2(n_2084),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2156),
.A2(n_2096),
.B1(n_2116),
.B2(n_2095),
.C(n_2109),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2150),
.Y(n_2172)
);

AOI32xp33_ASAP7_75t_L g2173 ( 
.A1(n_2128),
.A2(n_2084),
.A3(n_2108),
.B1(n_2041),
.B2(n_2024),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_2120),
.Y(n_2174)
);

OAI21xp33_ASAP7_75t_L g2175 ( 
.A1(n_2129),
.A2(n_1928),
.B(n_1927),
.Y(n_2175)
);

O2A1O1Ixp33_ASAP7_75t_L g2176 ( 
.A1(n_2119),
.A2(n_2148),
.B(n_2151),
.C(n_2125),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2121),
.B(n_2114),
.Y(n_2177)
);

AOI221xp5_ASAP7_75t_L g2178 ( 
.A1(n_2120),
.A2(n_2112),
.B1(n_2111),
.B2(n_2110),
.C(n_2103),
.Y(n_2178)
);

AOI221x1_ASAP7_75t_L g2179 ( 
.A1(n_2121),
.A2(n_2114),
.B1(n_1965),
.B2(n_2069),
.C(n_1994),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2126),
.Y(n_2180)
);

NAND3x1_ASAP7_75t_L g2181 ( 
.A(n_2158),
.B(n_1864),
.C(n_1795),
.Y(n_2181)
);

OAI221xp5_ASAP7_75t_L g2182 ( 
.A1(n_2133),
.A2(n_1941),
.B1(n_1983),
.B2(n_1896),
.C(n_2050),
.Y(n_2182)
);

OAI21xp33_ASAP7_75t_SL g2183 ( 
.A1(n_2158),
.A2(n_2123),
.B(n_2152),
.Y(n_2183)
);

NAND4xp25_ASAP7_75t_L g2184 ( 
.A(n_2138),
.B(n_1801),
.C(n_1837),
.D(n_1830),
.Y(n_2184)
);

INVxp67_ASAP7_75t_SL g2185 ( 
.A(n_2133),
.Y(n_2185)
);

AOI21xp33_ASAP7_75t_L g2186 ( 
.A1(n_2142),
.A2(n_1968),
.B(n_1985),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2131),
.B(n_2135),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2130),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2131),
.B(n_2080),
.Y(n_2189)
);

NAND2x1p5_ASAP7_75t_L g2190 ( 
.A(n_2177),
.B(n_1801),
.Y(n_2190)
);

O2A1O1Ixp33_ASAP7_75t_L g2191 ( 
.A1(n_2163),
.A2(n_2159),
.B(n_2134),
.C(n_2155),
.Y(n_2191)
);

OAI322xp33_ASAP7_75t_L g2192 ( 
.A1(n_2165),
.A2(n_2136),
.A3(n_2137),
.B1(n_2140),
.B2(n_2143),
.C1(n_2135),
.C2(n_2146),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2162),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2174),
.B(n_2142),
.Y(n_2194)
);

AOI211xp5_ASAP7_75t_L g2195 ( 
.A1(n_2164),
.A2(n_2123),
.B(n_2152),
.C(n_2153),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2164),
.A2(n_2153),
.B1(n_2150),
.B2(n_2141),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2187),
.Y(n_2197)
);

OAI321xp33_ASAP7_75t_L g2198 ( 
.A1(n_2171),
.A2(n_2136),
.A3(n_2146),
.B1(n_2141),
.B2(n_2154),
.C(n_2157),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2176),
.A2(n_2157),
.B(n_2154),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_SL g2200 ( 
.A(n_2167),
.B(n_2060),
.C(n_2050),
.Y(n_2200)
);

A2O1A1Ixp33_ASAP7_75t_L g2201 ( 
.A1(n_2160),
.A2(n_2053),
.B(n_2059),
.C(n_2028),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2169),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2161),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_2170),
.B(n_2053),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2180),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2166),
.B(n_2091),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2172),
.B(n_2076),
.Y(n_2207)
);

OAI322xp33_ASAP7_75t_L g2208 ( 
.A1(n_2188),
.A2(n_2060),
.A3(n_2045),
.B1(n_2047),
.B2(n_2051),
.C1(n_2037),
.C2(n_1942),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2189),
.Y(n_2209)
);

OAI21xp33_ASAP7_75t_L g2210 ( 
.A1(n_2168),
.A2(n_1918),
.B(n_1899),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2183),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2184),
.B(n_2079),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_SL g2213 ( 
.A1(n_2182),
.A2(n_1968),
.B1(n_1899),
.B2(n_1918),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2197),
.B(n_2178),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2209),
.B(n_2173),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2211),
.B(n_2184),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2207),
.B(n_2195),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2194),
.B(n_2185),
.Y(n_2218)
);

INVxp67_ASAP7_75t_SL g2219 ( 
.A(n_2190),
.Y(n_2219)
);

AOI222xp33_ASAP7_75t_L g2220 ( 
.A1(n_2193),
.A2(n_2175),
.B1(n_2179),
.B2(n_2041),
.C1(n_2024),
.C2(n_2042),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2192),
.A2(n_2186),
.B1(n_2041),
.B2(n_2042),
.C(n_2024),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2203),
.B(n_2042),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_2190),
.B(n_2181),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2202),
.Y(n_2224)
);

OAI32xp33_ASAP7_75t_L g2225 ( 
.A1(n_2190),
.A2(n_2051),
.A3(n_2037),
.B1(n_2047),
.B2(n_2045),
.Y(n_2225)
);

XOR2x1_ASAP7_75t_L g2226 ( 
.A(n_2205),
.B(n_1810),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2207),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2212),
.Y(n_2228)
);

XNOR2x1_ASAP7_75t_L g2229 ( 
.A(n_2206),
.B(n_1810),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2227),
.Y(n_2230)
);

AOI211xp5_ASAP7_75t_L g2231 ( 
.A1(n_2214),
.A2(n_2201),
.B(n_2198),
.C(n_2191),
.Y(n_2231)
);

NAND3xp33_ASAP7_75t_SL g2232 ( 
.A(n_2214),
.B(n_2201),
.C(n_2199),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2222),
.Y(n_2233)
);

NOR3xp33_ASAP7_75t_L g2234 ( 
.A(n_2228),
.B(n_2204),
.C(n_2210),
.Y(n_2234)
);

AOI211x1_ASAP7_75t_L g2235 ( 
.A1(n_2215),
.A2(n_2204),
.B(n_2196),
.C(n_2200),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2218),
.Y(n_2236)
);

NOR3xp33_ASAP7_75t_L g2237 ( 
.A(n_2216),
.B(n_2213),
.C(n_2208),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2217),
.B(n_2000),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2224),
.Y(n_2239)
);

NAND4xp25_ASAP7_75t_L g2240 ( 
.A(n_2220),
.B(n_1865),
.C(n_1935),
.D(n_1900),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2229),
.B(n_2000),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2238),
.B(n_2219),
.Y(n_2242)
);

AOI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2232),
.A2(n_2221),
.B1(n_2225),
.B2(n_2223),
.C(n_2220),
.Y(n_2243)
);

OAI221xp5_ASAP7_75t_SL g2244 ( 
.A1(n_2231),
.A2(n_2226),
.B1(n_1825),
.B2(n_2051),
.C(n_2037),
.Y(n_2244)
);

XNOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2236),
.B(n_1969),
.Y(n_2245)
);

AOI222xp33_ASAP7_75t_L g2246 ( 
.A1(n_2232),
.A2(n_1977),
.B1(n_1918),
.B2(n_1899),
.C1(n_1929),
.C2(n_1947),
.Y(n_2246)
);

NAND4xp25_ASAP7_75t_SL g2247 ( 
.A(n_2237),
.B(n_1872),
.C(n_1969),
.D(n_1971),
.Y(n_2247)
);

AOI211xp5_ASAP7_75t_L g2248 ( 
.A1(n_2234),
.A2(n_1786),
.B(n_1784),
.C(n_1787),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2242),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2245),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2244),
.Y(n_2251)
);

INVx1_ASAP7_75t_SL g2252 ( 
.A(n_2248),
.Y(n_2252)
);

INVxp33_ASAP7_75t_L g2253 ( 
.A(n_2243),
.Y(n_2253)
);

OAI211xp5_ASAP7_75t_L g2254 ( 
.A1(n_2246),
.A2(n_2235),
.B(n_2230),
.C(n_2233),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2247),
.B(n_2239),
.Y(n_2255)
);

NAND4xp75_ASAP7_75t_L g2256 ( 
.A(n_2249),
.B(n_2241),
.C(n_2240),
.D(n_1984),
.Y(n_2256)
);

NAND4xp75_ASAP7_75t_L g2257 ( 
.A(n_2250),
.B(n_1984),
.C(n_2043),
.D(n_2048),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_2252),
.B(n_2023),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2254),
.B(n_2023),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2255),
.B(n_2043),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2252),
.Y(n_2261)
);

NAND3xp33_ASAP7_75t_L g2262 ( 
.A(n_2261),
.B(n_2253),
.C(n_2251),
.Y(n_2262)
);

NAND3xp33_ASAP7_75t_L g2263 ( 
.A(n_2259),
.B(n_1771),
.C(n_2056),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2258),
.B(n_2023),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2262),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2265),
.A2(n_2256),
.B1(n_2257),
.B2(n_2260),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2266),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2266),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2268),
.Y(n_2269)
);

AOI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2267),
.A2(n_2264),
.B1(n_2263),
.B2(n_2023),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2269),
.Y(n_2271)
);

AOI221xp5_ASAP7_75t_L g2272 ( 
.A1(n_2270),
.A2(n_2048),
.B1(n_2056),
.B2(n_2015),
.C(n_2018),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2271),
.A2(n_2015),
.B1(n_2018),
.B2(n_2020),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2273),
.Y(n_2274)
);

XNOR2xp5_ASAP7_75t_L g2275 ( 
.A(n_2274),
.B(n_2272),
.Y(n_2275)
);

OAI221xp5_ASAP7_75t_R g2276 ( 
.A1(n_2275),
.A2(n_1673),
.B1(n_2015),
.B2(n_2018),
.C(n_2020),
.Y(n_2276)
);

AOI211xp5_ASAP7_75t_L g2277 ( 
.A1(n_2276),
.A2(n_1784),
.B(n_1786),
.C(n_2056),
.Y(n_2277)
);


endmodule