module fake_jpeg_23589_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_56;
wire n_131;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_40),
.B(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_25),
.B(n_0),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_32),
.C(n_31),
.Y(n_74)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_26),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_55),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_34),
.B1(n_20),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_62),
.B1(n_81),
.B2(n_23),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_17),
.B(n_22),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_74),
.B(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_19),
.B1(n_20),
.B2(n_27),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_4),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_20),
.B1(n_35),
.B2(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_35),
.B1(n_33),
.B2(n_32),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_4),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_29),
.B1(n_17),
.B2(n_3),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_82),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_40),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_84),
.B(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_94),
.B1(n_5),
.B2(n_7),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_67),
.B(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_16),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_2),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_79),
.B1(n_68),
.B2(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_82),
.B1(n_79),
.B2(n_49),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_5),
.B(n_7),
.Y(n_123)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_52),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_118),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_82),
.B(n_79),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_86),
.B(n_84),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_86),
.A3(n_110),
.B1(n_96),
.B2(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_53),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_53),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_127),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_102),
.B1(n_114),
.B2(n_87),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_72),
.B1(n_49),
.B2(n_57),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_128),
.B1(n_99),
.B2(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_77),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_75),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_57),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_93),
.B(n_5),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_110),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_78),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_70),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_145),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_87),
.B(n_72),
.C(n_71),
.Y(n_142)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_155),
.B1(n_163),
.B2(n_135),
.C(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_92),
.B(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_153),
.B(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_116),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_8),
.C(n_9),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_87),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_164),
.B1(n_121),
.B2(n_115),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_100),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_8),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_107),
.B(n_109),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_96),
.B1(n_55),
.B2(n_58),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_173),
.B1(n_163),
.B2(n_155),
.C(n_142),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_113),
.B1(n_118),
.B2(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_174),
.B1(n_175),
.B2(n_151),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_180),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_8),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_112),
.B1(n_70),
.B2(n_88),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_112),
.B1(n_88),
.B2(n_91),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_164),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_138),
.C(n_124),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_161),
.C(n_149),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_124),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_177),
.B(n_153),
.C(n_143),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_198),
.C(n_186),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_190),
.B(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_143),
.B1(n_153),
.B2(n_160),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_179),
.C(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_166),
.C(n_168),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_169),
.Y(n_203)
);

OAI322xp33_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_152),
.A3(n_158),
.B1(n_147),
.B2(n_142),
.C1(n_145),
.C2(n_144),
.Y(n_197)
);

OAI322xp33_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_172),
.A3(n_167),
.B1(n_165),
.B2(n_169),
.C1(n_178),
.C2(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

BUFx4f_ASAP7_75t_SL g211 ( 
.A(n_199),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_203),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_185),
.B1(n_191),
.B2(n_205),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_182),
.B(n_184),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_208),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_170),
.C(n_140),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_140),
.C(n_168),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_189),
.B1(n_193),
.B2(n_191),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_216),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_167),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_190),
.B(n_180),
.C(n_188),
.Y(n_215)
);

OAI31xp33_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_211),
.A3(n_184),
.B(n_187),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_221),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_194),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_9),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_207),
.C(n_200),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_124),
.B(n_130),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_228),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_213),
.Y(n_232)
);

OAI221xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_215),
.B1(n_216),
.B2(n_220),
.C(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_230),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_213),
.B1(n_130),
.B2(n_131),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_232),
.A2(n_225),
.B1(n_228),
.B2(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_130),
.C(n_131),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_237),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_224),
.B(n_226),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_235),
.B(n_12),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_239),
.C(n_15),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_11),
.CI(n_12),
.CON(n_239),
.SN(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_11),
.B(n_14),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);


endmodule