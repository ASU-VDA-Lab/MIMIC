module fake_jpeg_7202_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_35),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_21),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_29),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_16),
.C(n_26),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_34),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_27),
.B1(n_23),
.B2(n_21),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_12),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_33),
.B1(n_25),
.B2(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_25),
.B1(n_33),
.B2(n_31),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_35),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_28),
.B1(n_34),
.B2(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_107),
.B1(n_59),
.B2(n_57),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_76),
.B(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_108),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_81),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_29),
.B(n_17),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_41),
.B(n_22),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_96),
.B1(n_104),
.B2(n_109),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_48),
.B(n_66),
.C(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_35),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g128 ( 
.A(n_90),
.Y(n_128)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_17),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_12),
.B(n_15),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g138 ( 
.A(n_94),
.B(n_100),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_17),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_101),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_22),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_106),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_22),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_27),
.B1(n_45),
.B2(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_29),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_44),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_122),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_41),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_100),
.B(n_108),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_57),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_101),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_36),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_44),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_105),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_80),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_141),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_148),
.B(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_102),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_143),
.B(n_157),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_145),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_151),
.C(n_43),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_155),
.B(n_126),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_73),
.B(n_81),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_90),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_133),
.B1(n_116),
.B2(n_122),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_154),
.B1(n_158),
.B2(n_59),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_83),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_153),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_83),
.B(n_78),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_86),
.B1(n_99),
.B2(n_91),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_83),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_117),
.B(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_165),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_36),
.A3(n_45),
.B1(n_44),
.B2(n_22),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_153),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_36),
.A3(n_45),
.B1(n_22),
.B2(n_43),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_172),
.A2(n_170),
.B1(n_168),
.B2(n_140),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_133),
.B1(n_122),
.B2(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_186),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_120),
.B1(n_112),
.B2(n_125),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_112),
.B1(n_115),
.B2(n_123),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_189),
.B(n_161),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_43),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_43),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_159),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_157),
.B1(n_139),
.B2(n_141),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_117),
.B1(n_129),
.B2(n_137),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_22),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_63),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_43),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_143),
.A2(n_129),
.B1(n_96),
.B2(n_36),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_144),
.B(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_63),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_155),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_129),
.B1(n_45),
.B2(n_36),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_203),
.A2(n_204),
.B1(n_84),
.B2(n_45),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_45),
.B1(n_43),
.B2(n_67),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_163),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_220),
.Y(n_251)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_185),
.B1(n_186),
.B2(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_208),
.A2(n_211),
.B(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_188),
.B(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_169),
.B(n_1),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_226),
.Y(n_244)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_127),
.C(n_74),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

BUFx12f_ASAP7_75t_SL g228 ( 
.A(n_193),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_231),
.B1(n_190),
.B2(n_175),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_74),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_220),
.B1(n_217),
.B2(n_226),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_239),
.B1(n_242),
.B2(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_190),
.B1(n_175),
.B2(n_176),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_178),
.B1(n_172),
.B2(n_174),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_247),
.B1(n_230),
.B2(n_219),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_196),
.C(n_184),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_213),
.C(n_209),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_177),
.B1(n_194),
.B2(n_191),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_194),
.B1(n_201),
.B2(n_187),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_197),
.B1(n_202),
.B2(n_195),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_200),
.B1(n_183),
.B2(n_204),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_252),
.B1(n_254),
.B2(n_243),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_127),
.B1(n_130),
.B2(n_45),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_215),
.A2(n_127),
.B1(n_130),
.B2(n_74),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_262),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_209),
.C(n_225),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_259),
.B(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_253),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_207),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_205),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_268),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_207),
.C(n_224),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_237),
.B1(n_245),
.B2(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_67),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_238),
.A2(n_223),
.B1(n_9),
.B2(n_10),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_257),
.B(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_233),
.B1(n_239),
.B2(n_252),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_249),
.B(n_232),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_249),
.B(n_240),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_253),
.B1(n_246),
.B2(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_273),
.B(n_268),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_280),
.A2(n_258),
.B(n_1),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_0),
.Y(n_301)
);

INVx11_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_273),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_260),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_88),
.B1(n_1),
.B2(n_2),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_260),
.C(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_290),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_271),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

OAI21x1_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_259),
.B(n_262),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_281),
.B1(n_286),
.B2(n_279),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_8),
.B(n_15),
.Y(n_297)
);

BUFx12f_ASAP7_75t_SL g298 ( 
.A(n_287),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_283),
.B(n_8),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_43),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_284),
.B1(n_285),
.B2(n_282),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_301),
.B1(n_2),
.B2(n_3),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_307),
.C(n_311),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_288),
.B1(n_275),
.B2(n_278),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_296),
.B(n_10),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_283),
.C(n_63),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_294),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_7),
.C(n_13),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_7),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_318),
.A3(n_313),
.B1(n_304),
.B2(n_13),
.C1(n_11),
.C2(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_13),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_321),
.B(n_2),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_306),
.A3(n_311),
.B1(n_302),
.B2(n_63),
.C1(n_1),
.C2(n_4),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_3),
.B(n_4),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_3),
.Y(n_327)
);


endmodule