module fake_netlist_6_2490_n_3618 (n_992, n_52, n_591, n_435, n_1115, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_1079, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_1103, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_1061, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_1044, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_1072, n_677, n_969, n_988, n_805, n_396, n_495, n_1065, n_815, n_350, n_1100, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_1128, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_1071, n_628, n_1067, n_883, n_557, n_823, n_1132, n_349, n_643, n_233, n_617, n_698, n_898, n_1074, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_1138, n_893, n_214, n_925, n_485, n_1099, n_67, n_15, n_1026, n_443, n_1101, n_246, n_892, n_768, n_1097, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_1130, n_59, n_181, n_1127, n_182, n_238, n_1095, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_1120, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_1139, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_1105, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_1140, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_1114, n_56, n_763, n_1057, n_1147, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_1143, n_536, n_895, n_1126, n_866, n_622, n_147, n_191, n_340, n_710, n_1108, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_1119, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_1056, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_1116, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_1094, n_494, n_539, n_493, n_397, n_155, n_1022, n_1083, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_1112, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_1117, n_1087, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_1049, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1043, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_1088, n_708, n_196, n_919, n_1081, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_1084, n_107, n_1104, n_907, n_854, n_6, n_1058, n_417, n_14, n_446, n_498, n_662, n_1122, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_1109, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_1148, n_293, n_1054, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_1070, n_1085, n_232, n_650, n_998, n_16, n_1046, n_163, n_717, n_46, n_1145, n_330, n_771, n_1121, n_470, n_475, n_924, n_1102, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1073, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_1062, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_1090, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_1142, n_503, n_716, n_152, n_623, n_1048, n_1123, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_1078, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_1137, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_1144, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_1068, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_1075, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_1110, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_1133, n_635, n_95, n_787, n_311, n_10, n_1064, n_403, n_1080, n_723, n_253, n_634, n_1051, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_1141, n_1146, n_249, n_201, n_386, n_764, n_1039, n_556, n_159, n_1034, n_1086, n_1066, n_157, n_162, n_692, n_733, n_754, n_1136, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_1125, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_1107, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_1092, n_441, n_221, n_811, n_882, n_1060, n_444, n_586, n_423, n_146, n_737, n_318, n_1111, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_1053, n_530, n_277, n_520, n_1029, n_418, n_1093, n_113, n_618, n_1055, n_790, n_1106, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_1069, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1047, n_1010, n_355, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_1131, n_54, n_1052, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_1045, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_1089, n_1135, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_1096, n_1063, n_729, n_1091, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_1124, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_1059, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_1077, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_1082, n_259, n_177, n_1113, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_1098, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_1050, n_379, n_170, n_778, n_1025, n_1134, n_332, n_891, n_336, n_12, n_398, n_410, n_1129, n_566, n_554, n_602, n_1013, n_1023, n_1076, n_1118, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_3618);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1115;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_1079;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_1103;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_1061;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_1044;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_1072;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_1065;
input n_815;
input n_350;
input n_1100;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_1128;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_1071;
input n_628;
input n_1067;
input n_883;
input n_557;
input n_823;
input n_1132;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1074;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_1138;
input n_893;
input n_214;
input n_925;
input n_485;
input n_1099;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_1101;
input n_246;
input n_892;
input n_768;
input n_1097;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_1130;
input n_59;
input n_181;
input n_1127;
input n_182;
input n_238;
input n_1095;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_1120;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_1139;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_1105;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_1140;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1057;
input n_1147;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_1143;
input n_536;
input n_895;
input n_1126;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_1108;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_1119;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_1116;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_1094;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_1083;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_1112;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_1117;
input n_1087;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_1049;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1043;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_1088;
input n_708;
input n_196;
input n_919;
input n_1081;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_1084;
input n_107;
input n_1104;
input n_907;
input n_854;
input n_6;
input n_1058;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_1122;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_1109;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_1148;
input n_293;
input n_1054;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_1070;
input n_1085;
input n_232;
input n_650;
input n_998;
input n_16;
input n_1046;
input n_163;
input n_717;
input n_46;
input n_1145;
input n_330;
input n_771;
input n_1121;
input n_470;
input n_475;
input n_924;
input n_1102;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1073;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_1062;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_1090;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_1142;
input n_503;
input n_716;
input n_152;
input n_623;
input n_1048;
input n_1123;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_1078;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_1137;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_1144;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_1068;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_1075;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_1110;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_1064;
input n_403;
input n_1080;
input n_723;
input n_253;
input n_634;
input n_1051;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_1141;
input n_1146;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_556;
input n_159;
input n_1034;
input n_1086;
input n_1066;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_1136;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_1125;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_1107;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_1092;
input n_441;
input n_221;
input n_811;
input n_882;
input n_1060;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_1111;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_1053;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_1093;
input n_113;
input n_618;
input n_1055;
input n_790;
input n_1106;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_1069;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1047;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_1131;
input n_54;
input n_1052;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_1045;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_1089;
input n_1135;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_1096;
input n_1063;
input n_729;
input n_1091;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_1124;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_1059;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_1077;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_1082;
input n_259;
input n_177;
input n_1113;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_1098;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_1050;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_1134;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_1129;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_3618;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1581;
wire n_1237;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3251;
wire n_3316;
wire n_2212;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1471;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_3368;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_1658;
wire n_2593;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_1193;
wire n_1967;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_1302;
wire n_1599;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_1873;
wire n_3518;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_2068;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3247;
wire n_3069;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_1214;
wire n_2347;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_3415;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_3510;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3500;
wire n_3526;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_2271;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_3209;
wire n_3450;
wire n_2622;
wire n_1858;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2750;
wire n_2558;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1627;
wire n_1295;
wire n_1164;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2684;
wire n_2712;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_1952;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_1932;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_3179;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_2537;
wire n_2554;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3537;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2667;
wire n_2539;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3325;
wire n_3203;
wire n_2238;
wire n_2368;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_2849;
wire n_1774;
wire n_1475;
wire n_3103;
wire n_1398;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_1837;
wire n_1314;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_3244;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_3306;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_2329;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_2990;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_2249;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3284;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3205;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_2315;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_3566;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_2201;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3276;
wire n_3194;
wire n_1934;
wire n_3250;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_3548;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3550;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_2412;
wire n_1997;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_2305;
wire n_2120;
wire n_2050;
wire n_1472;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3379;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1741;
wire n_1746;
wire n_1325;
wire n_1949;
wire n_3398;
wire n_3524;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_2516;
wire n_3391;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_2949;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_2969;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_1785;
wire n_1848;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_1737;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_3584;
wire n_3486;
wire n_2649;
wire n_2721;
wire n_3556;
wire n_2034;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_1821;
wire n_1537;
wire n_1500;
wire n_2205;
wire n_3204;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3290;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1156;
wire n_1362;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_2071;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1194;
wire n_3374;
wire n_2742;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3330;
wire n_1479;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_3444;
wire n_2553;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_2512;
wire n_3433;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_1322;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_3504;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx14_ASAP7_75t_R g1149 ( 
.A(n_954),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_873),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_860),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_109),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_815),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_502),
.Y(n_1154)
);

CKINVDCx16_ASAP7_75t_R g1155 ( 
.A(n_844),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1047),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_552),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_137),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_854),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_653),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_659),
.Y(n_1161)
);

CKINVDCx16_ASAP7_75t_R g1162 ( 
.A(n_1087),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1017),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_833),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_402),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_866),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_863),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_730),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_904),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_834),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_202),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_482),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1141),
.B(n_440),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_267),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_417),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_858),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1118),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1009),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_908),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_823),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_752),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1014),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_398),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_982),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_789),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_593),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_172),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_753),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_419),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_252),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_498),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_903),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_138),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_669),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_485),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_211),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_674),
.Y(n_1198)
);

BUFx2_ASAP7_75t_SL g1199 ( 
.A(n_841),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_968),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_731),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_494),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_724),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_908),
.B(n_453),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_185),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_969),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_253),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_754),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_163),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_864),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_385),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_60),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_402),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_4),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_667),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_161),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_722),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_986),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_846),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_553),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_216),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_323),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_244),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_632),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_876),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_381),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1095),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_959),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_373),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_11),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_967),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_834),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_541),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_903),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_64),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_727),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_405),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_329),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_61),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_313),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_297),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1114),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_89),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_127),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_689),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_907),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1115),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_201),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_394),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_862),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_743),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_366),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_548),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1025),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_316),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_56),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_513),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1027),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_217),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1016),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_732),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_630),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1134),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_381),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_290),
.B(n_1042),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_297),
.Y(n_1266)
);

CKINVDCx16_ASAP7_75t_R g1267 ( 
.A(n_577),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_305),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_677),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_844),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_396),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_154),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_418),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_449),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_302),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_217),
.Y(n_1276)
);

CKINVDCx16_ASAP7_75t_R g1277 ( 
.A(n_891),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_524),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_840),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_219),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_463),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_712),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_175),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_42),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_790),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_934),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_880),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_565),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_663),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_231),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_698),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_119),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_693),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_347),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1073),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_881),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_394),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_857),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_758),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1116),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_360),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_460),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_751),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_475),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_861),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_819),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_871),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_25),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_345),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_233),
.Y(n_1310)
);

INVxp33_ASAP7_75t_L g1311 ( 
.A(n_617),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_60),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1000),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_504),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_594),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_694),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_816),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_917),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_27),
.B(n_891),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_52),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_852),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_845),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1061),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1012),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_804),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_35),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_515),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_89),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_820),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1102),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_632),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_502),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_816),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_784),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_195),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_438),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_140),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_485),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1132),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_392),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_185),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1060),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_826),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_938),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_870),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_721),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1048),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_757),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_765),
.B(n_536),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_225),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_349),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_877),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_717),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_824),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_110),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_878),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_615),
.B(n_296),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_780),
.Y(n_1358)
);

NOR2xp67_ASAP7_75t_L g1359 ( 
.A(n_252),
.B(n_101),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_652),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_433),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_126),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_612),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_655),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_991),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_874),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1138),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_132),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_680),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_215),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_745),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_831),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_616),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1020),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_514),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_556),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_607),
.Y(n_1377)
);

BUFx10_ASAP7_75t_L g1378 ( 
.A(n_272),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_720),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_371),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_702),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_91),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_661),
.Y(n_1383)
);

BUFx8_ASAP7_75t_SL g1384 ( 
.A(n_424),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1136),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1049),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_885),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_517),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_851),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_575),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_482),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_813),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1023),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_197),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_872),
.Y(n_1395)
);

BUFx10_ASAP7_75t_L g1396 ( 
.A(n_835),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_25),
.Y(n_1397)
);

INVxp67_ASAP7_75t_SL g1398 ( 
.A(n_842),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_679),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_166),
.Y(n_1400)
);

CKINVDCx16_ASAP7_75t_R g1401 ( 
.A(n_607),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_567),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_822),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_355),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_970),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_856),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_451),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_125),
.Y(n_1408)
);

BUFx10_ASAP7_75t_L g1409 ( 
.A(n_323),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_881),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_732),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_108),
.Y(n_1412)
);

CKINVDCx16_ASAP7_75t_R g1413 ( 
.A(n_1090),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_692),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1065),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_509),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_345),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_935),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_298),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_930),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1098),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1113),
.B(n_1004),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_818),
.B(n_726),
.Y(n_1423)
);

BUFx5_ASAP7_75t_L g1424 ( 
.A(n_957),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_534),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_500),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_288),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_915),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_985),
.B(n_830),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1097),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_622),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_998),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_1026),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_120),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_647),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_948),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_18),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_755),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_829),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_20),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_879),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_222),
.Y(n_1442)
);

CKINVDCx16_ASAP7_75t_R g1443 ( 
.A(n_1024),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_855),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1133),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_572),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_236),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_918),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_636),
.Y(n_1449)
);

CKINVDCx16_ASAP7_75t_R g1450 ( 
.A(n_403),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_774),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_955),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_30),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_868),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_396),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_836),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_222),
.Y(n_1457)
);

CKINVDCx16_ASAP7_75t_R g1458 ( 
.A(n_3),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_907),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_843),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_414),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_576),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1033),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_518),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_711),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_233),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_850),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_617),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_535),
.B(n_119),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_480),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_649),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_261),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_45),
.Y(n_1473)
);

CKINVDCx14_ASAP7_75t_R g1474 ( 
.A(n_856),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_475),
.Y(n_1475)
);

BUFx10_ASAP7_75t_L g1476 ( 
.A(n_867),
.Y(n_1476)
);

INVxp33_ASAP7_75t_L g1477 ( 
.A(n_424),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_14),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_224),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_167),
.Y(n_1480)
);

CKINVDCx16_ASAP7_75t_R g1481 ( 
.A(n_730),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_118),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_407),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_429),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_884),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_976),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1068),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_868),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_133),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_145),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_699),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_496),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_357),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_937),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_700),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_646),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1001),
.B(n_1037),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_76),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_960),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_805),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_369),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1063),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_788),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_131),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_88),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_279),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_567),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_247),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_165),
.B(n_801),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_9),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_898),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_512),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_521),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_870),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_183),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_154),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_360),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1021),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_445),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_418),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_931),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_993),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_852),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_581),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_555),
.Y(n_1526)
);

CKINVDCx16_ASAP7_75t_R g1527 ( 
.A(n_882),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_135),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_615),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_675),
.Y(n_1530)
);

BUFx5_ASAP7_75t_L g1531 ( 
.A(n_601),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1106),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_624),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1019),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_128),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_875),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_825),
.B(n_564),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_563),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_540),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_878),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_403),
.Y(n_1541)
);

INVxp33_ASAP7_75t_L g1542 ( 
.A(n_210),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_906),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_633),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_926),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_328),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_979),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_839),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_450),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_112),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_341),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_810),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_977),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1062),
.Y(n_1554)
);

BUFx5_ASAP7_75t_L g1555 ( 
.A(n_274),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_848),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_853),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_460),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_832),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_544),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_506),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_382),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_459),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_363),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_9),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_32),
.Y(n_1566)
);

CKINVDCx16_ASAP7_75t_R g1567 ( 
.A(n_92),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_122),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_865),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_7),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_7),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_434),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_821),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_348),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_740),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_827),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_549),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_849),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1137),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_591),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_21),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_88),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_584),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_404),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_919),
.Y(n_1585)
);

CKINVDCx14_ASAP7_75t_R g1586 ( 
.A(n_859),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_899),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_643),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_883),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_837),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_544),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_888),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_850),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_642),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_543),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_847),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_838),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_258),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_815),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_34),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_192),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1081),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_313),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_430),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_455),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_946),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_650),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_522),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_133),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_672),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_869),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_828),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_384),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_335),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_175),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_456),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_817),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_390),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1531),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1531),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1193),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1531),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1198),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1198),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1236),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1384),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1531),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1531),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1155),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1163),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1198),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1474),
.B(n_0),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1555),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1218),
.Y(n_1634)
);

AND2x6_ASAP7_75t_L g1635 ( 
.A(n_1423),
.B(n_920),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1554),
.B(n_1),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1202),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1242),
.A2(n_922),
.B(n_921),
.Y(n_1638)
);

CKINVDCx6p67_ASAP7_75t_R g1639 ( 
.A(n_1248),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1286),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1586),
.B(n_0),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1165),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1300),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1555),
.Y(n_1644)
);

INVx5_ASAP7_75t_L g1645 ( 
.A(n_1165),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1156),
.A2(n_924),
.B(n_923),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1579),
.A2(n_927),
.B(n_925),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1555),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1165),
.Y(n_1649)
);

INVx5_ASAP7_75t_L g1650 ( 
.A(n_1534),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1555),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1202),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1555),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1202),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1238),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1205),
.Y(n_1656)
);

BUFx8_ASAP7_75t_SL g1657 ( 
.A(n_1257),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1152),
.Y(n_1658)
);

INVx6_ASAP7_75t_L g1659 ( 
.A(n_1282),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1519),
.B(n_1),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1152),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1522),
.B(n_2),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1553),
.B(n_2),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1205),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1282),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1205),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1283),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1274),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1149),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1618),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1534),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1178),
.A2(n_929),
.B(n_928),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1274),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1173),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1301),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1185),
.B(n_6),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1179),
.A2(n_933),
.B(n_932),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1183),
.A2(n_939),
.B(n_936),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1618),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1162),
.B(n_8),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1274),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1309),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1368),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1337),
.B(n_10),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1309),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1390),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1309),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1322),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1267),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1206),
.A2(n_941),
.B(n_940),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1493),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1322),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1228),
.B(n_10),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1277),
.B(n_11),
.Y(n_1695)
);

INVx6_ASAP7_75t_L g1696 ( 
.A(n_1327),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1341),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1413),
.B(n_12),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1322),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1352),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1231),
.B(n_12),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1352),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1352),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1362),
.Y(n_1704)
);

XOR2xp5_ASAP7_75t_L g1705 ( 
.A(n_1299),
.B(n_13),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1362),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1362),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1311),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1363),
.Y(n_1709)
);

NAND2xp33_ASAP7_75t_L g1710 ( 
.A(n_1349),
.B(n_15),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1327),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1363),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1363),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1516),
.Y(n_1714)
);

OAI22x1_ASAP7_75t_R g1715 ( 
.A1(n_1184),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1247),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1465),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1465),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1465),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1563),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1360),
.B(n_16),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1401),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1433),
.B(n_17),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1563),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1200),
.Y(n_1725)
);

AND2x2_ASAP7_75t_SL g1726 ( 
.A(n_1443),
.B(n_19),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1563),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1578),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1578),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1410),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1578),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1431),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1566),
.B(n_19),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1450),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1583),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1583),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1583),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1254),
.A2(n_943),
.B(n_942),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1258),
.B(n_20),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1424),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1260),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1560),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1477),
.B(n_1542),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1344),
.B(n_21),
.Y(n_1744)
);

AND2x6_ASAP7_75t_L g1745 ( 
.A(n_1534),
.B(n_944),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1365),
.B(n_22),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1604),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1458),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1378),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1623),
.Y(n_1750)
);

AND2x2_ASAP7_75t_SL g1751 ( 
.A(n_1726),
.B(n_1481),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1629),
.B(n_1527),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1641),
.B(n_1227),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_L g1754 ( 
.A(n_1681),
.B(n_1357),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1659),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1630),
.B(n_1265),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1623),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1624),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1624),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1631),
.Y(n_1760)
);

INVxp33_ASAP7_75t_L g1761 ( 
.A(n_1743),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1685),
.A2(n_1601),
.B1(n_1569),
.B2(n_1219),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1631),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1654),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1637),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1749),
.B(n_1550),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1634),
.B(n_1367),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1696),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1656),
.Y(n_1769)
);

BUFx10_ASAP7_75t_L g1770 ( 
.A(n_1666),
.Y(n_1770)
);

NOR2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1639),
.B(n_1469),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1690),
.B(n_1567),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1716),
.B(n_1385),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1660),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1722),
.B(n_1182),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1637),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1667),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1734),
.Y(n_1778)
);

INVx4_ASAP7_75t_L g1779 ( 
.A(n_1741),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1632),
.B(n_1174),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1725),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1671),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1711),
.B(n_1429),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1680),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1652),
.Y(n_1785)
);

BUFx8_ASAP7_75t_SL g1786 ( 
.A(n_1626),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1640),
.B(n_1386),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1683),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1730),
.B(n_1199),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1652),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1698),
.B(n_1393),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1723),
.B(n_1405),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1636),
.B(n_1509),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1748),
.A2(n_1537),
.B1(n_1594),
.B2(n_1172),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1693),
.Y(n_1795)
);

BUFx10_ASAP7_75t_L g1796 ( 
.A(n_1742),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1700),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1699),
.Y(n_1798)
);

INVx8_ASAP7_75t_L g1799 ( 
.A(n_1657),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1643),
.B(n_1418),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1702),
.Y(n_1801)
);

AOI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1619),
.A2(n_1445),
.B(n_1436),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1699),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1677),
.B(n_1448),
.Y(n_1804)
);

CKINVDCx16_ASAP7_75t_R g1805 ( 
.A(n_1687),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1721),
.A2(n_1317),
.B1(n_1403),
.B2(n_1216),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1709),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1704),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1714),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_R g1810 ( 
.A(n_1733),
.B(n_1646),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1706),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1709),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1745),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_SL g1814 ( 
.A(n_1747),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1713),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1668),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1713),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1707),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1717),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1712),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1719),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1720),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1717),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1727),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1645),
.B(n_1463),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1658),
.B(n_1203),
.Y(n_1826)
);

BUFx10_ASAP7_75t_L g1827 ( 
.A(n_1661),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1731),
.Y(n_1828)
);

BUFx10_ASAP7_75t_L g1829 ( 
.A(n_1663),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1718),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1621),
.Y(n_1831)
);

INVx8_ASAP7_75t_L g1832 ( 
.A(n_1635),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1718),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1831),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1761),
.B(n_1697),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1764),
.Y(n_1836)
);

INVx8_ASAP7_75t_L g1837 ( 
.A(n_1799),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1780),
.B(n_1664),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1753),
.B(n_1732),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1791),
.B(n_1792),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1767),
.B(n_1645),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1809),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1769),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1774),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1777),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1773),
.B(n_1756),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1804),
.B(n_1650),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1793),
.A2(n_1635),
.B1(n_1710),
.B2(n_1701),
.Y(n_1848)
);

INVx4_ASAP7_75t_L g1849 ( 
.A(n_1832),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1813),
.B(n_1650),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1762),
.B(n_1695),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1782),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1784),
.Y(n_1853)
);

OAI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1806),
.A2(n_1744),
.B(n_1739),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1788),
.B(n_1642),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1795),
.B(n_1649),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1797),
.B(n_1672),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1794),
.A2(n_1746),
.B1(n_1190),
.B2(n_1287),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1801),
.B(n_1694),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1808),
.B(n_1620),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1750),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1811),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1751),
.B(n_1313),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1805),
.B(n_1323),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1832),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1779),
.B(n_1625),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_SL g1867 ( 
.A(n_1816),
.B(n_1374),
.Y(n_1867)
);

O2A1O1Ixp33_ASAP7_75t_L g1868 ( 
.A1(n_1754),
.A2(n_1662),
.B(n_1708),
.C(n_1628),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1766),
.B(n_1263),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1775),
.B(n_1655),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1818),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1778),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1752),
.B(n_1676),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1820),
.B(n_1622),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1821),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1822),
.Y(n_1876)
);

AO221x1_ASAP7_75t_L g1877 ( 
.A1(n_1810),
.A2(n_1670),
.B1(n_1675),
.B2(n_1606),
.C(n_1153),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1796),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1772),
.B(n_1684),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_SL g1880 ( 
.A1(n_1789),
.A2(n_1194),
.B1(n_1273),
.B2(n_1211),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1824),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1828),
.B(n_1644),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1759),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1760),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1763),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1790),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1770),
.B(n_1295),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1798),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1787),
.B(n_1648),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1800),
.B(n_1651),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1781),
.Y(n_1891)
);

INVx4_ASAP7_75t_L g1892 ( 
.A(n_1814),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1825),
.B(n_1653),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1783),
.B(n_1692),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1789),
.B(n_1735),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1771),
.A2(n_1204),
.B1(n_1398),
.B2(n_1359),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1826),
.B(n_1627),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1803),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1799),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1826),
.B(n_1633),
.Y(n_1900)
);

INVx4_ASAP7_75t_L g1901 ( 
.A(n_1827),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1807),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1829),
.B(n_1724),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1817),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1823),
.B(n_1745),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1750),
.B(n_1724),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1830),
.B(n_1736),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1833),
.A2(n_1332),
.B1(n_1348),
.B2(n_1276),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1757),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1802),
.B(n_1740),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1765),
.B(n_1776),
.Y(n_1911)
);

CKINVDCx16_ASAP7_75t_R g1912 ( 
.A(n_1755),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1768),
.A2(n_1319),
.B1(n_1249),
.B2(n_1289),
.Y(n_1913)
);

AND2x6_ASAP7_75t_SL g1914 ( 
.A(n_1786),
.B(n_1150),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1757),
.B(n_1729),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1819),
.B(n_1665),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1758),
.B(n_1318),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1758),
.B(n_1324),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1812),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1785),
.B(n_1669),
.Y(n_1920)
);

INVxp67_ASAP7_75t_SL g1921 ( 
.A(n_1812),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1840),
.B(n_1502),
.Y(n_1922)
);

A2O1A1Ixp33_ASAP7_75t_SL g1923 ( 
.A1(n_1848),
.A2(n_1585),
.B(n_1532),
.C(n_1338),
.Y(n_1923)
);

NOR3xp33_ASAP7_75t_L g1924 ( 
.A(n_1846),
.B(n_1444),
.C(n_1307),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1854),
.A2(n_1691),
.B(n_1679),
.C(n_1647),
.Y(n_1925)
);

OAI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1910),
.A2(n_1838),
.B(n_1897),
.Y(n_1926)
);

A2O1A1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1868),
.A2(n_1638),
.B(n_1497),
.C(n_1422),
.Y(n_1927)
);

O2A1O1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1851),
.A2(n_1456),
.B(n_1154),
.C(n_1158),
.Y(n_1928)
);

O2A1O1Ixp33_ASAP7_75t_SL g1929 ( 
.A1(n_1889),
.A2(n_1890),
.B(n_1893),
.C(n_1905),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1900),
.B(n_1330),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1870),
.B(n_1339),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1859),
.A2(n_1678),
.B(n_1673),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1835),
.B(n_1815),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1860),
.A2(n_1738),
.B(n_1606),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1879),
.A2(n_1347),
.B1(n_1415),
.B2(n_1342),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1872),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1850),
.A2(n_1882),
.B(n_1874),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1841),
.A2(n_1606),
.B(n_1421),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1899),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1863),
.A2(n_1430),
.B1(n_1432),
.B2(n_1420),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1858),
.A2(n_1159),
.B(n_1160),
.C(n_1151),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1855),
.A2(n_1486),
.B(n_1452),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1836),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1839),
.A2(n_1487),
.B1(n_1499),
.B2(n_1494),
.Y(n_1944)
);

O2A1O1Ixp33_ASAP7_75t_L g1945 ( 
.A1(n_1869),
.A2(n_1166),
.B(n_1167),
.C(n_1164),
.Y(n_1945)
);

OAI21xp33_ASAP7_75t_L g1946 ( 
.A1(n_1896),
.A2(n_1538),
.B(n_1507),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1862),
.Y(n_1947)
);

NOR2xp67_ASAP7_75t_L g1948 ( 
.A(n_1865),
.B(n_1674),
.Y(n_1948)
);

NAND2x1p5_ASAP7_75t_L g1949 ( 
.A(n_1849),
.B(n_1729),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1873),
.A2(n_1523),
.B1(n_1547),
.B2(n_1545),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1871),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1881),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1856),
.A2(n_1602),
.B(n_1688),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1911),
.B(n_1682),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1843),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1842),
.B(n_1378),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1861),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1866),
.B(n_1424),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1911),
.B(n_1686),
.Y(n_1959)
);

NOR3xp33_ASAP7_75t_L g1960 ( 
.A(n_1864),
.B(n_1296),
.C(n_1188),
.Y(n_1960)
);

O2A1O1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1907),
.A2(n_1171),
.B(n_1175),
.C(n_1169),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1849),
.B(n_1424),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_R g1963 ( 
.A(n_1837),
.B(n_1275),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1857),
.A2(n_1845),
.B(n_1844),
.Y(n_1964)
);

OAI21xp33_ASAP7_75t_L g1965 ( 
.A1(n_1894),
.A2(n_1574),
.B(n_1539),
.Y(n_1965)
);

NAND2x1_ASAP7_75t_L g1966 ( 
.A(n_1852),
.B(n_1689),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1837),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1895),
.A2(n_1442),
.B1(n_1533),
.B2(n_1428),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1834),
.A2(n_1568),
.B1(n_1161),
.B2(n_1168),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1861),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1853),
.A2(n_1728),
.B(n_1703),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1875),
.B(n_1424),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1917),
.A2(n_1187),
.B(n_1191),
.C(n_1186),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1876),
.A2(n_1737),
.B(n_1195),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1913),
.A2(n_1170),
.B1(n_1176),
.B2(n_1157),
.Y(n_1975)
);

O2A1O1Ixp5_ASAP7_75t_L g1976 ( 
.A1(n_1847),
.A2(n_1411),
.B(n_1457),
.C(n_1380),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1901),
.A2(n_1180),
.B1(n_1181),
.B2(n_1177),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1883),
.B(n_1424),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1884),
.B(n_1737),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1908),
.A2(n_1201),
.B1(n_1208),
.B2(n_1189),
.Y(n_1980)
);

O2A1O1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1918),
.A2(n_1196),
.B(n_1197),
.C(n_1192),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1916),
.A2(n_1212),
.B(n_1207),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1920),
.A2(n_1215),
.B(n_1213),
.Y(n_1983)
);

O2A1O1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1886),
.A2(n_1223),
.B(n_1224),
.C(n_1221),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1902),
.A2(n_1226),
.B(n_1225),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1904),
.Y(n_1986)
);

A2O1A1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1903),
.A2(n_1475),
.B(n_1488),
.C(n_1459),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1891),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1885),
.A2(n_1233),
.B(n_1232),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1867),
.B(n_1209),
.Y(n_1990)
);

OAI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1887),
.A2(n_1235),
.B(n_1234),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1888),
.A2(n_1239),
.B(n_1237),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1878),
.B(n_1705),
.Y(n_1993)
);

AOI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1898),
.A2(n_1241),
.B(n_1240),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1880),
.A2(n_1214),
.B1(n_1217),
.B2(n_1210),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1921),
.B(n_1220),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1912),
.B(n_1396),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1861),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1909),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1877),
.B(n_1222),
.Y(n_2000)
);

OAI22x1_ASAP7_75t_L g2001 ( 
.A1(n_1892),
.A2(n_1715),
.B1(n_1230),
.B2(n_1244),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1919),
.B(n_1229),
.Y(n_2002)
);

OAI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1906),
.A2(n_1315),
.B1(n_1343),
.B2(n_1284),
.Y(n_2003)
);

OAI21xp33_ASAP7_75t_L g2004 ( 
.A1(n_1915),
.A2(n_1246),
.B(n_1243),
.Y(n_2004)
);

AO21x1_ASAP7_75t_L g2005 ( 
.A1(n_1914),
.A2(n_1252),
.B(n_1251),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1840),
.B(n_1245),
.Y(n_2006)
);

AOI22x1_ASAP7_75t_L g2007 ( 
.A1(n_1873),
.A2(n_1261),
.B1(n_1262),
.B2(n_1250),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1840),
.B(n_1264),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1910),
.A2(n_1255),
.B(n_1253),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1840),
.A2(n_1259),
.B(n_1256),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1891),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1840),
.B(n_1270),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1910),
.A2(n_1268),
.B(n_1266),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1840),
.B(n_1271),
.Y(n_2014)
);

AO21x1_ASAP7_75t_L g2015 ( 
.A1(n_1846),
.A2(n_1272),
.B(n_1269),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1840),
.A2(n_1529),
.B(n_1543),
.C(n_1514),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1836),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1910),
.A2(n_1279),
.B(n_1278),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1840),
.B(n_1291),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1910),
.A2(n_1281),
.B(n_1280),
.Y(n_2020)
);

AOI21xp33_ASAP7_75t_L g2021 ( 
.A1(n_1840),
.A2(n_1304),
.B(n_1302),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1861),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1840),
.B(n_1305),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1872),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1840),
.B(n_1312),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1910),
.A2(n_1288),
.B(n_1285),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1910),
.A2(n_1292),
.B(n_1290),
.Y(n_2027)
);

AOI33xp33_ASAP7_75t_L g2028 ( 
.A1(n_1880),
.A2(n_1482),
.A3(n_1371),
.B1(n_1506),
.B2(n_1425),
.B3(n_1303),
.Y(n_2028)
);

NOR2x1p5_ASAP7_75t_L g2029 ( 
.A(n_1840),
.B(n_1314),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1910),
.A2(n_1294),
.B(n_1293),
.Y(n_2030)
);

OAI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1840),
.A2(n_1298),
.B(n_1297),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1910),
.A2(n_1308),
.B(n_1306),
.Y(n_2032)
);

A2O1A1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1840),
.A2(n_1605),
.B(n_1588),
.C(n_1320),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1840),
.B(n_1316),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1840),
.B(n_1325),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1910),
.A2(n_1321),
.B(n_1310),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1836),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1910),
.A2(n_1329),
.B(n_1328),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_SL g2039 ( 
.A(n_1878),
.B(n_1379),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1840),
.B(n_1326),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1840),
.A2(n_1335),
.B(n_1331),
.Y(n_2041)
);

INVx4_ASAP7_75t_L g2042 ( 
.A(n_1849),
.Y(n_2042)
);

A2O1A1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1840),
.A2(n_1350),
.B(n_1351),
.C(n_1346),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1872),
.Y(n_2044)
);

NOR2xp67_ASAP7_75t_L g2045 ( 
.A(n_1865),
.B(n_945),
.Y(n_2045)
);

A2O1A1Ixp33_ASAP7_75t_SL g2046 ( 
.A1(n_1840),
.A2(n_1356),
.B(n_1361),
.C(n_1353),
.Y(n_2046)
);

AOI21x1_ASAP7_75t_L g2047 ( 
.A1(n_1910),
.A2(n_1369),
.B(n_1364),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1840),
.B(n_1333),
.Y(n_2048)
);

INVx3_ASAP7_75t_L g2049 ( 
.A(n_1861),
.Y(n_2049)
);

INVx4_ASAP7_75t_L g2050 ( 
.A(n_1849),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1910),
.A2(n_1373),
.B(n_1372),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1836),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1861),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_L g2054 ( 
.A(n_1840),
.B(n_1334),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1836),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1836),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1870),
.B(n_1396),
.Y(n_2057)
);

INVx3_ASAP7_75t_L g2058 ( 
.A(n_1861),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1840),
.A2(n_1381),
.B1(n_1383),
.B2(n_1375),
.Y(n_2059)
);

O2A1O1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_1840),
.A2(n_1391),
.B(n_1392),
.C(n_1388),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1840),
.A2(n_1397),
.B1(n_1404),
.B2(n_1394),
.Y(n_2061)
);

AO32x2_ASAP7_75t_L g2062 ( 
.A1(n_1995),
.A2(n_26),
.A3(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_2062)
);

OAI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1926),
.A2(n_1414),
.B(n_1408),
.Y(n_2063)
);

OA22x2_ASAP7_75t_L g2064 ( 
.A1(n_2001),
.A2(n_1340),
.B1(n_1345),
.B2(n_1336),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2048),
.B(n_1354),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_1937),
.A2(n_1427),
.B(n_1416),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1967),
.B(n_1439),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_SL g2068 ( 
.A1(n_1925),
.A2(n_949),
.B(n_947),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1932),
.A2(n_1964),
.B(n_2047),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_SL g2070 ( 
.A1(n_1927),
.A2(n_951),
.B(n_950),
.Y(n_2070)
);

NAND3xp33_ASAP7_75t_SL g2071 ( 
.A(n_2010),
.B(n_2041),
.C(n_2031),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1929),
.A2(n_1451),
.B(n_1447),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1930),
.A2(n_1460),
.B(n_1454),
.Y(n_2073)
);

AO31x2_ASAP7_75t_L g2074 ( 
.A1(n_2015),
.A2(n_1467),
.A3(n_1468),
.B(n_1466),
.Y(n_2074)
);

BUFx5_ASAP7_75t_L g2075 ( 
.A(n_1955),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1931),
.A2(n_1490),
.B(n_1485),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1922),
.B(n_1355),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1934),
.A2(n_1492),
.B(n_1491),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_2044),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1954),
.B(n_1496),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2057),
.B(n_1409),
.Y(n_2081)
);

AO21x2_ASAP7_75t_L g2082 ( 
.A1(n_1958),
.A2(n_1501),
.B(n_1498),
.Y(n_2082)
);

OAI21x1_ASAP7_75t_L g2083 ( 
.A1(n_2009),
.A2(n_1511),
.B(n_1504),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1986),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_2013),
.A2(n_1515),
.B(n_1513),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2006),
.B(n_2008),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_L g2087 ( 
.A1(n_2018),
.A2(n_1524),
.B(n_1520),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1959),
.B(n_1525),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1933),
.B(n_2012),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_2014),
.B(n_1419),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2019),
.B(n_1358),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1996),
.A2(n_1541),
.B(n_1535),
.Y(n_2092)
);

A2O1A1Ixp33_ASAP7_75t_L g2093 ( 
.A1(n_2021),
.A2(n_1548),
.B(n_1551),
.C(n_1544),
.Y(n_2093)
);

OAI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2023),
.A2(n_1558),
.B(n_1557),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_2020),
.A2(n_1561),
.B(n_1559),
.Y(n_2095)
);

O2A1O1Ixp5_ASAP7_75t_L g2096 ( 
.A1(n_1962),
.A2(n_1573),
.B(n_1584),
.C(n_1565),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2000),
.A2(n_2054),
.B1(n_2029),
.B2(n_2035),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2034),
.B(n_1366),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_2026),
.A2(n_1593),
.B(n_1589),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2040),
.B(n_1370),
.Y(n_2100)
);

NOR2x1_ASAP7_75t_SL g2101 ( 
.A(n_1957),
.B(n_1597),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1943),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1988),
.Y(n_2103)
);

AO31x2_ASAP7_75t_L g2104 ( 
.A1(n_2016),
.A2(n_1600),
.A3(n_1608),
.B(n_1599),
.Y(n_2104)
);

AO22x2_ASAP7_75t_L g2105 ( 
.A1(n_1924),
.A2(n_1611),
.B1(n_1613),
.B2(n_1609),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_2027),
.A2(n_1617),
.B(n_953),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_L g2107 ( 
.A1(n_1928),
.A2(n_1377),
.B(n_1382),
.C(n_1376),
.Y(n_2107)
);

OAI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2025),
.A2(n_1616),
.B(n_1615),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_2030),
.A2(n_956),
.B(n_952),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1951),
.A2(n_1389),
.B(n_1387),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1952),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1947),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1970),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2017),
.A2(n_1399),
.B(n_1395),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2055),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2037),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2052),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1939),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2056),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1972),
.A2(n_1402),
.B(n_1400),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_2024),
.Y(n_2121)
);

AOI31xp67_ASAP7_75t_L g2122 ( 
.A1(n_1978),
.A2(n_961),
.A3(n_962),
.B(n_958),
.Y(n_2122)
);

INVx2_ASAP7_75t_SL g2123 ( 
.A(n_1936),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1999),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_2002),
.A2(n_1407),
.B(n_1406),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_2032),
.A2(n_2038),
.B(n_2036),
.Y(n_2126)
);

BUFx10_ASAP7_75t_L g2127 ( 
.A(n_1993),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2003),
.B(n_1434),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1979),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1966),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1957),
.Y(n_2131)
);

AO31x2_ASAP7_75t_L g2132 ( 
.A1(n_2033),
.A2(n_29),
.A3(n_26),
.B(n_28),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_2051),
.A2(n_964),
.B(n_963),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_2011),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_1923),
.A2(n_1417),
.B(n_1412),
.Y(n_2135)
);

OAI21xp33_ASAP7_75t_L g2136 ( 
.A1(n_2059),
.A2(n_1435),
.B(n_1426),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1935),
.B(n_1437),
.Y(n_2137)
);

AO22x2_ASAP7_75t_L g2138 ( 
.A1(n_1968),
.A2(n_1590),
.B1(n_1489),
.B2(n_1556),
.Y(n_2138)
);

OAI21x1_ASAP7_75t_L g2139 ( 
.A1(n_1976),
.A2(n_966),
.B(n_965),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1956),
.B(n_1438),
.Y(n_2140)
);

AO31x2_ASAP7_75t_L g2141 ( 
.A1(n_2043),
.A2(n_30),
.A3(n_28),
.B(n_29),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1957),
.Y(n_2142)
);

NOR2xp67_ASAP7_75t_L g2143 ( 
.A(n_2042),
.B(n_971),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2061),
.B(n_1440),
.Y(n_2144)
);

AOI21x1_ASAP7_75t_L g2145 ( 
.A1(n_1942),
.A2(n_973),
.B(n_972),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_2022),
.A2(n_2058),
.B(n_2049),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1946),
.B(n_1441),
.Y(n_2147)
);

BUFx3_ASAP7_75t_L g2148 ( 
.A(n_1998),
.Y(n_2148)
);

AO31x2_ASAP7_75t_L g2149 ( 
.A1(n_1987),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_1969),
.B(n_1582),
.Y(n_2150)
);

AO31x2_ASAP7_75t_L g2151 ( 
.A1(n_1985),
.A2(n_34),
.A3(n_31),
.B(n_33),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_L g2152 ( 
.A1(n_1971),
.A2(n_975),
.B(n_974),
.Y(n_2152)
);

BUFx2_ASAP7_75t_L g2153 ( 
.A(n_1998),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1998),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2053),
.Y(n_2155)
);

AOI211x1_ASAP7_75t_L g2156 ( 
.A1(n_1982),
.A2(n_1476),
.B(n_1483),
.C(n_1409),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_1940),
.A2(n_1607),
.B(n_1603),
.Y(n_2157)
);

AO31x2_ASAP7_75t_L g2158 ( 
.A1(n_1938),
.A2(n_1983),
.A3(n_1977),
.B(n_1975),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_2050),
.B(n_1521),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1950),
.B(n_1446),
.Y(n_2160)
);

OAI21x1_ASAP7_75t_L g2161 ( 
.A1(n_1949),
.A2(n_980),
.B(n_978),
.Y(n_2161)
);

OAI21x1_ASAP7_75t_L g2162 ( 
.A1(n_1989),
.A2(n_983),
.B(n_981),
.Y(n_2162)
);

OAI21x1_ASAP7_75t_L g2163 ( 
.A1(n_1992),
.A2(n_987),
.B(n_984),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_2045),
.A2(n_990),
.B(n_989),
.Y(n_2164)
);

BUFx3_ASAP7_75t_L g2165 ( 
.A(n_2053),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1953),
.A2(n_1453),
.B(n_1449),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2053),
.Y(n_2167)
);

AOI221x1_ASAP7_75t_L g2168 ( 
.A1(n_1960),
.A2(n_995),
.B1(n_996),
.B2(n_994),
.C(n_992),
.Y(n_2168)
);

INVx1_ASAP7_75t_SL g2169 ( 
.A(n_1997),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_1948),
.A2(n_1461),
.B(n_1455),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1991),
.B(n_1462),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1990),
.B(n_1564),
.Y(n_2172)
);

OAI21x1_ASAP7_75t_L g2173 ( 
.A1(n_1994),
.A2(n_999),
.B(n_997),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1965),
.B(n_1464),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1945),
.A2(n_1471),
.B(n_1470),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_1973),
.A2(n_1473),
.B(n_1472),
.Y(n_2176)
);

BUFx4_ASAP7_75t_SL g2177 ( 
.A(n_1963),
.Y(n_2177)
);

AO21x2_ASAP7_75t_L g2178 ( 
.A1(n_2046),
.A2(n_1944),
.B(n_2004),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2007),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2039),
.B(n_1476),
.Y(n_2180)
);

INVx3_ASAP7_75t_L g2181 ( 
.A(n_1984),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_1981),
.A2(n_1479),
.B(n_1478),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2028),
.B(n_1480),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1941),
.B(n_2060),
.Y(n_2184)
);

OAI21x1_ASAP7_75t_L g2185 ( 
.A1(n_1974),
.A2(n_1003),
.B(n_1002),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1980),
.B(n_1484),
.Y(n_2186)
);

OAI21x1_ASAP7_75t_L g2187 ( 
.A1(n_1961),
.A2(n_1006),
.B(n_1005),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2005),
.B(n_1495),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2048),
.A2(n_1612),
.B1(n_1614),
.B2(n_1580),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2048),
.B(n_1483),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1988),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1986),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2048),
.A2(n_1503),
.B1(n_1505),
.B2(n_1500),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2048),
.B(n_1508),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_1937),
.A2(n_1008),
.B(n_1007),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2048),
.B(n_1510),
.Y(n_2196)
);

AO21x2_ASAP7_75t_L g2197 ( 
.A1(n_1926),
.A2(n_1011),
.B(n_1010),
.Y(n_2197)
);

CKINVDCx8_ASAP7_75t_R g2198 ( 
.A(n_1988),
.Y(n_2198)
);

INVx4_ASAP7_75t_SL g2199 ( 
.A(n_1967),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_SL g2200 ( 
.A(n_2010),
.B(n_1512),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_1936),
.B(n_1517),
.Y(n_2201)
);

BUFx3_ASAP7_75t_L g2202 ( 
.A(n_1967),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_2044),
.Y(n_2203)
);

AOI221x1_ASAP7_75t_L g2204 ( 
.A1(n_1927),
.A2(n_1018),
.B1(n_1022),
.B2(n_1015),
.C(n_1013),
.Y(n_2204)
);

AOI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_1926),
.A2(n_1526),
.B(n_1518),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2048),
.B(n_1528),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2048),
.B(n_1530),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1986),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_1926),
.A2(n_1540),
.B(n_1536),
.Y(n_2209)
);

AOI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_1926),
.A2(n_1549),
.B(n_1546),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_1926),
.A2(n_1562),
.B(n_1552),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2024),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2048),
.B(n_1570),
.Y(n_2213)
);

AOI21x1_ASAP7_75t_SL g2214 ( 
.A1(n_2000),
.A2(n_1572),
.B(n_1571),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_1926),
.A2(n_1576),
.B(n_1575),
.Y(n_2215)
);

INVx4_ASAP7_75t_L g2216 ( 
.A(n_1967),
.Y(n_2216)
);

OAI21x1_ASAP7_75t_L g2217 ( 
.A1(n_1937),
.A2(n_1029),
.B(n_1028),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2048),
.A2(n_1581),
.B1(n_1587),
.B2(n_1577),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1957),
.Y(n_2219)
);

OAI21x1_ASAP7_75t_L g2220 ( 
.A1(n_1937),
.A2(n_1031),
.B(n_1030),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2048),
.A2(n_1592),
.B1(n_1595),
.B2(n_1591),
.Y(n_2221)
);

AO31x2_ASAP7_75t_L g2222 ( 
.A1(n_1925),
.A2(n_37),
.A3(n_35),
.B(n_36),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_1936),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_1937),
.A2(n_1034),
.B(n_1032),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_SL g2225 ( 
.A1(n_2048),
.A2(n_1598),
.B(n_1596),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2048),
.B(n_1610),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_2044),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_1926),
.A2(n_1036),
.B(n_1035),
.Y(n_2228)
);

A2O1A1Ixp33_ASAP7_75t_L g2229 ( 
.A1(n_2048),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_2229)
);

OAI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_1926),
.A2(n_1039),
.B(n_1038),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1986),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1986),
.Y(n_2232)
);

NAND2x1p5_ASAP7_75t_L g2233 ( 
.A(n_2042),
.B(n_1040),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1937),
.A2(n_1043),
.B(n_1041),
.Y(n_2234)
);

AOI21xp5_ASAP7_75t_SL g2235 ( 
.A1(n_1925),
.A2(n_1045),
.B(n_1044),
.Y(n_2235)
);

OAI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_1926),
.A2(n_1050),
.B(n_1046),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2048),
.B(n_38),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_1967),
.B(n_1051),
.Y(n_2238)
);

OA21x2_ASAP7_75t_L g2239 ( 
.A1(n_1932),
.A2(n_1053),
.B(n_1052),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2111),
.Y(n_2240)
);

OAI21x1_ASAP7_75t_L g2241 ( 
.A1(n_2066),
.A2(n_2069),
.B(n_2078),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_SL g2242 ( 
.A1(n_2230),
.A2(n_1055),
.B(n_1054),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_2079),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2089),
.B(n_39),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2084),
.Y(n_2245)
);

OAI21x1_ASAP7_75t_L g2246 ( 
.A1(n_2146),
.A2(n_1057),
.B(n_1056),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2202),
.B(n_1058),
.Y(n_2247)
);

OAI21xp33_ASAP7_75t_SL g2248 ( 
.A1(n_2086),
.A2(n_39),
.B(n_40),
.Y(n_2248)
);

OA21x2_ASAP7_75t_L g2249 ( 
.A1(n_2236),
.A2(n_1064),
.B(n_1059),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_2199),
.B(n_1066),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2090),
.B(n_40),
.Y(n_2251)
);

AO21x2_ASAP7_75t_L g2252 ( 
.A1(n_2071),
.A2(n_1069),
.B(n_1067),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2192),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2115),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2203),
.Y(n_2255)
);

OR2x6_ASAP7_75t_L g2256 ( 
.A(n_2123),
.B(n_41),
.Y(n_2256)
);

OAI21x1_ASAP7_75t_L g2257 ( 
.A1(n_2126),
.A2(n_1071),
.B(n_1070),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2070),
.A2(n_1074),
.B(n_1072),
.Y(n_2258)
);

OAI21x1_ASAP7_75t_L g2259 ( 
.A1(n_2195),
.A2(n_2234),
.B(n_2220),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_2219),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2119),
.Y(n_2261)
);

OAI21x1_ASAP7_75t_L g2262 ( 
.A1(n_2217),
.A2(n_1076),
.B(n_1075),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2227),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2199),
.B(n_1077),
.Y(n_2264)
);

OA21x2_ASAP7_75t_L g2265 ( 
.A1(n_2204),
.A2(n_1079),
.B(n_1078),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2208),
.Y(n_2266)
);

OAI21x1_ASAP7_75t_L g2267 ( 
.A1(n_2224),
.A2(n_1082),
.B(n_1080),
.Y(n_2267)
);

HB1xp67_ASAP7_75t_L g2268 ( 
.A(n_2212),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_2223),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2065),
.B(n_2194),
.Y(n_2270)
);

AO21x2_ASAP7_75t_L g2271 ( 
.A1(n_2063),
.A2(n_1084),
.B(n_1083),
.Y(n_2271)
);

OAI21x1_ASAP7_75t_L g2272 ( 
.A1(n_2106),
.A2(n_2139),
.B(n_2133),
.Y(n_2272)
);

OAI21x1_ASAP7_75t_L g2273 ( 
.A1(n_2109),
.A2(n_1086),
.B(n_1085),
.Y(n_2273)
);

BUFx2_ASAP7_75t_L g2274 ( 
.A(n_2103),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2216),
.B(n_2121),
.Y(n_2275)
);

OR2x6_ASAP7_75t_L g2276 ( 
.A(n_2238),
.B(n_41),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2152),
.A2(n_1089),
.B(n_1088),
.Y(n_2277)
);

AO31x2_ASAP7_75t_L g2278 ( 
.A1(n_2072),
.A2(n_1130),
.A3(n_1131),
.B(n_1129),
.Y(n_2278)
);

AO21x2_ASAP7_75t_L g2279 ( 
.A1(n_2228),
.A2(n_1092),
.B(n_1091),
.Y(n_2279)
);

AOI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2068),
.A2(n_1094),
.B(n_1093),
.Y(n_2280)
);

OAI21x1_ASAP7_75t_SL g2281 ( 
.A1(n_2101),
.A2(n_1099),
.B(n_1096),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2134),
.B(n_42),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2196),
.B(n_43),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2219),
.Y(n_2284)
);

NOR2xp67_ASAP7_75t_L g2285 ( 
.A(n_2191),
.B(n_2118),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2231),
.Y(n_2286)
);

OA21x2_ASAP7_75t_L g2287 ( 
.A1(n_2179),
.A2(n_1101),
.B(n_1100),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2153),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_2198),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2097),
.B(n_1103),
.Y(n_2290)
);

OAI21x1_ASAP7_75t_L g2291 ( 
.A1(n_2162),
.A2(n_1105),
.B(n_1104),
.Y(n_2291)
);

OA21x2_ASAP7_75t_L g2292 ( 
.A1(n_2083),
.A2(n_1108),
.B(n_1107),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2232),
.Y(n_2293)
);

NAND2x1p5_ASAP7_75t_L g2294 ( 
.A(n_2148),
.B(n_1109),
.Y(n_2294)
);

OAI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2237),
.A2(n_1111),
.B(n_1110),
.Y(n_2295)
);

BUFx3_ASAP7_75t_L g2296 ( 
.A(n_2165),
.Y(n_2296)
);

A2O1A1Ixp33_ASAP7_75t_L g2297 ( 
.A1(n_2094),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2102),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2112),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_2067),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2206),
.B(n_44),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2207),
.B(n_2213),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2081),
.B(n_46),
.Y(n_2303)
);

OR2x2_ASAP7_75t_L g2304 ( 
.A(n_2201),
.B(n_2169),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2235),
.A2(n_1117),
.B(n_1112),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2226),
.B(n_46),
.Y(n_2306)
);

AND2x6_ASAP7_75t_L g2307 ( 
.A(n_2181),
.B(n_1119),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2116),
.Y(n_2308)
);

OA21x2_ASAP7_75t_L g2309 ( 
.A1(n_2085),
.A2(n_1121),
.B(n_1120),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2117),
.Y(n_2310)
);

OAI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2205),
.A2(n_1123),
.B(n_1122),
.Y(n_2311)
);

OAI21x1_ASAP7_75t_L g2312 ( 
.A1(n_2163),
.A2(n_1125),
.B(n_1124),
.Y(n_2312)
);

AO21x2_ASAP7_75t_L g2313 ( 
.A1(n_2197),
.A2(n_1127),
.B(n_1126),
.Y(n_2313)
);

OAI21x1_ASAP7_75t_L g2314 ( 
.A1(n_2173),
.A2(n_1135),
.B(n_1128),
.Y(n_2314)
);

OA21x2_ASAP7_75t_L g2315 ( 
.A1(n_2087),
.A2(n_1140),
.B(n_1139),
.Y(n_2315)
);

INVx4_ASAP7_75t_L g2316 ( 
.A(n_2113),
.Y(n_2316)
);

BUFx2_ASAP7_75t_L g2317 ( 
.A(n_2142),
.Y(n_2317)
);

AO222x2_ASAP7_75t_L g2318 ( 
.A1(n_2172),
.A2(n_49),
.B1(n_51),
.B2(n_47),
.C1(n_48),
.C2(n_50),
.Y(n_2318)
);

OAI21x1_ASAP7_75t_L g2319 ( 
.A1(n_2185),
.A2(n_1143),
.B(n_1142),
.Y(n_2319)
);

AO21x2_ASAP7_75t_L g2320 ( 
.A1(n_2209),
.A2(n_1145),
.B(n_1144),
.Y(n_2320)
);

OAI21x1_ASAP7_75t_L g2321 ( 
.A1(n_2214),
.A2(n_1147),
.B(n_1146),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2167),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2124),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_2080),
.Y(n_2324)
);

OAI21x1_ASAP7_75t_L g2325 ( 
.A1(n_2161),
.A2(n_1148),
.B(n_47),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_2088),
.B(n_48),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2131),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2075),
.Y(n_2328)
);

OA21x2_ASAP7_75t_L g2329 ( 
.A1(n_2095),
.A2(n_49),
.B(n_50),
.Y(n_2329)
);

BUFx2_ASAP7_75t_SL g2330 ( 
.A(n_2159),
.Y(n_2330)
);

BUFx2_ASAP7_75t_R g2331 ( 
.A(n_2178),
.Y(n_2331)
);

INVx1_ASAP7_75t_SL g2332 ( 
.A(n_2177),
.Y(n_2332)
);

OAI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_2210),
.A2(n_51),
.B(n_52),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_2099),
.A2(n_53),
.B(n_54),
.Y(n_2334)
);

OAI21x1_ASAP7_75t_L g2335 ( 
.A1(n_2145),
.A2(n_53),
.B(n_54),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2129),
.B(n_55),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2190),
.B(n_55),
.Y(n_2337)
);

OA21x2_ASAP7_75t_L g2338 ( 
.A1(n_2187),
.A2(n_56),
.B(n_57),
.Y(n_2338)
);

BUFx3_ASAP7_75t_L g2339 ( 
.A(n_2127),
.Y(n_2339)
);

OAI21x1_ASAP7_75t_L g2340 ( 
.A1(n_2130),
.A2(n_57),
.B(n_58),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2091),
.B(n_58),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2180),
.B(n_59),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2189),
.B(n_914),
.Y(n_2343)
);

AO31x2_ASAP7_75t_L g2344 ( 
.A1(n_2168),
.A2(n_62),
.A3(n_59),
.B(n_61),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2154),
.Y(n_2345)
);

OAI21x1_ASAP7_75t_L g2346 ( 
.A1(n_2239),
.A2(n_62),
.B(n_63),
.Y(n_2346)
);

AOI21xp5_ASAP7_75t_L g2347 ( 
.A1(n_2098),
.A2(n_63),
.B(n_64),
.Y(n_2347)
);

NOR2xp67_ASAP7_75t_L g2348 ( 
.A(n_2140),
.B(n_65),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2155),
.Y(n_2349)
);

OAI21x1_ASAP7_75t_L g2350 ( 
.A1(n_2233),
.A2(n_2076),
.B(n_2096),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2100),
.A2(n_65),
.B(n_66),
.Y(n_2351)
);

A2O1A1Ixp33_ASAP7_75t_L g2352 ( 
.A1(n_2157),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_2062),
.Y(n_2353)
);

BUFx2_ASAP7_75t_L g2354 ( 
.A(n_2064),
.Y(n_2354)
);

OAI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2211),
.A2(n_67),
.B(n_68),
.Y(n_2355)
);

AOI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2215),
.A2(n_69),
.B(n_70),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2104),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2104),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2077),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2128),
.B(n_909),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2143),
.A2(n_71),
.B(n_72),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2075),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2075),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2075),
.Y(n_2364)
);

BUFx12f_ASAP7_75t_L g2365 ( 
.A(n_2150),
.Y(n_2365)
);

INVx4_ASAP7_75t_SL g2366 ( 
.A(n_2151),
.Y(n_2366)
);

CKINVDCx8_ASAP7_75t_R g2367 ( 
.A(n_2138),
.Y(n_2367)
);

OAI21x1_ASAP7_75t_L g2368 ( 
.A1(n_2073),
.A2(n_72),
.B(n_73),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_2186),
.B(n_73),
.Y(n_2369)
);

OAI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2184),
.A2(n_74),
.B(n_75),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_2147),
.A2(n_74),
.B(n_75),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_SL g2372 ( 
.A1(n_2164),
.A2(n_76),
.B(n_77),
.Y(n_2372)
);

INVxp67_ASAP7_75t_SL g2373 ( 
.A(n_2188),
.Y(n_2373)
);

CKINVDCx6p67_ASAP7_75t_R g2374 ( 
.A(n_2183),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2225),
.B(n_77),
.Y(n_2375)
);

NAND2x1p5_ASAP7_75t_L g2376 ( 
.A(n_2200),
.B(n_78),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2074),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2171),
.B(n_78),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2137),
.A2(n_79),
.B(n_80),
.Y(n_2379)
);

OR2x6_ASAP7_75t_L g2380 ( 
.A(n_2330),
.B(n_2156),
.Y(n_2380)
);

AO21x2_ASAP7_75t_L g2381 ( 
.A1(n_2241),
.A2(n_2082),
.B(n_2092),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2245),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2270),
.B(n_2074),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2253),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2275),
.Y(n_2385)
);

OAI21x1_ASAP7_75t_L g2386 ( 
.A1(n_2259),
.A2(n_2114),
.B(n_2110),
.Y(n_2386)
);

AO21x2_ASAP7_75t_L g2387 ( 
.A1(n_2272),
.A2(n_2093),
.B(n_2107),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_2243),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2293),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2304),
.B(n_2144),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2251),
.B(n_2105),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2255),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2268),
.Y(n_2393)
);

AOI21x1_ASAP7_75t_L g2394 ( 
.A1(n_2290),
.A2(n_2120),
.B(n_2174),
.Y(n_2394)
);

INVx3_ASAP7_75t_L g2395 ( 
.A(n_2296),
.Y(n_2395)
);

OR2x2_ASAP7_75t_L g2396 ( 
.A(n_2244),
.B(n_2160),
.Y(n_2396)
);

AO21x2_ASAP7_75t_L g2397 ( 
.A1(n_2377),
.A2(n_2229),
.B(n_2125),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2266),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2298),
.Y(n_2399)
);

OAI21x1_ASAP7_75t_L g2400 ( 
.A1(n_2257),
.A2(n_2135),
.B(n_2166),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2286),
.Y(n_2401)
);

BUFx2_ASAP7_75t_L g2402 ( 
.A(n_2269),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2308),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2299),
.Y(n_2404)
);

AOI21xp33_ASAP7_75t_SL g2405 ( 
.A1(n_2343),
.A2(n_2221),
.B(n_2193),
.Y(n_2405)
);

HB1xp67_ASAP7_75t_L g2406 ( 
.A(n_2263),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2360),
.B(n_2108),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2310),
.Y(n_2408)
);

INVx5_ASAP7_75t_L g2409 ( 
.A(n_2260),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2323),
.Y(n_2410)
);

OR2x6_ASAP7_75t_L g2411 ( 
.A(n_2285),
.B(n_2175),
.Y(n_2411)
);

INVx4_ASAP7_75t_L g2412 ( 
.A(n_2260),
.Y(n_2412)
);

BUFx2_ASAP7_75t_L g2413 ( 
.A(n_2288),
.Y(n_2413)
);

OAI21x1_ASAP7_75t_L g2414 ( 
.A1(n_2319),
.A2(n_2170),
.B(n_2176),
.Y(n_2414)
);

AO21x2_ASAP7_75t_L g2415 ( 
.A1(n_2357),
.A2(n_2182),
.B(n_2122),
.Y(n_2415)
);

INVx2_ASAP7_75t_SL g2416 ( 
.A(n_2300),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2261),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2240),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2324),
.B(n_2158),
.Y(n_2419)
);

BUFx6f_ASAP7_75t_L g2420 ( 
.A(n_2284),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2254),
.Y(n_2421)
);

BUFx3_ASAP7_75t_L g2422 ( 
.A(n_2274),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2317),
.Y(n_2423)
);

OAI21x1_ASAP7_75t_L g2424 ( 
.A1(n_2246),
.A2(n_2218),
.B(n_2222),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2289),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2302),
.B(n_2136),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_2300),
.Y(n_2427)
);

INVxp33_ASAP7_75t_L g2428 ( 
.A(n_2282),
.Y(n_2428)
);

OA21x2_ASAP7_75t_L g2429 ( 
.A1(n_2346),
.A2(n_2222),
.B(n_2149),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2327),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_2322),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2284),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2345),
.Y(n_2433)
);

INVx3_ASAP7_75t_L g2434 ( 
.A(n_2316),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2336),
.Y(n_2435)
);

OAI21x1_ASAP7_75t_L g2436 ( 
.A1(n_2262),
.A2(n_2158),
.B(n_2149),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2349),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2354),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2358),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2328),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2340),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2364),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2333),
.A2(n_2062),
.B(n_2132),
.Y(n_2443)
);

INVxp67_ASAP7_75t_L g2444 ( 
.A(n_2342),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2362),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2378),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2303),
.B(n_2141),
.Y(n_2447)
);

BUFx2_ASAP7_75t_L g2448 ( 
.A(n_2339),
.Y(n_2448)
);

AOI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2363),
.A2(n_2132),
.B(n_2141),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2355),
.Y(n_2450)
);

OR2x6_ASAP7_75t_L g2451 ( 
.A(n_2276),
.B(n_2151),
.Y(n_2451)
);

INVxp67_ASAP7_75t_SL g2452 ( 
.A(n_2373),
.Y(n_2452)
);

INVxp67_ASAP7_75t_SL g2453 ( 
.A(n_2341),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2369),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2366),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2368),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2370),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2356),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2247),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2325),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2332),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2283),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2287),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2301),
.Y(n_2464)
);

AOI22xp33_ASAP7_75t_L g2465 ( 
.A1(n_2375),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2350),
.Y(n_2466)
);

OA21x2_ASAP7_75t_L g2467 ( 
.A1(n_2335),
.A2(n_81),
.B(n_82),
.Y(n_2467)
);

HB1xp67_ASAP7_75t_L g2468 ( 
.A(n_2276),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2326),
.B(n_901),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2306),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2353),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2337),
.B(n_82),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_2365),
.Y(n_2473)
);

OA21x2_ASAP7_75t_L g2474 ( 
.A1(n_2291),
.A2(n_83),
.B(n_84),
.Y(n_2474)
);

HB1xp67_ASAP7_75t_L g2475 ( 
.A(n_2256),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2256),
.Y(n_2476)
);

NAND2x1p5_ASAP7_75t_L g2477 ( 
.A(n_2250),
.B(n_83),
.Y(n_2477)
);

BUFx6f_ASAP7_75t_L g2478 ( 
.A(n_2264),
.Y(n_2478)
);

BUFx2_ASAP7_75t_L g2479 ( 
.A(n_2374),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2353),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2348),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2352),
.Y(n_2482)
);

INVx3_ASAP7_75t_L g2483 ( 
.A(n_2294),
.Y(n_2483)
);

CKINVDCx11_ASAP7_75t_R g2484 ( 
.A(n_2367),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2376),
.Y(n_2485)
);

OA21x2_ASAP7_75t_L g2486 ( 
.A1(n_2312),
.A2(n_84),
.B(n_85),
.Y(n_2486)
);

HB1xp67_ASAP7_75t_L g2487 ( 
.A(n_2248),
.Y(n_2487)
);

AND2x4_ASAP7_75t_L g2488 ( 
.A(n_2307),
.B(n_85),
.Y(n_2488)
);

AOI21x1_ASAP7_75t_L g2489 ( 
.A1(n_2242),
.A2(n_86),
.B(n_87),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2359),
.B(n_906),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2307),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2307),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2334),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2278),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2297),
.B(n_86),
.Y(n_2495)
);

OR2x2_ASAP7_75t_L g2496 ( 
.A(n_2347),
.B(n_87),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2344),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2344),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2277),
.Y(n_2499)
);

NOR2x1_ASAP7_75t_SL g2500 ( 
.A(n_2279),
.B(n_90),
.Y(n_2500)
);

AO31x2_ASAP7_75t_L g2501 ( 
.A1(n_2280),
.A2(n_92),
.A3(n_90),
.B(n_91),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_2320),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2321),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2351),
.B(n_914),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2331),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2329),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2252),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2273),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2371),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_2281),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2379),
.B(n_93),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2258),
.B(n_93),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2314),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2295),
.B(n_94),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2278),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2338),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2361),
.Y(n_2517)
);

AO21x2_ASAP7_75t_L g2518 ( 
.A1(n_2311),
.A2(n_94),
.B(n_95),
.Y(n_2518)
);

OAI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2305),
.A2(n_95),
.B(n_96),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2267),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2313),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2271),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2265),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2249),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2292),
.Y(n_2525)
);

INVx3_ASAP7_75t_L g2526 ( 
.A(n_2309),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2372),
.B(n_96),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2315),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2318),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2270),
.B(n_97),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2270),
.B(n_97),
.Y(n_2531)
);

INVx2_ASAP7_75t_SL g2532 ( 
.A(n_2409),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2407),
.B(n_98),
.Y(n_2533)
);

INVx4_ASAP7_75t_L g2534 ( 
.A(n_2409),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2454),
.B(n_98),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_2402),
.Y(n_2536)
);

INVxp33_ASAP7_75t_SL g2537 ( 
.A(n_2461),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2530),
.B(n_99),
.Y(n_2538)
);

INVx4_ASAP7_75t_L g2539 ( 
.A(n_2420),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2382),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2398),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2384),
.Y(n_2542)
);

OAI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2529),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2401),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2389),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2399),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2404),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2388),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2392),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2396),
.B(n_100),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2408),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2530),
.B(n_102),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2403),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2531),
.B(n_102),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2531),
.B(n_103),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2422),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2410),
.Y(n_2557)
);

OAI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2405),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2430),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2417),
.Y(n_2560)
);

OA21x2_ASAP7_75t_L g2561 ( 
.A1(n_2436),
.A2(n_104),
.B(n_105),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2437),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2421),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2433),
.Y(n_2564)
);

BUFx2_ASAP7_75t_L g2565 ( 
.A(n_2471),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2439),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2462),
.B(n_106),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2418),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2480),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2440),
.Y(n_2570)
);

AO21x2_ASAP7_75t_L g2571 ( 
.A1(n_2522),
.A2(n_106),
.B(n_107),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2442),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2445),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2496),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2464),
.B(n_107),
.Y(n_2575)
);

OR2x2_ASAP7_75t_L g2576 ( 
.A(n_2390),
.B(n_108),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2470),
.B(n_2446),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2511),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2509),
.Y(n_2579)
);

INVx2_ASAP7_75t_SL g2580 ( 
.A(n_2420),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2391),
.B(n_109),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2453),
.B(n_110),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2490),
.B(n_111),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2413),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2487),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2517),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2431),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2469),
.B(n_111),
.Y(n_2588)
);

CKINVDCx20_ASAP7_75t_R g2589 ( 
.A(n_2484),
.Y(n_2589)
);

INVx1_ASAP7_75t_SL g2590 ( 
.A(n_2423),
.Y(n_2590)
);

AO31x2_ASAP7_75t_L g2591 ( 
.A1(n_2457),
.A2(n_114),
.A3(n_112),
.B(n_113),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2449),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2497),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2426),
.B(n_113),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2498),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2458),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2393),
.B(n_114),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2406),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2441),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2506),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2419),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2432),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2516),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2452),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2504),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2383),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2435),
.Y(n_2607)
);

INVx1_ASAP7_75t_SL g2608 ( 
.A(n_2425),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2383),
.Y(n_2609)
);

BUFx2_ASAP7_75t_L g2610 ( 
.A(n_2451),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2495),
.Y(n_2611)
);

INVx3_ASAP7_75t_L g2612 ( 
.A(n_2395),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2456),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2501),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2463),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2447),
.B(n_115),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2448),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2523),
.Y(n_2618)
);

AO31x2_ASAP7_75t_L g2619 ( 
.A1(n_2493),
.A2(n_117),
.A3(n_115),
.B(n_116),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2438),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2460),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2447),
.B(n_116),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2472),
.B(n_117),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2478),
.Y(n_2624)
);

HB1xp67_ASAP7_75t_L g2625 ( 
.A(n_2475),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_2476),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2429),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2501),
.Y(n_2628)
);

NOR2x1_ASAP7_75t_L g2629 ( 
.A(n_2434),
.B(n_2491),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2451),
.Y(n_2630)
);

OAI21xp33_ASAP7_75t_L g2631 ( 
.A1(n_2514),
.A2(n_118),
.B(n_120),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2455),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2482),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2397),
.Y(n_2634)
);

OR2x2_ASAP7_75t_L g2635 ( 
.A(n_2428),
.B(n_121),
.Y(n_2635)
);

INVxp33_ASAP7_75t_L g2636 ( 
.A(n_2468),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2485),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2479),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_2412),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2459),
.B(n_121),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2467),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2512),
.Y(n_2642)
);

AO21x2_ASAP7_75t_L g2643 ( 
.A1(n_2466),
.A2(n_122),
.B(n_123),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2505),
.B(n_123),
.Y(n_2644)
);

INVxp67_ASAP7_75t_SL g2645 ( 
.A(n_2385),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2527),
.B(n_124),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2481),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2444),
.B(n_124),
.Y(n_2648)
);

OR2x2_ASAP7_75t_L g2649 ( 
.A(n_2478),
.B(n_2483),
.Y(n_2649)
);

BUFx2_ASAP7_75t_L g2650 ( 
.A(n_2494),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2527),
.B(n_125),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2500),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2416),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2474),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2486),
.Y(n_2655)
);

INVxp67_ASAP7_75t_SL g2656 ( 
.A(n_2492),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2488),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2518),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2450),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2465),
.B(n_126),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2477),
.B(n_127),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2489),
.Y(n_2662)
);

HB1xp67_ASAP7_75t_L g2663 ( 
.A(n_2427),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2381),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2510),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2387),
.Y(n_2666)
);

HB1xp67_ASAP7_75t_L g2667 ( 
.A(n_2411),
.Y(n_2667)
);

OR2x2_ASAP7_75t_L g2668 ( 
.A(n_2380),
.B(n_128),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2380),
.B(n_129),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2411),
.Y(n_2670)
);

BUFx6f_ASAP7_75t_L g2671 ( 
.A(n_2473),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2519),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2549),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2616),
.B(n_2443),
.Y(n_2674)
);

AND2x6_ASAP7_75t_SL g2675 ( 
.A(n_2550),
.B(n_129),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2577),
.B(n_2524),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2574),
.B(n_2578),
.Y(n_2677)
);

OR2x2_ASAP7_75t_L g2678 ( 
.A(n_2605),
.B(n_2515),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2622),
.B(n_2415),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2646),
.B(n_2424),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2566),
.Y(n_2681)
);

AND2x4_ASAP7_75t_L g2682 ( 
.A(n_2556),
.B(n_2386),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2651),
.B(n_2538),
.Y(n_2683)
);

INVxp67_ASAP7_75t_L g2684 ( 
.A(n_2598),
.Y(n_2684)
);

HB1xp67_ASAP7_75t_L g2685 ( 
.A(n_2620),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2642),
.A2(n_2631),
.B1(n_2657),
.B2(n_2611),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2552),
.B(n_2394),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2554),
.B(n_2521),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2590),
.B(n_2594),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2555),
.B(n_2502),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2593),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2581),
.B(n_2414),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2582),
.B(n_2507),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2583),
.B(n_2503),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2533),
.B(n_2503),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2595),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2606),
.B(n_2525),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2562),
.B(n_130),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2541),
.B(n_130),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2544),
.B(n_131),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2553),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2560),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2536),
.B(n_2499),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_2672),
.A2(n_2508),
.B1(n_2513),
.B2(n_2520),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2600),
.Y(n_2705)
);

AND2x4_ASAP7_75t_L g2706 ( 
.A(n_2584),
.B(n_2400),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2579),
.Y(n_2707)
);

NAND2xp33_ASAP7_75t_R g2708 ( 
.A(n_2638),
.B(n_2526),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2563),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2537),
.B(n_132),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2540),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2609),
.B(n_2528),
.Y(n_2712)
);

CKINVDCx16_ASAP7_75t_R g2713 ( 
.A(n_2589),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2587),
.B(n_2585),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2570),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2640),
.B(n_134),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2647),
.B(n_134),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2542),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2576),
.B(n_135),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2604),
.B(n_2623),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2601),
.B(n_136),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2572),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2548),
.B(n_136),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2629),
.B(n_137),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2660),
.B(n_138),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2567),
.B(n_139),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2534),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2545),
.Y(n_2728)
);

HB1xp67_ASAP7_75t_L g2729 ( 
.A(n_2565),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2644),
.B(n_139),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2575),
.B(n_140),
.Y(n_2731)
);

INVx2_ASAP7_75t_SL g2732 ( 
.A(n_2639),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2665),
.B(n_141),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_2650),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2630),
.B(n_141),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2546),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2565),
.B(n_142),
.Y(n_2737)
);

AND2x4_ASAP7_75t_SL g2738 ( 
.A(n_2612),
.B(n_142),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2547),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2650),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2588),
.B(n_143),
.Y(n_2741)
);

OR2x6_ASAP7_75t_SL g2742 ( 
.A(n_2668),
.B(n_143),
.Y(n_2742)
);

AND2x4_ASAP7_75t_L g2743 ( 
.A(n_2610),
.B(n_144),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2573),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2568),
.Y(n_2745)
);

OR2x2_ASAP7_75t_L g2746 ( 
.A(n_2551),
.B(n_144),
.Y(n_2746)
);

INVx2_ASAP7_75t_SL g2747 ( 
.A(n_2617),
.Y(n_2747)
);

NAND2x1p5_ASAP7_75t_L g2748 ( 
.A(n_2608),
.B(n_145),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2557),
.Y(n_2749)
);

INVxp67_ASAP7_75t_L g2750 ( 
.A(n_2607),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2559),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2569),
.B(n_146),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2610),
.B(n_146),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2564),
.Y(n_2754)
);

INVx2_ASAP7_75t_SL g2755 ( 
.A(n_2532),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2625),
.B(n_147),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2626),
.B(n_147),
.Y(n_2757)
);

NAND2x1p5_ASAP7_75t_L g2758 ( 
.A(n_2649),
.B(n_148),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2670),
.B(n_2667),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2602),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2618),
.Y(n_2761)
);

AND2x4_ASAP7_75t_L g2762 ( 
.A(n_2656),
.B(n_148),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2586),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2674),
.B(n_2652),
.Y(n_2764)
);

AND2x4_ASAP7_75t_SL g2765 ( 
.A(n_2747),
.B(n_2671),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2694),
.B(n_2669),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2759),
.B(n_2636),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2691),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2734),
.B(n_2614),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2696),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2673),
.B(n_2633),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2759),
.B(n_2658),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2685),
.B(n_2596),
.Y(n_2773)
);

AND2x4_ASAP7_75t_SL g2774 ( 
.A(n_2760),
.B(n_2671),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2744),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2676),
.B(n_2603),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2715),
.Y(n_2777)
);

NAND4xp25_ASAP7_75t_L g2778 ( 
.A(n_2726),
.B(n_2635),
.C(n_2535),
.D(n_2597),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2734),
.B(n_2628),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2707),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2720),
.B(n_2637),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2679),
.B(n_2661),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2683),
.B(n_2632),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2681),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2740),
.B(n_2599),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2706),
.B(n_2729),
.Y(n_2786)
);

OAI211xp5_ASAP7_75t_L g2787 ( 
.A1(n_2686),
.A2(n_2725),
.B(n_2731),
.C(n_2733),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2682),
.B(n_2613),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2680),
.B(n_2645),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2722),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2690),
.B(n_2662),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2711),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2695),
.B(n_2663),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2688),
.B(n_2571),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2714),
.B(n_2634),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2750),
.B(n_2615),
.Y(n_2796)
);

INVxp67_ASAP7_75t_SL g2797 ( 
.A(n_2678),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2745),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2689),
.B(n_2659),
.Y(n_2799)
);

INVx1_ASAP7_75t_SL g2800 ( 
.A(n_2732),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2692),
.B(n_2624),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2687),
.B(n_2703),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2693),
.B(n_2684),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2718),
.Y(n_2804)
);

INVxp67_ASAP7_75t_SL g2805 ( 
.A(n_2697),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2728),
.B(n_2621),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2677),
.B(n_2591),
.Y(n_2807)
);

OR2x2_ASAP7_75t_L g2808 ( 
.A(n_2736),
.B(n_2641),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2739),
.B(n_2749),
.Y(n_2809)
);

NAND2x1p5_ASAP7_75t_L g2810 ( 
.A(n_2727),
.B(n_2539),
.Y(n_2810)
);

NOR2x1_ASAP7_75t_L g2811 ( 
.A(n_2701),
.B(n_2643),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2763),
.B(n_2591),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2751),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2754),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2753),
.B(n_2619),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2702),
.B(n_2619),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2705),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2716),
.B(n_2648),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2761),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2712),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2709),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2719),
.B(n_2654),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2708),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2699),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2698),
.Y(n_2825)
);

OR2x2_ASAP7_75t_L g2826 ( 
.A(n_2756),
.B(n_2666),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2700),
.Y(n_2827)
);

OR2x2_ASAP7_75t_L g2828 ( 
.A(n_2746),
.B(n_2627),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2723),
.B(n_2592),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2737),
.B(n_2653),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2752),
.Y(n_2831)
);

OR2x2_ASAP7_75t_L g2832 ( 
.A(n_2735),
.B(n_2664),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2717),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2757),
.B(n_2655),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2762),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2721),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2762),
.B(n_2558),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2743),
.B(n_2580),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2704),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2743),
.Y(n_2840)
);

AND2x2_ASAP7_75t_SL g2841 ( 
.A(n_2713),
.B(n_2561),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2742),
.A2(n_2543),
.B1(n_2561),
.B2(n_151),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2755),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2741),
.B(n_900),
.Y(n_2844)
);

AND2x4_ASAP7_75t_SL g2845 ( 
.A(n_2724),
.B(n_2730),
.Y(n_2845)
);

NAND4xp25_ASAP7_75t_L g2846 ( 
.A(n_2778),
.B(n_2710),
.C(n_2675),
.D(n_2748),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2797),
.B(n_2758),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2820),
.B(n_2738),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2764),
.B(n_149),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2803),
.B(n_149),
.Y(n_2850)
);

NAND2x1p5_ASAP7_75t_L g2851 ( 
.A(n_2811),
.B(n_150),
.Y(n_2851)
);

OR2x2_ASAP7_75t_L g2852 ( 
.A(n_2769),
.B(n_150),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2809),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2768),
.Y(n_2854)
);

AND2x4_ASAP7_75t_L g2855 ( 
.A(n_2786),
.B(n_151),
.Y(n_2855)
);

INVxp67_ASAP7_75t_L g2856 ( 
.A(n_2793),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2823),
.B(n_152),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2770),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2805),
.B(n_152),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2791),
.B(n_153),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2794),
.B(n_153),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2780),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2784),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2814),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2782),
.B(n_910),
.Y(n_2865)
);

NAND2x2_ASAP7_75t_L g2866 ( 
.A(n_2837),
.B(n_155),
.Y(n_2866)
);

HB1xp67_ASAP7_75t_L g2867 ( 
.A(n_2779),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2826),
.B(n_155),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2819),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2802),
.B(n_911),
.Y(n_2870)
);

NAND4xp25_ASAP7_75t_L g2871 ( 
.A(n_2787),
.B(n_911),
.C(n_912),
.D(n_910),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2792),
.Y(n_2872)
);

OR2x2_ASAP7_75t_L g2873 ( 
.A(n_2807),
.B(n_156),
.Y(n_2873)
);

INVx2_ASAP7_75t_SL g2874 ( 
.A(n_2774),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2771),
.B(n_156),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2804),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2798),
.Y(n_2877)
);

OAI21xp33_ASAP7_75t_L g2878 ( 
.A1(n_2842),
.A2(n_157),
.B(n_158),
.Y(n_2878)
);

NOR2x1_ASAP7_75t_L g2879 ( 
.A(n_2829),
.B(n_157),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2835),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_SL g2881 ( 
.A(n_2800),
.B(n_159),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2766),
.B(n_160),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2786),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2813),
.Y(n_2884)
);

AOI22xp33_ASAP7_75t_L g2885 ( 
.A1(n_2840),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2817),
.Y(n_2886)
);

NOR2xp67_ASAP7_75t_L g2887 ( 
.A(n_2843),
.B(n_162),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_2781),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2834),
.B(n_164),
.Y(n_2889)
);

INVx3_ASAP7_75t_SL g2890 ( 
.A(n_2765),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2767),
.B(n_899),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2772),
.B(n_900),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2773),
.B(n_2775),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2808),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2777),
.B(n_164),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2790),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2789),
.B(n_902),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2822),
.B(n_165),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2801),
.B(n_2815),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2785),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2812),
.Y(n_2901)
);

INVx1_ASAP7_75t_SL g2902 ( 
.A(n_2838),
.Y(n_2902)
);

OR2x2_ASAP7_75t_L g2903 ( 
.A(n_2795),
.B(n_166),
.Y(n_2903)
);

NAND2x1_ASAP7_75t_L g2904 ( 
.A(n_2806),
.B(n_167),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2816),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2830),
.B(n_909),
.Y(n_2906)
);

INVxp67_ASAP7_75t_L g2907 ( 
.A(n_2783),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2785),
.B(n_168),
.Y(n_2908)
);

INVx1_ASAP7_75t_SL g2909 ( 
.A(n_2845),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2799),
.B(n_2821),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2806),
.Y(n_2911)
);

A2O1A1Ixp33_ASAP7_75t_L g2912 ( 
.A1(n_2841),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2796),
.Y(n_2913)
);

INVxp67_ASAP7_75t_SL g2914 ( 
.A(n_2832),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2828),
.B(n_169),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2818),
.B(n_915),
.Y(n_2916)
);

NAND3xp33_ASAP7_75t_L g2917 ( 
.A(n_2839),
.B(n_2776),
.C(n_2825),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2831),
.B(n_170),
.Y(n_2918)
);

OR2x2_ASAP7_75t_L g2919 ( 
.A(n_2824),
.B(n_171),
.Y(n_2919)
);

OR2x2_ASAP7_75t_L g2920 ( 
.A(n_2833),
.B(n_171),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2788),
.Y(n_2921)
);

AND2x2_ASAP7_75t_L g2922 ( 
.A(n_2827),
.B(n_2836),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2788),
.B(n_172),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2844),
.B(n_173),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2810),
.B(n_173),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2768),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2782),
.B(n_893),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2782),
.B(n_893),
.Y(n_2928)
);

OAI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2787),
.A2(n_174),
.B(n_176),
.Y(n_2929)
);

INVx1_ASAP7_75t_SL g2930 ( 
.A(n_2800),
.Y(n_2930)
);

OAI322xp33_ASAP7_75t_L g2931 ( 
.A1(n_2888),
.A2(n_200),
.A3(n_183),
.B1(n_208),
.B2(n_216),
.C1(n_192),
.C2(n_174),
.Y(n_2931)
);

NAND4xp25_ASAP7_75t_L g2932 ( 
.A(n_2871),
.B(n_178),
.C(n_176),
.D(n_177),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2913),
.B(n_177),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2914),
.B(n_178),
.Y(n_2934)
);

INVx3_ASAP7_75t_L g2935 ( 
.A(n_2853),
.Y(n_2935)
);

AND2x2_ASAP7_75t_SL g2936 ( 
.A(n_2855),
.B(n_179),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2854),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2901),
.B(n_179),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2858),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2862),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2893),
.B(n_2905),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2883),
.B(n_180),
.Y(n_2942)
);

NAND4xp25_ASAP7_75t_L g2943 ( 
.A(n_2929),
.B(n_182),
.C(n_180),
.D(n_181),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2863),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2878),
.A2(n_184),
.B1(n_181),
.B2(n_182),
.Y(n_2945)
);

OR2x2_ASAP7_75t_L g2946 ( 
.A(n_2867),
.B(n_913),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2910),
.B(n_184),
.Y(n_2947)
);

OR2x2_ASAP7_75t_L g2948 ( 
.A(n_2894),
.B(n_916),
.Y(n_2948)
);

NOR2xp67_ASAP7_75t_SL g2949 ( 
.A(n_2846),
.B(n_186),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2872),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2866),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2951)
);

NOR2xp33_ASAP7_75t_L g2952 ( 
.A(n_2890),
.B(n_2909),
.Y(n_2952)
);

INVx2_ASAP7_75t_SL g2953 ( 
.A(n_2930),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2899),
.B(n_187),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2876),
.Y(n_2955)
);

AOI22xp5_ASAP7_75t_L g2956 ( 
.A1(n_2912),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2917),
.B(n_890),
.Y(n_2957)
);

AO221x1_ASAP7_75t_L g2958 ( 
.A1(n_2884),
.A2(n_2926),
.B1(n_2921),
.B2(n_2896),
.C(n_2856),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2879),
.B(n_890),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_L g2960 ( 
.A(n_2873),
.B(n_189),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2886),
.Y(n_2961)
);

AOI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2898),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2864),
.Y(n_2963)
);

AOI21xp33_ASAP7_75t_L g2964 ( 
.A1(n_2904),
.A2(n_191),
.B(n_193),
.Y(n_2964)
);

AOI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_2847),
.A2(n_194),
.B(n_195),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2869),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2877),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2900),
.Y(n_2968)
);

BUFx2_ASAP7_75t_L g2969 ( 
.A(n_2911),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2922),
.Y(n_2970)
);

OAI21xp33_ASAP7_75t_SL g2971 ( 
.A1(n_2861),
.A2(n_194),
.B(n_196),
.Y(n_2971)
);

OAI22xp33_ASAP7_75t_L g2972 ( 
.A1(n_2851),
.A2(n_2880),
.B1(n_2849),
.B2(n_2852),
.Y(n_2972)
);

AOI211xp5_ASAP7_75t_L g2973 ( 
.A1(n_2881),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2907),
.B(n_198),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2902),
.B(n_199),
.Y(n_2975)
);

AOI21xp33_ASAP7_75t_L g2976 ( 
.A1(n_2925),
.A2(n_2868),
.B(n_2859),
.Y(n_2976)
);

NOR2xp67_ASAP7_75t_L g2977 ( 
.A(n_2874),
.B(n_2875),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2903),
.Y(n_2978)
);

AOI322xp5_ASAP7_75t_L g2979 ( 
.A1(n_2857),
.A2(n_204),
.A3(n_203),
.B1(n_201),
.B2(n_199),
.C1(n_200),
.C2(n_202),
.Y(n_2979)
);

AOI321xp33_ASAP7_75t_L g2980 ( 
.A1(n_2885),
.A2(n_205),
.A3(n_207),
.B1(n_203),
.B2(n_204),
.C(n_206),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2889),
.B(n_2915),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2848),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2919),
.Y(n_2983)
);

OAI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2887),
.A2(n_205),
.B(n_206),
.Y(n_2984)
);

OAI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2923),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2860),
.B(n_209),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2895),
.Y(n_2987)
);

OAI21xp33_ASAP7_75t_L g2988 ( 
.A1(n_2908),
.A2(n_2850),
.B(n_2918),
.Y(n_2988)
);

AO21x1_ASAP7_75t_L g2989 ( 
.A1(n_2855),
.A2(n_210),
.B(n_211),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2920),
.Y(n_2990)
);

AOI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2891),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2892),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2897),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2865),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2870),
.B(n_212),
.Y(n_2995)
);

AOI222xp33_ASAP7_75t_L g2996 ( 
.A1(n_2924),
.A2(n_215),
.B1(n_219),
.B2(n_213),
.C1(n_214),
.C2(n_218),
.Y(n_2996)
);

INVxp67_ASAP7_75t_SL g2997 ( 
.A(n_2927),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2928),
.B(n_218),
.Y(n_2998)
);

INVxp67_ASAP7_75t_SL g2999 ( 
.A(n_2882),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2916),
.Y(n_3000)
);

AOI21xp5_ASAP7_75t_SL g3001 ( 
.A1(n_2906),
.A2(n_220),
.B(n_221),
.Y(n_3001)
);

OR2x2_ASAP7_75t_L g3002 ( 
.A(n_2914),
.B(n_916),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2853),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2854),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2883),
.B(n_220),
.Y(n_3005)
);

NAND2xp33_ASAP7_75t_SL g3006 ( 
.A(n_2890),
.B(n_221),
.Y(n_3006)
);

OAI221xp5_ASAP7_75t_L g3007 ( 
.A1(n_2929),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.C(n_226),
.Y(n_3007)
);

OAI32xp33_ASAP7_75t_L g3008 ( 
.A1(n_2871),
.A2(n_227),
.A3(n_223),
.B1(n_226),
.B2(n_228),
.Y(n_3008)
);

AOI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2871),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_3009)
);

INVxp67_ASAP7_75t_L g3010 ( 
.A(n_2867),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2888),
.B(n_229),
.Y(n_3011)
);

A2O1A1Ixp33_ASAP7_75t_SL g3012 ( 
.A1(n_2929),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2854),
.Y(n_3013)
);

INVxp67_ASAP7_75t_L g3014 ( 
.A(n_2867),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2854),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2883),
.B(n_230),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2883),
.B(n_232),
.Y(n_3017)
);

O2A1O1Ixp33_ASAP7_75t_L g3018 ( 
.A1(n_2912),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_3018)
);

INVxp67_ASAP7_75t_L g3019 ( 
.A(n_2867),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2854),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2854),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2854),
.Y(n_3022)
);

AOI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2871),
.A2(n_237),
.B1(n_234),
.B2(n_235),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2854),
.Y(n_3024)
);

A2O1A1Ixp33_ASAP7_75t_L g3025 ( 
.A1(n_2929),
.A2(n_239),
.B(n_240),
.C(n_238),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2888),
.B(n_237),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2914),
.B(n_238),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2854),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2888),
.B(n_239),
.Y(n_3029)
);

OAI21xp5_ASAP7_75t_SL g3030 ( 
.A1(n_2929),
.A2(n_240),
.B(n_241),
.Y(n_3030)
);

AOI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2871),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2878),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2888),
.B(n_245),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2883),
.B(n_245),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2883),
.B(n_246),
.Y(n_3035)
);

AOI21xp33_ASAP7_75t_L g3036 ( 
.A1(n_2929),
.A2(n_246),
.B(n_247),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2888),
.B(n_248),
.Y(n_3037)
);

OAI31xp33_ASAP7_75t_L g3038 ( 
.A1(n_2912),
.A2(n_250),
.A3(n_248),
.B(n_249),
.Y(n_3038)
);

OA21x2_ASAP7_75t_L g3039 ( 
.A1(n_2917),
.A2(n_249),
.B(n_250),
.Y(n_3039)
);

AOI221xp5_ASAP7_75t_L g3040 ( 
.A1(n_3008),
.A2(n_3007),
.B1(n_2931),
.B2(n_3018),
.C(n_2985),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2987),
.B(n_251),
.Y(n_3041)
);

OR2x2_ASAP7_75t_L g3042 ( 
.A(n_3010),
.B(n_251),
.Y(n_3042)
);

OAI222xp33_ASAP7_75t_L g3043 ( 
.A1(n_2949),
.A2(n_2957),
.B1(n_2962),
.B2(n_3023),
.C1(n_3031),
.C2(n_3009),
.Y(n_3043)
);

OAI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_3030),
.A2(n_2956),
.B1(n_3025),
.B2(n_2945),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_3014),
.B(n_253),
.Y(n_3045)
);

OAI21xp33_ASAP7_75t_L g3046 ( 
.A1(n_2943),
.A2(n_256),
.B(n_255),
.Y(n_3046)
);

AOI211xp5_ASAP7_75t_SL g3047 ( 
.A1(n_3036),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_3019),
.B(n_254),
.Y(n_3048)
);

OAI21xp33_ASAP7_75t_SL g3049 ( 
.A1(n_2958),
.A2(n_257),
.B(n_258),
.Y(n_3049)
);

OR2x2_ASAP7_75t_L g3050 ( 
.A(n_2970),
.B(n_257),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2939),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_3012),
.A2(n_259),
.B(n_260),
.Y(n_3052)
);

AOI322xp5_ASAP7_75t_L g3053 ( 
.A1(n_2971),
.A2(n_264),
.A3(n_263),
.B1(n_261),
.B2(n_259),
.C1(n_260),
.C2(n_262),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_2932),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2941),
.B(n_265),
.Y(n_3055)
);

OAI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2965),
.A2(n_265),
.B(n_266),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2944),
.Y(n_3057)
);

NAND4xp25_ASAP7_75t_L g3058 ( 
.A(n_2996),
.B(n_268),
.C(n_266),
.D(n_267),
.Y(n_3058)
);

AOI222xp33_ASAP7_75t_L g3059 ( 
.A1(n_3032),
.A2(n_270),
.B1(n_272),
.B2(n_268),
.C1(n_269),
.C2(n_271),
.Y(n_3059)
);

O2A1O1Ixp33_ASAP7_75t_L g3060 ( 
.A1(n_2959),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_3060)
);

AOI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_3006),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3061)
);

AOI221xp5_ASAP7_75t_L g3062 ( 
.A1(n_3001),
.A2(n_2972),
.B1(n_3038),
.B2(n_2976),
.C(n_2973),
.Y(n_3062)
);

OAI222xp33_ASAP7_75t_L g3063 ( 
.A1(n_2991),
.A2(n_276),
.B1(n_278),
.B2(n_273),
.C1(n_275),
.C2(n_277),
.Y(n_3063)
);

OR2x2_ASAP7_75t_L g3064 ( 
.A(n_2978),
.B(n_276),
.Y(n_3064)
);

OAI21xp33_ASAP7_75t_L g3065 ( 
.A1(n_2979),
.A2(n_279),
.B(n_278),
.Y(n_3065)
);

A2O1A1Ixp33_ASAP7_75t_L g3066 ( 
.A1(n_2980),
.A2(n_2984),
.B(n_2960),
.C(n_2951),
.Y(n_3066)
);

AOI221xp5_ASAP7_75t_L g3067 ( 
.A1(n_2988),
.A2(n_281),
.B1(n_277),
.B2(n_280),
.C(n_282),
.Y(n_3067)
);

OAI22xp33_ASAP7_75t_L g3068 ( 
.A1(n_3039),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3068)
);

AO22x1_ASAP7_75t_L g3069 ( 
.A1(n_2942),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_3069)
);

OAI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2977),
.A2(n_3039),
.B(n_2981),
.Y(n_3070)
);

AOI221xp5_ASAP7_75t_L g3071 ( 
.A1(n_2989),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2936),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_3072)
);

AO21x1_ASAP7_75t_L g3073 ( 
.A1(n_2942),
.A2(n_287),
.B(n_289),
.Y(n_3073)
);

AOI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2964),
.A2(n_289),
.B(n_290),
.Y(n_3074)
);

OAI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_2986),
.A2(n_291),
.B(n_292),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_3011),
.A2(n_291),
.B(n_292),
.Y(n_3076)
);

OAI22xp33_ASAP7_75t_SL g3077 ( 
.A1(n_2934),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_3077)
);

OAI222xp33_ASAP7_75t_L g3078 ( 
.A1(n_2954),
.A2(n_295),
.B1(n_298),
.B2(n_293),
.C1(n_294),
.C2(n_296),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2990),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3079)
);

NAND3xp33_ASAP7_75t_L g3080 ( 
.A(n_2933),
.B(n_299),
.C(n_300),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2955),
.Y(n_3081)
);

AOI211x1_ASAP7_75t_SL g3082 ( 
.A1(n_2938),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_3082)
);

INVxp67_ASAP7_75t_L g3083 ( 
.A(n_3026),
.Y(n_3083)
);

AOI32xp33_ASAP7_75t_L g3084 ( 
.A1(n_3005),
.A2(n_305),
.A3(n_303),
.B1(n_304),
.B2(n_306),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3004),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_SL g3086 ( 
.A1(n_2952),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.Y(n_3086)
);

OAI211xp5_ASAP7_75t_L g3087 ( 
.A1(n_3037),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_3087)
);

OR2x6_ASAP7_75t_L g3088 ( 
.A(n_2953),
.B(n_308),
.Y(n_3088)
);

NOR4xp25_ASAP7_75t_L g3089 ( 
.A(n_3029),
.B(n_311),
.C(n_312),
.D(n_310),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_2982),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_3033),
.A2(n_312),
.B(n_314),
.Y(n_3091)
);

AOI211xp5_ASAP7_75t_L g3092 ( 
.A1(n_2947),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_3092)
);

OAI32xp33_ASAP7_75t_L g3093 ( 
.A1(n_3002),
.A2(n_318),
.A3(n_315),
.B1(n_317),
.B2(n_319),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2975),
.A2(n_317),
.B(n_318),
.Y(n_3094)
);

AOI221xp5_ASAP7_75t_L g3095 ( 
.A1(n_2974),
.A2(n_2999),
.B1(n_2997),
.B2(n_2993),
.C(n_3000),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_3013),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2983),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_3097)
);

O2A1O1Ixp33_ASAP7_75t_L g3098 ( 
.A1(n_2946),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_3098)
);

OAI211xp5_ASAP7_75t_SL g3099 ( 
.A1(n_2998),
.A2(n_325),
.B(n_322),
.C(n_324),
.Y(n_3099)
);

AOI32xp33_ASAP7_75t_L g3100 ( 
.A1(n_3016),
.A2(n_326),
.A3(n_324),
.B1(n_325),
.B2(n_327),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_3003),
.B(n_326),
.Y(n_3101)
);

OAI32xp33_ASAP7_75t_L g3102 ( 
.A1(n_3027),
.A2(n_329),
.A3(n_327),
.B1(n_328),
.B2(n_330),
.Y(n_3102)
);

OAI31xp33_ASAP7_75t_L g3103 ( 
.A1(n_3017),
.A2(n_332),
.A3(n_330),
.B(n_331),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2994),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_3104)
);

OAI32xp33_ASAP7_75t_L g3105 ( 
.A1(n_2948),
.A2(n_335),
.A3(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_3105)
);

AOI321xp33_ASAP7_75t_L g3106 ( 
.A1(n_3034),
.A2(n_337),
.A3(n_339),
.B1(n_334),
.B2(n_336),
.C(n_338),
.Y(n_3106)
);

AOI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2992),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_3107)
);

NOR3xp33_ASAP7_75t_L g3108 ( 
.A(n_3035),
.B(n_340),
.C(n_341),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_3020),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3021),
.Y(n_3110)
);

OAI22x1_ASAP7_75t_L g3111 ( 
.A1(n_2969),
.A2(n_343),
.B1(n_340),
.B2(n_342),
.Y(n_3111)
);

AOI32xp33_ASAP7_75t_SL g3112 ( 
.A1(n_3028),
.A2(n_344),
.A3(n_342),
.B1(n_343),
.B2(n_346),
.Y(n_3112)
);

OAI211xp5_ASAP7_75t_L g3113 ( 
.A1(n_2995),
.A2(n_347),
.B(n_344),
.C(n_346),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_2935),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3114)
);

AOI22xp5_ASAP7_75t_L g3115 ( 
.A1(n_3003),
.A2(n_3024),
.B1(n_3022),
.B2(n_2968),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2937),
.Y(n_3116)
);

OAI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2940),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3117)
);

AOI221xp5_ASAP7_75t_L g3118 ( 
.A1(n_2961),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.C(n_354),
.Y(n_3118)
);

AOI22xp5_ASAP7_75t_L g3119 ( 
.A1(n_2967),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3119)
);

INVxp67_ASAP7_75t_L g3120 ( 
.A(n_2950),
.Y(n_3120)
);

AOI222xp33_ASAP7_75t_L g3121 ( 
.A1(n_2963),
.A2(n_358),
.B1(n_361),
.B2(n_356),
.C1(n_357),
.C2(n_359),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2966),
.A2(n_359),
.B1(n_356),
.B2(n_358),
.Y(n_3122)
);

AOI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_3015),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2937),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2939),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2939),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2957),
.A2(n_362),
.B(n_364),
.Y(n_3127)
);

AOI222xp33_ASAP7_75t_L g3128 ( 
.A1(n_3030),
.A2(n_366),
.B1(n_368),
.B2(n_364),
.C1(n_365),
.C2(n_367),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2988),
.B(n_901),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2939),
.Y(n_3130)
);

AOI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_3030),
.A2(n_368),
.B1(n_365),
.B2(n_367),
.Y(n_3131)
);

OAI21xp33_ASAP7_75t_L g3132 ( 
.A1(n_3030),
.A2(n_371),
.B(n_370),
.Y(n_3132)
);

OAI211xp5_ASAP7_75t_L g3133 ( 
.A1(n_2996),
.A2(n_372),
.B(n_369),
.C(n_370),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2937),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2939),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2939),
.Y(n_3136)
);

AOI221x1_ASAP7_75t_L g3137 ( 
.A1(n_3001),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.C(n_375),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2957),
.A2(n_374),
.B(n_375),
.Y(n_3138)
);

AOI21xp33_ASAP7_75t_L g3139 ( 
.A1(n_2996),
.A2(n_376),
.B(n_377),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2939),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2987),
.B(n_376),
.Y(n_3141)
);

HB1xp67_ASAP7_75t_L g3142 ( 
.A(n_3010),
.Y(n_3142)
);

OAI21xp33_ASAP7_75t_L g3143 ( 
.A1(n_3030),
.A2(n_379),
.B(n_378),
.Y(n_3143)
);

INVx1_ASAP7_75t_SL g3144 ( 
.A(n_2953),
.Y(n_3144)
);

INVxp67_ASAP7_75t_L g3145 ( 
.A(n_2981),
.Y(n_3145)
);

AOI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2957),
.A2(n_377),
.B(n_378),
.Y(n_3146)
);

INVx1_ASAP7_75t_SL g3147 ( 
.A(n_2953),
.Y(n_3147)
);

NAND3xp33_ASAP7_75t_L g3148 ( 
.A(n_3038),
.B(n_379),
.C(n_380),
.Y(n_3148)
);

AOI321xp33_ASAP7_75t_L g3149 ( 
.A1(n_3007),
.A2(n_383),
.A3(n_385),
.B1(n_380),
.B2(n_382),
.C(n_384),
.Y(n_3149)
);

AOI22xp5_ASAP7_75t_SL g3150 ( 
.A1(n_2942),
.A2(n_387),
.B1(n_388),
.B2(n_386),
.Y(n_3150)
);

OA33x2_ASAP7_75t_L g3151 ( 
.A1(n_2985),
.A2(n_387),
.A3(n_389),
.B1(n_383),
.B2(n_386),
.B3(n_388),
.Y(n_3151)
);

OAI211xp5_ASAP7_75t_SL g3152 ( 
.A1(n_2996),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_2988),
.B(n_888),
.Y(n_3153)
);

AOI221x1_ASAP7_75t_L g3154 ( 
.A1(n_3001),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.C(n_395),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2939),
.Y(n_3155)
);

NAND3xp33_ASAP7_75t_L g3156 ( 
.A(n_3038),
.B(n_393),
.C(n_395),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_SL g3157 ( 
.A1(n_3007),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2939),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_L g3159 ( 
.A(n_2988),
.B(n_897),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2939),
.Y(n_3160)
);

NOR3x1_ASAP7_75t_L g3161 ( 
.A(n_3030),
.B(n_397),
.C(n_399),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_3062),
.A2(n_400),
.B(n_401),
.Y(n_3162)
);

NOR3x1_ASAP7_75t_L g3163 ( 
.A(n_3058),
.B(n_400),
.C(n_401),
.Y(n_3163)
);

NOR3xp33_ASAP7_75t_L g3164 ( 
.A(n_3139),
.B(n_404),
.C(n_405),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_3083),
.B(n_406),
.Y(n_3165)
);

AOI221xp5_ASAP7_75t_L g3166 ( 
.A1(n_3089),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.C(n_409),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3051),
.Y(n_3167)
);

AOI22xp5_ASAP7_75t_L g3168 ( 
.A1(n_3148),
.A2(n_3156),
.B1(n_3133),
.B2(n_3044),
.Y(n_3168)
);

AOI322xp5_ASAP7_75t_L g3169 ( 
.A1(n_3065),
.A2(n_892),
.A3(n_887),
.B1(n_894),
.B2(n_895),
.C1(n_889),
.C2(n_886),
.Y(n_3169)
);

AOI221xp5_ASAP7_75t_L g3170 ( 
.A1(n_3049),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.C(n_411),
.Y(n_3170)
);

NAND4xp75_ASAP7_75t_L g3171 ( 
.A(n_3161),
.B(n_412),
.C(n_410),
.D(n_411),
.Y(n_3171)
);

NAND4xp25_ASAP7_75t_L g3172 ( 
.A(n_3149),
.B(n_414),
.C(n_412),
.D(n_413),
.Y(n_3172)
);

AOI211xp5_ASAP7_75t_L g3173 ( 
.A1(n_3043),
.A2(n_416),
.B(n_413),
.C(n_415),
.Y(n_3173)
);

NAND4xp25_ASAP7_75t_L g3174 ( 
.A(n_3106),
.B(n_417),
.C(n_415),
.D(n_416),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3057),
.Y(n_3175)
);

NAND3xp33_ASAP7_75t_SL g3176 ( 
.A(n_3040),
.B(n_419),
.C(n_420),
.Y(n_3176)
);

OAI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_3066),
.A2(n_420),
.B(n_421),
.Y(n_3177)
);

AOI22xp5_ASAP7_75t_SL g3178 ( 
.A1(n_3077),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3178)
);

NAND3xp33_ASAP7_75t_SL g3179 ( 
.A(n_3070),
.B(n_422),
.C(n_423),
.Y(n_3179)
);

OAI21xp5_ASAP7_75t_SL g3180 ( 
.A1(n_3131),
.A2(n_425),
.B(n_426),
.Y(n_3180)
);

OAI21xp33_ASAP7_75t_L g3181 ( 
.A1(n_3132),
.A2(n_425),
.B(n_426),
.Y(n_3181)
);

OAI21xp33_ASAP7_75t_L g3182 ( 
.A1(n_3143),
.A2(n_427),
.B(n_428),
.Y(n_3182)
);

NOR2xp67_ASAP7_75t_L g3183 ( 
.A(n_3142),
.B(n_886),
.Y(n_3183)
);

AOI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_3152),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_3184)
);

INVx1_ASAP7_75t_SL g3185 ( 
.A(n_3144),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_3056),
.A2(n_430),
.B(n_431),
.Y(n_3186)
);

A2O1A1Ixp33_ASAP7_75t_L g3187 ( 
.A1(n_3084),
.A2(n_433),
.B(n_431),
.C(n_432),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_3052),
.A2(n_3074),
.B(n_3098),
.Y(n_3188)
);

BUFx2_ASAP7_75t_SL g3189 ( 
.A(n_3147),
.Y(n_3189)
);

NAND3xp33_ASAP7_75t_SL g3190 ( 
.A(n_3092),
.B(n_432),
.C(n_434),
.Y(n_3190)
);

NAND4xp25_ASAP7_75t_L g3191 ( 
.A(n_3128),
.B(n_437),
.C(n_435),
.D(n_436),
.Y(n_3191)
);

AOI221xp5_ASAP7_75t_L g3192 ( 
.A1(n_3071),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.C(n_438),
.Y(n_3192)
);

NAND4xp25_ASAP7_75t_SL g3193 ( 
.A(n_3100),
.B(n_441),
.C(n_439),
.D(n_440),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_SL g3194 ( 
.A(n_3095),
.B(n_439),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3145),
.B(n_441),
.Y(n_3195)
);

AOI221xp5_ASAP7_75t_L g3196 ( 
.A1(n_3129),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.C(n_445),
.Y(n_3196)
);

AOI221xp5_ASAP7_75t_L g3197 ( 
.A1(n_3153),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.C(n_446),
.Y(n_3197)
);

O2A1O1Ixp5_ASAP7_75t_L g3198 ( 
.A1(n_3073),
.A2(n_448),
.B(n_446),
.C(n_447),
.Y(n_3198)
);

OAI211xp5_ASAP7_75t_L g3199 ( 
.A1(n_3137),
.A2(n_449),
.B(n_447),
.C(n_448),
.Y(n_3199)
);

AOI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_3157),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_3115),
.B(n_452),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_3120),
.B(n_453),
.Y(n_3202)
);

OAI32xp33_ASAP7_75t_L g3203 ( 
.A1(n_3082),
.A2(n_456),
.A3(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_3203)
);

OAI221xp5_ASAP7_75t_L g3204 ( 
.A1(n_3151),
.A2(n_458),
.B1(n_454),
.B2(n_457),
.C(n_459),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3081),
.Y(n_3205)
);

NAND4xp25_ASAP7_75t_L g3206 ( 
.A(n_3054),
.B(n_462),
.C(n_458),
.D(n_461),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3085),
.Y(n_3207)
);

AOI211xp5_ASAP7_75t_L g3208 ( 
.A1(n_3086),
.A2(n_463),
.B(n_461),
.C(n_462),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_3124),
.Y(n_3209)
);

OAI221xp5_ASAP7_75t_L g3210 ( 
.A1(n_3075),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.C(n_467),
.Y(n_3210)
);

OAI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3076),
.A2(n_464),
.B(n_465),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_3041),
.B(n_466),
.Y(n_3212)
);

OAI211xp5_ASAP7_75t_L g3213 ( 
.A1(n_3154),
.A2(n_469),
.B(n_467),
.C(n_468),
.Y(n_3213)
);

AOI221xp5_ASAP7_75t_L g3214 ( 
.A1(n_3159),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.C(n_471),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_3134),
.B(n_3116),
.Y(n_3215)
);

AOI21xp33_ASAP7_75t_L g3216 ( 
.A1(n_3121),
.A2(n_912),
.B(n_470),
.Y(n_3216)
);

OAI21xp33_ASAP7_75t_L g3217 ( 
.A1(n_3046),
.A2(n_472),
.B(n_473),
.Y(n_3217)
);

NAND4xp25_ASAP7_75t_L g3218 ( 
.A(n_3072),
.B(n_474),
.C(n_472),
.D(n_473),
.Y(n_3218)
);

NAND4xp25_ASAP7_75t_SL g3219 ( 
.A(n_3108),
.B(n_477),
.C(n_474),
.D(n_476),
.Y(n_3219)
);

NOR3x1_ASAP7_75t_L g3220 ( 
.A(n_3069),
.B(n_476),
.C(n_477),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_3068),
.A2(n_478),
.B(n_479),
.Y(n_3221)
);

OAI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_3091),
.A2(n_478),
.B(n_479),
.Y(n_3222)
);

A2O1A1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_3060),
.A2(n_483),
.B(n_480),
.C(n_481),
.Y(n_3223)
);

OAI221xp5_ASAP7_75t_L g3224 ( 
.A1(n_3103),
.A2(n_484),
.B1(n_481),
.B2(n_483),
.C(n_486),
.Y(n_3224)
);

AOI211xp5_ASAP7_75t_L g3225 ( 
.A1(n_3063),
.A2(n_487),
.B(n_484),
.C(n_486),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_3127),
.A2(n_487),
.B(n_488),
.Y(n_3226)
);

AOI221xp5_ASAP7_75t_L g3227 ( 
.A1(n_3067),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.C(n_491),
.Y(n_3227)
);

AOI222xp33_ASAP7_75t_L g3228 ( 
.A1(n_3099),
.A2(n_491),
.B1(n_493),
.B2(n_489),
.C1(n_490),
.C2(n_492),
.Y(n_3228)
);

AOI22xp5_ASAP7_75t_L g3229 ( 
.A1(n_3118),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_3229)
);

O2A1O1Ixp33_ASAP7_75t_L g3230 ( 
.A1(n_3078),
.A2(n_3087),
.B(n_3102),
.C(n_3093),
.Y(n_3230)
);

OAI21xp33_ASAP7_75t_L g3231 ( 
.A1(n_3053),
.A2(n_495),
.B(n_496),
.Y(n_3231)
);

AOI221xp5_ASAP7_75t_L g3232 ( 
.A1(n_3094),
.A2(n_498),
.B1(n_495),
.B2(n_497),
.C(n_499),
.Y(n_3232)
);

OAI31xp33_ASAP7_75t_L g3233 ( 
.A1(n_3113),
.A2(n_500),
.A3(n_497),
.B(n_499),
.Y(n_3233)
);

A2O1A1Ixp33_ASAP7_75t_L g3234 ( 
.A1(n_3138),
.A2(n_504),
.B(n_501),
.C(n_503),
.Y(n_3234)
);

AOI221xp5_ASAP7_75t_SL g3235 ( 
.A1(n_3111),
.A2(n_505),
.B1(n_501),
.B2(n_503),
.C(n_506),
.Y(n_3235)
);

OAI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_3080),
.A2(n_505),
.B(n_507),
.Y(n_3236)
);

OAI211xp5_ASAP7_75t_SL g3237 ( 
.A1(n_3141),
.A2(n_913),
.B(n_509),
.C(n_507),
.Y(n_3237)
);

NOR2xp33_ASAP7_75t_L g3238 ( 
.A(n_3055),
.B(n_508),
.Y(n_3238)
);

OAI22xp33_ASAP7_75t_L g3239 ( 
.A1(n_3047),
.A2(n_511),
.B1(n_508),
.B2(n_510),
.Y(n_3239)
);

NAND4xp75_ASAP7_75t_L g3240 ( 
.A(n_3061),
.B(n_512),
.C(n_510),
.D(n_511),
.Y(n_3240)
);

AOI21xp33_ASAP7_75t_SL g3241 ( 
.A1(n_3088),
.A2(n_513),
.B(n_514),
.Y(n_3241)
);

OAI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3146),
.A2(n_515),
.B(n_516),
.Y(n_3242)
);

NAND3xp33_ASAP7_75t_L g3243 ( 
.A(n_3059),
.B(n_905),
.C(n_516),
.Y(n_3243)
);

AOI21xp33_ASAP7_75t_L g3244 ( 
.A1(n_3105),
.A2(n_517),
.B(n_518),
.Y(n_3244)
);

NOR2x1_ASAP7_75t_L g3245 ( 
.A(n_3088),
.B(n_519),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_3088),
.Y(n_3246)
);

NAND3xp33_ASAP7_75t_L g3247 ( 
.A(n_3123),
.B(n_519),
.C(n_520),
.Y(n_3247)
);

AOI221xp5_ASAP7_75t_L g3248 ( 
.A1(n_3104),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.C(n_523),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3117),
.A2(n_523),
.B(n_524),
.Y(n_3249)
);

AOI22xp5_ASAP7_75t_L g3250 ( 
.A1(n_3114),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_3097),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.Y(n_3251)
);

OAI21xp5_ASAP7_75t_SL g3252 ( 
.A1(n_3079),
.A2(n_528),
.B(n_529),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3096),
.Y(n_3253)
);

AOI211xp5_ASAP7_75t_SL g3254 ( 
.A1(n_3119),
.A2(n_905),
.B(n_530),
.C(n_528),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_3109),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_3045),
.B(n_3048),
.Y(n_3256)
);

AOI221xp5_ASAP7_75t_L g3257 ( 
.A1(n_3090),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.C(n_532),
.Y(n_3257)
);

AOI211xp5_ASAP7_75t_SL g3258 ( 
.A1(n_3122),
.A2(n_904),
.B(n_533),
.C(n_531),
.Y(n_3258)
);

AOI221x1_ASAP7_75t_SL g3259 ( 
.A1(n_3112),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.C(n_535),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_SL g3260 ( 
.A1(n_3101),
.A2(n_536),
.B(n_537),
.Y(n_3260)
);

AOI221xp5_ASAP7_75t_L g3261 ( 
.A1(n_3107),
.A2(n_539),
.B1(n_537),
.B2(n_538),
.C(n_540),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_3042),
.B(n_538),
.Y(n_3262)
);

NAND3xp33_ASAP7_75t_L g3263 ( 
.A(n_3150),
.B(n_902),
.C(n_539),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3110),
.B(n_541),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_3160),
.B(n_542),
.Y(n_3265)
);

AOI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_3125),
.A2(n_545),
.B1(n_542),
.B2(n_543),
.Y(n_3266)
);

AOI22xp33_ASAP7_75t_SL g3267 ( 
.A1(n_3064),
.A2(n_547),
.B1(n_545),
.B2(n_546),
.Y(n_3267)
);

NAND3xp33_ASAP7_75t_L g3268 ( 
.A(n_3050),
.B(n_898),
.C(n_546),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3126),
.A2(n_547),
.B(n_548),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_SL g3270 ( 
.A(n_3130),
.B(n_549),
.Y(n_3270)
);

NAND2xp33_ASAP7_75t_SL g3271 ( 
.A(n_3135),
.B(n_3136),
.Y(n_3271)
);

NOR3x1_ASAP7_75t_L g3272 ( 
.A(n_3140),
.B(n_550),
.C(n_551),
.Y(n_3272)
);

AOI321xp33_ASAP7_75t_L g3273 ( 
.A1(n_3155),
.A2(n_552),
.A3(n_554),
.B1(n_550),
.B2(n_551),
.C(n_553),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3158),
.B(n_554),
.Y(n_3274)
);

OAI211xp5_ASAP7_75t_SL g3275 ( 
.A1(n_3062),
.A2(n_897),
.B(n_557),
.C(n_555),
.Y(n_3275)
);

NOR2x1_ASAP7_75t_L g3276 ( 
.A(n_3070),
.B(n_556),
.Y(n_3276)
);

AOI221xp5_ASAP7_75t_L g3277 ( 
.A1(n_3062),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.C(n_560),
.Y(n_3277)
);

AOI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3148),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_3278)
);

OAI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_3148),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3145),
.B(n_561),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3051),
.Y(n_3281)
);

AOI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_3148),
.A2(n_565),
.B1(n_562),
.B2(n_564),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3051),
.Y(n_3283)
);

NAND3xp33_ASAP7_75t_L g3284 ( 
.A(n_3062),
.B(n_896),
.C(n_566),
.Y(n_3284)
);

AOI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3148),
.A2(n_569),
.B1(n_566),
.B2(n_568),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3145),
.B(n_568),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_SL g3287 ( 
.A1(n_3062),
.A2(n_569),
.B(n_570),
.Y(n_3287)
);

AND4x1_ASAP7_75t_L g3288 ( 
.A(n_3062),
.B(n_572),
.C(n_570),
.D(n_571),
.Y(n_3288)
);

NAND3xp33_ASAP7_75t_L g3289 ( 
.A(n_3062),
.B(n_571),
.C(n_573),
.Y(n_3289)
);

NAND4xp25_ASAP7_75t_L g3290 ( 
.A(n_3149),
.B(n_575),
.C(n_573),
.D(n_574),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_3083),
.B(n_574),
.Y(n_3291)
);

NAND4xp25_ASAP7_75t_L g3292 ( 
.A(n_3149),
.B(n_578),
.C(n_576),
.D(n_577),
.Y(n_3292)
);

OAI21xp33_ASAP7_75t_L g3293 ( 
.A1(n_3065),
.A2(n_578),
.B(n_579),
.Y(n_3293)
);

AOI211xp5_ASAP7_75t_L g3294 ( 
.A1(n_3062),
.A2(n_581),
.B(n_579),
.C(n_580),
.Y(n_3294)
);

AND4x1_ASAP7_75t_L g3295 ( 
.A(n_3062),
.B(n_583),
.C(n_580),
.D(n_582),
.Y(n_3295)
);

AOI322xp5_ASAP7_75t_L g3296 ( 
.A1(n_3065),
.A2(n_587),
.A3(n_586),
.B1(n_584),
.B2(n_582),
.C1(n_583),
.C2(n_585),
.Y(n_3296)
);

NAND4xp75_ASAP7_75t_L g3297 ( 
.A(n_3161),
.B(n_587),
.C(n_585),
.D(n_586),
.Y(n_3297)
);

AOI221xp5_ASAP7_75t_L g3298 ( 
.A1(n_3062),
.A2(n_590),
.B1(n_588),
.B2(n_589),
.C(n_591),
.Y(n_3298)
);

O2A1O1Ixp33_ASAP7_75t_L g3299 ( 
.A1(n_3043),
.A2(n_590),
.B(n_588),
.C(n_589),
.Y(n_3299)
);

OAI221xp5_ASAP7_75t_L g3300 ( 
.A1(n_3062),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.C(n_595),
.Y(n_3300)
);

AO21x1_ASAP7_75t_L g3301 ( 
.A1(n_3070),
.A2(n_592),
.B(n_595),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3148),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.Y(n_3302)
);

NOR3xp33_ASAP7_75t_L g3303 ( 
.A(n_3139),
.B(n_596),
.C(n_597),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3049),
.B(n_598),
.Y(n_3304)
);

OAI311xp33_ASAP7_75t_L g3305 ( 
.A1(n_3058),
.A2(n_896),
.A3(n_601),
.B1(n_599),
.C1(n_600),
.Y(n_3305)
);

NAND4xp25_ASAP7_75t_L g3306 ( 
.A(n_3149),
.B(n_602),
.C(n_599),
.D(n_600),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3145),
.B(n_602),
.Y(n_3307)
);

AOI221xp5_ASAP7_75t_L g3308 ( 
.A1(n_3062),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.C(n_606),
.Y(n_3308)
);

AOI221xp5_ASAP7_75t_L g3309 ( 
.A1(n_3062),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.C(n_606),
.Y(n_3309)
);

NOR4xp25_ASAP7_75t_L g3310 ( 
.A(n_3133),
.B(n_610),
.C(n_608),
.D(n_609),
.Y(n_3310)
);

O2A1O1Ixp5_ASAP7_75t_L g3311 ( 
.A1(n_3070),
.A2(n_610),
.B(n_608),
.C(n_609),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_3083),
.B(n_611),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3062),
.A2(n_611),
.B(n_612),
.Y(n_3313)
);

NAND3xp33_ASAP7_75t_L g3314 ( 
.A(n_3062),
.B(n_895),
.C(n_613),
.Y(n_3314)
);

NAND4xp25_ASAP7_75t_L g3315 ( 
.A(n_3149),
.B(n_616),
.C(n_613),
.D(n_614),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3145),
.B(n_614),
.Y(n_3316)
);

OAI211xp5_ASAP7_75t_L g3317 ( 
.A1(n_3062),
.A2(n_620),
.B(n_618),
.C(n_619),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3051),
.Y(n_3318)
);

AOI221xp5_ASAP7_75t_L g3319 ( 
.A1(n_3062),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.C(n_621),
.Y(n_3319)
);

AOI221xp5_ASAP7_75t_L g3320 ( 
.A1(n_3062),
.A2(n_623),
.B1(n_621),
.B2(n_622),
.C(n_624),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_L g3321 ( 
.A(n_3083),
.B(n_623),
.Y(n_3321)
);

OA21x2_ASAP7_75t_SL g3322 ( 
.A1(n_3151),
.A2(n_625),
.B(n_626),
.Y(n_3322)
);

NOR3xp33_ASAP7_75t_L g3323 ( 
.A(n_3139),
.B(n_625),
.C(n_626),
.Y(n_3323)
);

OAI21xp33_ASAP7_75t_L g3324 ( 
.A1(n_3065),
.A2(n_627),
.B(n_628),
.Y(n_3324)
);

AOI221xp5_ASAP7_75t_L g3325 ( 
.A1(n_3062),
.A2(n_629),
.B1(n_627),
.B2(n_628),
.C(n_630),
.Y(n_3325)
);

OAI21xp33_ASAP7_75t_L g3326 ( 
.A1(n_3065),
.A2(n_629),
.B(n_631),
.Y(n_3326)
);

OAI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3049),
.A2(n_631),
.B(n_633),
.Y(n_3327)
);

AOI211xp5_ASAP7_75t_L g3328 ( 
.A1(n_3062),
.A2(n_636),
.B(n_634),
.C(n_635),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3051),
.Y(n_3329)
);

NAND4xp25_ASAP7_75t_L g3330 ( 
.A(n_3149),
.B(n_637),
.C(n_634),
.D(n_635),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3051),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3145),
.B(n_637),
.Y(n_3332)
);

AOI322xp5_ASAP7_75t_L g3333 ( 
.A1(n_3065),
.A2(n_638),
.A3(n_639),
.B1(n_640),
.B2(n_641),
.C1(n_642),
.C2(n_643),
.Y(n_3333)
);

OAI221xp5_ASAP7_75t_L g3334 ( 
.A1(n_3062),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.C(n_641),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3287),
.A2(n_644),
.B(n_645),
.Y(n_3335)
);

NAND3xp33_ASAP7_75t_SL g3336 ( 
.A(n_3173),
.B(n_644),
.C(n_645),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_3189),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3276),
.B(n_646),
.Y(n_3338)
);

AND2x2_ASAP7_75t_L g3339 ( 
.A(n_3185),
.B(n_647),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3301),
.B(n_648),
.Y(n_3340)
);

NOR2x1_ASAP7_75t_L g3341 ( 
.A(n_3183),
.B(n_648),
.Y(n_3341)
);

NAND4xp25_ASAP7_75t_L g3342 ( 
.A(n_3322),
.B(n_651),
.C(n_649),
.D(n_650),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3177),
.A2(n_651),
.B(n_652),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3168),
.B(n_3284),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3194),
.B(n_3246),
.Y(n_3345)
);

NOR3xp33_ASAP7_75t_L g3346 ( 
.A(n_3179),
.B(n_653),
.C(n_654),
.Y(n_3346)
);

OAI221xp5_ASAP7_75t_L g3347 ( 
.A1(n_3294),
.A2(n_656),
.B1(n_654),
.B2(n_655),
.C(n_657),
.Y(n_3347)
);

OAI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3289),
.A2(n_656),
.B(n_657),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3167),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3256),
.B(n_658),
.Y(n_3350)
);

NOR3x1_ASAP7_75t_L g3351 ( 
.A(n_3314),
.B(n_658),
.C(n_659),
.Y(n_3351)
);

OAI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3204),
.A2(n_662),
.B1(n_660),
.B2(n_661),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3215),
.B(n_660),
.Y(n_3353)
);

NAND2xp33_ASAP7_75t_L g3354 ( 
.A(n_3171),
.B(n_662),
.Y(n_3354)
);

AND4x1_ASAP7_75t_L g3355 ( 
.A(n_3328),
.B(n_665),
.C(n_663),
.D(n_664),
.Y(n_3355)
);

NOR3xp33_ASAP7_75t_L g3356 ( 
.A(n_3317),
.B(n_3299),
.C(n_3176),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3304),
.A2(n_664),
.B(n_665),
.Y(n_3357)
);

AOI21xp5_ASAP7_75t_L g3358 ( 
.A1(n_3188),
.A2(n_666),
.B(n_667),
.Y(n_3358)
);

NAND3xp33_ASAP7_75t_L g3359 ( 
.A(n_3277),
.B(n_3308),
.C(n_3298),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3175),
.Y(n_3360)
);

NAND4xp25_ASAP7_75t_L g3361 ( 
.A(n_3259),
.B(n_669),
.C(n_666),
.D(n_668),
.Y(n_3361)
);

NAND3xp33_ASAP7_75t_L g3362 ( 
.A(n_3309),
.B(n_668),
.C(n_670),
.Y(n_3362)
);

AOI211xp5_ASAP7_75t_L g3363 ( 
.A1(n_3300),
.A2(n_672),
.B(n_670),
.C(n_671),
.Y(n_3363)
);

NOR3x1_ASAP7_75t_L g3364 ( 
.A(n_3174),
.B(n_671),
.C(n_673),
.Y(n_3364)
);

NAND4xp25_ASAP7_75t_L g3365 ( 
.A(n_3172),
.B(n_675),
.C(n_673),
.D(n_674),
.Y(n_3365)
);

INVxp67_ASAP7_75t_L g3366 ( 
.A(n_3245),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3162),
.B(n_676),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3205),
.Y(n_3368)
);

XNOR2xp5_ASAP7_75t_L g3369 ( 
.A(n_3288),
.B(n_676),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3313),
.B(n_677),
.Y(n_3370)
);

O2A1O1Ixp33_ASAP7_75t_L g3371 ( 
.A1(n_3305),
.A2(n_3201),
.B(n_3187),
.C(n_3334),
.Y(n_3371)
);

NOR3xp33_ASAP7_75t_L g3372 ( 
.A(n_3190),
.B(n_3320),
.C(n_3319),
.Y(n_3372)
);

NOR3xp33_ASAP7_75t_L g3373 ( 
.A(n_3325),
.B(n_3292),
.C(n_3290),
.Y(n_3373)
);

NAND3xp33_ASAP7_75t_L g3374 ( 
.A(n_3295),
.B(n_678),
.C(n_679),
.Y(n_3374)
);

AOI22xp5_ASAP7_75t_L g3375 ( 
.A1(n_3306),
.A2(n_681),
.B1(n_678),
.B2(n_680),
.Y(n_3375)
);

NOR3xp33_ASAP7_75t_L g3376 ( 
.A(n_3315),
.B(n_681),
.C(n_682),
.Y(n_3376)
);

OAI211xp5_ASAP7_75t_SL g3377 ( 
.A1(n_3169),
.A2(n_684),
.B(n_682),
.C(n_683),
.Y(n_3377)
);

NOR4xp25_ASAP7_75t_L g3378 ( 
.A(n_3330),
.B(n_685),
.C(n_683),
.D(n_684),
.Y(n_3378)
);

NOR3x1_ASAP7_75t_L g3379 ( 
.A(n_3327),
.B(n_685),
.C(n_686),
.Y(n_3379)
);

AOI211xp5_ASAP7_75t_L g3380 ( 
.A1(n_3310),
.A2(n_688),
.B(n_686),
.C(n_687),
.Y(n_3380)
);

AOI221xp5_ASAP7_75t_L g3381 ( 
.A1(n_3170),
.A2(n_689),
.B1(n_687),
.B2(n_688),
.C(n_690),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3209),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3311),
.B(n_3273),
.Y(n_3383)
);

AOI221xp5_ASAP7_75t_L g3384 ( 
.A1(n_3216),
.A2(n_692),
.B1(n_690),
.B2(n_691),
.C(n_693),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3207),
.Y(n_3385)
);

NAND4xp25_ASAP7_75t_L g3386 ( 
.A(n_3163),
.B(n_3225),
.C(n_3208),
.D(n_3191),
.Y(n_3386)
);

NAND3xp33_ASAP7_75t_L g3387 ( 
.A(n_3192),
.B(n_3166),
.C(n_3233),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3253),
.Y(n_3388)
);

NAND4xp25_ASAP7_75t_L g3389 ( 
.A(n_3296),
.B(n_695),
.C(n_691),
.D(n_694),
.Y(n_3389)
);

NAND4xp25_ASAP7_75t_L g3390 ( 
.A(n_3333),
.B(n_697),
.C(n_695),
.D(n_696),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_L g3391 ( 
.A(n_3195),
.B(n_696),
.Y(n_3391)
);

NOR4xp25_ASAP7_75t_L g3392 ( 
.A(n_3193),
.B(n_699),
.C(n_697),
.D(n_698),
.Y(n_3392)
);

NOR3xp33_ASAP7_75t_L g3393 ( 
.A(n_3231),
.B(n_700),
.C(n_701),
.Y(n_3393)
);

NOR2x1_ASAP7_75t_L g3394 ( 
.A(n_3260),
.B(n_894),
.Y(n_3394)
);

OAI211xp5_ASAP7_75t_SL g3395 ( 
.A1(n_3293),
.A2(n_703),
.B(n_701),
.C(n_702),
.Y(n_3395)
);

NAND4xp25_ASAP7_75t_L g3396 ( 
.A(n_3220),
.B(n_705),
.C(n_703),
.D(n_704),
.Y(n_3396)
);

AOI21xp33_ASAP7_75t_L g3397 ( 
.A1(n_3230),
.A2(n_704),
.B(n_705),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3235),
.B(n_706),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3202),
.B(n_706),
.Y(n_3399)
);

INVxp67_ASAP7_75t_SL g3400 ( 
.A(n_3272),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3263),
.B(n_707),
.Y(n_3401)
);

AOI211xp5_ASAP7_75t_L g3402 ( 
.A1(n_3180),
.A2(n_709),
.B(n_707),
.C(n_708),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3165),
.B(n_708),
.Y(n_3403)
);

OAI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3243),
.A2(n_3186),
.B(n_3198),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3255),
.B(n_3281),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_SL g3406 ( 
.A(n_3241),
.B(n_709),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3283),
.Y(n_3407)
);

AND3x1_ASAP7_75t_L g3408 ( 
.A(n_3324),
.B(n_892),
.C(n_710),
.Y(n_3408)
);

O2A1O1Ixp33_ASAP7_75t_L g3409 ( 
.A1(n_3275),
.A2(n_712),
.B(n_710),
.C(n_711),
.Y(n_3409)
);

NAND4xp75_ASAP7_75t_L g3410 ( 
.A(n_3227),
.B(n_715),
.C(n_713),
.D(n_714),
.Y(n_3410)
);

OAI21xp33_ASAP7_75t_L g3411 ( 
.A1(n_3326),
.A2(n_713),
.B(n_714),
.Y(n_3411)
);

NAND3xp33_ASAP7_75t_L g3412 ( 
.A(n_3254),
.B(n_715),
.C(n_716),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3318),
.B(n_716),
.Y(n_3413)
);

OAI211xp5_ASAP7_75t_L g3414 ( 
.A1(n_3252),
.A2(n_719),
.B(n_717),
.C(n_718),
.Y(n_3414)
);

NAND3xp33_ASAP7_75t_L g3415 ( 
.A(n_3258),
.B(n_718),
.C(n_719),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3199),
.A2(n_722),
.B1(n_720),
.B2(n_721),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3291),
.B(n_723),
.Y(n_3417)
);

AOI221xp5_ASAP7_75t_L g3418 ( 
.A1(n_3279),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.C(n_726),
.Y(n_3418)
);

OA211x2_ASAP7_75t_L g3419 ( 
.A1(n_3219),
.A2(n_728),
.B(n_725),
.C(n_727),
.Y(n_3419)
);

NOR2x1_ASAP7_75t_L g3420 ( 
.A(n_3268),
.B(n_728),
.Y(n_3420)
);

NOR3xp33_ASAP7_75t_L g3421 ( 
.A(n_3210),
.B(n_729),
.C(n_731),
.Y(n_3421)
);

NOR2x1_ASAP7_75t_L g3422 ( 
.A(n_3280),
.B(n_729),
.Y(n_3422)
);

NOR4xp25_ASAP7_75t_L g3423 ( 
.A(n_3213),
.B(n_735),
.C(n_733),
.D(n_734),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3329),
.Y(n_3424)
);

NOR4xp25_ASAP7_75t_L g3425 ( 
.A(n_3237),
.B(n_735),
.C(n_733),
.D(n_734),
.Y(n_3425)
);

NAND4xp25_ASAP7_75t_L g3426 ( 
.A(n_3228),
.B(n_738),
.C(n_736),
.D(n_737),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3312),
.B(n_736),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3321),
.B(n_737),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3178),
.B(n_738),
.Y(n_3429)
);

NAND4xp25_ASAP7_75t_L g3430 ( 
.A(n_3206),
.B(n_3197),
.C(n_3214),
.D(n_3196),
.Y(n_3430)
);

NAND3xp33_ASAP7_75t_L g3431 ( 
.A(n_3232),
.B(n_739),
.C(n_740),
.Y(n_3431)
);

NOR3xp33_ASAP7_75t_L g3432 ( 
.A(n_3211),
.B(n_739),
.C(n_741),
.Y(n_3432)
);

OAI211xp5_ASAP7_75t_L g3433 ( 
.A1(n_3278),
.A2(n_743),
.B(n_741),
.C(n_742),
.Y(n_3433)
);

NOR2x1p5_ASAP7_75t_SL g3434 ( 
.A(n_3331),
.B(n_742),
.Y(n_3434)
);

AOI221xp5_ASAP7_75t_L g3435 ( 
.A1(n_3302),
.A2(n_746),
.B1(n_744),
.B2(n_745),
.C(n_747),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3264),
.B(n_744),
.Y(n_3436)
);

O2A1O1Ixp33_ASAP7_75t_L g3437 ( 
.A1(n_3223),
.A2(n_748),
.B(n_746),
.C(n_747),
.Y(n_3437)
);

OAI21xp5_ASAP7_75t_SL g3438 ( 
.A1(n_3282),
.A2(n_748),
.B(n_749),
.Y(n_3438)
);

NAND3x1_ASAP7_75t_L g3439 ( 
.A(n_3286),
.B(n_889),
.C(n_749),
.Y(n_3439)
);

AOI22x1_ASAP7_75t_L g3440 ( 
.A1(n_3221),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_L g3441 ( 
.A(n_3307),
.B(n_750),
.Y(n_3441)
);

NAND2xp33_ASAP7_75t_L g3442 ( 
.A(n_3297),
.B(n_753),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3316),
.B(n_754),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_3332),
.B(n_3262),
.Y(n_3444)
);

NOR3xp33_ASAP7_75t_L g3445 ( 
.A(n_3222),
.B(n_755),
.C(n_756),
.Y(n_3445)
);

NAND3xp33_ASAP7_75t_L g3446 ( 
.A(n_3164),
.B(n_756),
.C(n_757),
.Y(n_3446)
);

CKINVDCx16_ASAP7_75t_R g3447 ( 
.A(n_3285),
.Y(n_3447)
);

NAND3xp33_ASAP7_75t_L g3448 ( 
.A(n_3303),
.B(n_758),
.C(n_759),
.Y(n_3448)
);

AOI211xp5_ASAP7_75t_L g3449 ( 
.A1(n_3239),
.A2(n_761),
.B(n_759),
.C(n_760),
.Y(n_3449)
);

NAND3xp33_ASAP7_75t_L g3450 ( 
.A(n_3323),
.B(n_760),
.C(n_761),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3265),
.B(n_762),
.Y(n_3451)
);

A2O1A1Ixp33_ASAP7_75t_L g3452 ( 
.A1(n_3181),
.A2(n_3182),
.B(n_3247),
.C(n_3184),
.Y(n_3452)
);

OAI211xp5_ASAP7_75t_SL g3453 ( 
.A1(n_3236),
.A2(n_3217),
.B(n_3229),
.C(n_3261),
.Y(n_3453)
);

NOR4xp25_ASAP7_75t_L g3454 ( 
.A(n_3224),
.B(n_3218),
.C(n_3244),
.D(n_3234),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_SL g3455 ( 
.A(n_3271),
.B(n_762),
.Y(n_3455)
);

NAND4xp75_ASAP7_75t_L g3456 ( 
.A(n_3200),
.B(n_765),
.C(n_763),
.D(n_764),
.Y(n_3456)
);

AOI21xp33_ASAP7_75t_L g3457 ( 
.A1(n_3242),
.A2(n_763),
.B(n_764),
.Y(n_3457)
);

NOR3xp33_ASAP7_75t_L g3458 ( 
.A(n_3226),
.B(n_766),
.C(n_767),
.Y(n_3458)
);

AOI211xp5_ASAP7_75t_L g3459 ( 
.A1(n_3203),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3274),
.B(n_768),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_3212),
.B(n_769),
.Y(n_3461)
);

NAND3xp33_ASAP7_75t_L g3462 ( 
.A(n_3380),
.B(n_3248),
.C(n_3250),
.Y(n_3462)
);

INVxp67_ASAP7_75t_L g3463 ( 
.A(n_3337),
.Y(n_3463)
);

NOR3xp33_ASAP7_75t_L g3464 ( 
.A(n_3447),
.B(n_3257),
.C(n_3240),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_3366),
.B(n_3238),
.Y(n_3465)
);

O2A1O1Ixp33_ASAP7_75t_L g3466 ( 
.A1(n_3383),
.A2(n_3270),
.B(n_3269),
.C(n_3249),
.Y(n_3466)
);

NOR2x1_ASAP7_75t_L g3467 ( 
.A(n_3341),
.B(n_3267),
.Y(n_3467)
);

OAI211xp5_ASAP7_75t_L g3468 ( 
.A1(n_3361),
.A2(n_3378),
.B(n_3392),
.C(n_3342),
.Y(n_3468)
);

HB1xp67_ASAP7_75t_L g3469 ( 
.A(n_3345),
.Y(n_3469)
);

NOR3xp33_ASAP7_75t_L g3470 ( 
.A(n_3397),
.B(n_3266),
.C(n_3251),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3349),
.Y(n_3471)
);

NAND4xp25_ASAP7_75t_L g3472 ( 
.A(n_3344),
.B(n_771),
.C(n_769),
.D(n_770),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3400),
.B(n_770),
.Y(n_3473)
);

NOR3xp33_ASAP7_75t_L g3474 ( 
.A(n_3347),
.B(n_771),
.C(n_772),
.Y(n_3474)
);

NOR2x1p5_ASAP7_75t_L g3475 ( 
.A(n_3396),
.B(n_772),
.Y(n_3475)
);

NOR2x1_ASAP7_75t_L g3476 ( 
.A(n_3394),
.B(n_3340),
.Y(n_3476)
);

NOR3xp33_ASAP7_75t_L g3477 ( 
.A(n_3426),
.B(n_773),
.C(n_774),
.Y(n_3477)
);

NOR2x1_ASAP7_75t_L g3478 ( 
.A(n_3455),
.B(n_773),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3444),
.B(n_3356),
.Y(n_3479)
);

NOR3xp33_ASAP7_75t_L g3480 ( 
.A(n_3387),
.B(n_775),
.C(n_776),
.Y(n_3480)
);

NOR2x1_ASAP7_75t_L g3481 ( 
.A(n_3422),
.B(n_775),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3404),
.B(n_776),
.Y(n_3482)
);

NOR2x1_ASAP7_75t_L g3483 ( 
.A(n_3429),
.B(n_777),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3360),
.Y(n_3484)
);

NOR2x1_ASAP7_75t_L g3485 ( 
.A(n_3420),
.B(n_777),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_3386),
.B(n_778),
.Y(n_3486)
);

NOR3xp33_ASAP7_75t_SL g3487 ( 
.A(n_3336),
.B(n_778),
.C(n_779),
.Y(n_3487)
);

NOR2xp33_ASAP7_75t_L g3488 ( 
.A(n_3350),
.B(n_779),
.Y(n_3488)
);

NOR2x1p5_ASAP7_75t_L g3489 ( 
.A(n_3374),
.B(n_780),
.Y(n_3489)
);

A2O1A1Ixp33_ASAP7_75t_L g3490 ( 
.A1(n_3371),
.A2(n_783),
.B(n_781),
.C(n_782),
.Y(n_3490)
);

OAI211xp5_ASAP7_75t_L g3491 ( 
.A1(n_3423),
.A2(n_3335),
.B(n_3454),
.C(n_3390),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_3339),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3358),
.A2(n_781),
.B(n_782),
.Y(n_3493)
);

NOR2x1_ASAP7_75t_L g3494 ( 
.A(n_3412),
.B(n_783),
.Y(n_3494)
);

NOR2x1_ASAP7_75t_L g3495 ( 
.A(n_3415),
.B(n_784),
.Y(n_3495)
);

AND2x4_ASAP7_75t_L g3496 ( 
.A(n_3405),
.B(n_785),
.Y(n_3496)
);

O2A1O1Ixp33_ASAP7_75t_L g3497 ( 
.A1(n_3398),
.A2(n_787),
.B(n_785),
.C(n_786),
.Y(n_3497)
);

NAND4xp75_ASAP7_75t_L g3498 ( 
.A(n_3351),
.B(n_788),
.C(n_786),
.D(n_787),
.Y(n_3498)
);

NAND4xp25_ASAP7_75t_L g3499 ( 
.A(n_3373),
.B(n_791),
.C(n_789),
.D(n_790),
.Y(n_3499)
);

AOI21xp5_ASAP7_75t_L g3500 ( 
.A1(n_3343),
.A2(n_791),
.B(n_792),
.Y(n_3500)
);

AOI211x1_ASAP7_75t_L g3501 ( 
.A1(n_3359),
.A2(n_794),
.B(n_792),
.C(n_793),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3425),
.B(n_3372),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3439),
.B(n_793),
.Y(n_3503)
);

NAND3xp33_ASAP7_75t_SL g3504 ( 
.A(n_3376),
.B(n_794),
.C(n_795),
.Y(n_3504)
);

NOR2xp67_ASAP7_75t_L g3505 ( 
.A(n_3382),
.B(n_795),
.Y(n_3505)
);

NOR2x1_ASAP7_75t_L g3506 ( 
.A(n_3338),
.B(n_796),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3368),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3385),
.Y(n_3508)
);

AOI211x1_ASAP7_75t_SL g3509 ( 
.A1(n_3453),
.A2(n_798),
.B(n_796),
.C(n_797),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_3354),
.A2(n_797),
.B(n_798),
.Y(n_3510)
);

NOR2x1_ASAP7_75t_L g3511 ( 
.A(n_3401),
.B(n_799),
.Y(n_3511)
);

NOR2x1_ASAP7_75t_L g3512 ( 
.A(n_3431),
.B(n_799),
.Y(n_3512)
);

NOR2x1_ASAP7_75t_L g3513 ( 
.A(n_3362),
.B(n_800),
.Y(n_3513)
);

NAND4xp75_ASAP7_75t_L g3514 ( 
.A(n_3364),
.B(n_802),
.C(n_800),
.D(n_801),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3353),
.B(n_802),
.Y(n_3515)
);

NAND4xp25_ASAP7_75t_L g3516 ( 
.A(n_3430),
.B(n_805),
.C(n_803),
.D(n_804),
.Y(n_3516)
);

NOR2x1_ASAP7_75t_L g3517 ( 
.A(n_3446),
.B(n_803),
.Y(n_3517)
);

NAND3x2_ASAP7_75t_L g3518 ( 
.A(n_3355),
.B(n_806),
.C(n_807),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3413),
.B(n_806),
.Y(n_3519)
);

NOR3xp33_ASAP7_75t_SL g3520 ( 
.A(n_3389),
.B(n_807),
.C(n_808),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_L g3521 ( 
.A1(n_3393),
.A2(n_887),
.B1(n_810),
.B2(n_808),
.Y(n_3521)
);

NOR3xp33_ASAP7_75t_SL g3522 ( 
.A(n_3414),
.B(n_809),
.C(n_811),
.Y(n_3522)
);

NOR3xp33_ASAP7_75t_L g3523 ( 
.A(n_3457),
.B(n_809),
.C(n_811),
.Y(n_3523)
);

INVxp67_ASAP7_75t_SL g3524 ( 
.A(n_3379),
.Y(n_3524)
);

NOR2xp67_ASAP7_75t_L g3525 ( 
.A(n_3388),
.B(n_812),
.Y(n_3525)
);

NAND2x1p5_ASAP7_75t_L g3526 ( 
.A(n_3481),
.B(n_3406),
.Y(n_3526)
);

OR3x2_ASAP7_75t_L g3527 ( 
.A(n_3516),
.B(n_3365),
.C(n_3407),
.Y(n_3527)
);

NOR3xp33_ASAP7_75t_L g3528 ( 
.A(n_3479),
.B(n_3384),
.C(n_3433),
.Y(n_3528)
);

NOR3xp33_ASAP7_75t_SL g3529 ( 
.A(n_3491),
.B(n_3438),
.C(n_3377),
.Y(n_3529)
);

NOR2x1p5_ASAP7_75t_L g3530 ( 
.A(n_3524),
.B(n_3456),
.Y(n_3530)
);

INVxp67_ASAP7_75t_SL g3531 ( 
.A(n_3505),
.Y(n_3531)
);

CKINVDCx6p67_ASAP7_75t_R g3532 ( 
.A(n_3492),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_3463),
.B(n_3443),
.Y(n_3533)
);

AND3x4_ASAP7_75t_L g3534 ( 
.A(n_3464),
.B(n_3421),
.C(n_3346),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3469),
.B(n_3424),
.Y(n_3535)
);

NAND4xp75_ASAP7_75t_L g3536 ( 
.A(n_3476),
.B(n_3419),
.C(n_3348),
.D(n_3408),
.Y(n_3536)
);

INVxp67_ASAP7_75t_L g3537 ( 
.A(n_3483),
.Y(n_3537)
);

NAND3xp33_ASAP7_75t_L g3538 ( 
.A(n_3502),
.B(n_3459),
.C(n_3363),
.Y(n_3538)
);

NOR2xp67_ASAP7_75t_L g3539 ( 
.A(n_3492),
.B(n_3357),
.Y(n_3539)
);

NOR2xp67_ASAP7_75t_L g3540 ( 
.A(n_3492),
.B(n_3369),
.Y(n_3540)
);

NOR2x1_ASAP7_75t_L g3541 ( 
.A(n_3467),
.B(n_3448),
.Y(n_3541)
);

NAND4xp25_ASAP7_75t_L g3542 ( 
.A(n_3468),
.B(n_3375),
.C(n_3402),
.D(n_3449),
.Y(n_3542)
);

NOR3x1_ASAP7_75t_L g3543 ( 
.A(n_3514),
.B(n_3352),
.C(n_3410),
.Y(n_3543)
);

OAI22xp5_ASAP7_75t_L g3544 ( 
.A1(n_3462),
.A2(n_3452),
.B1(n_3416),
.B2(n_3450),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3490),
.B(n_3367),
.Y(n_3545)
);

NOR3x2_ASAP7_75t_L g3546 ( 
.A(n_3498),
.B(n_3434),
.C(n_3442),
.Y(n_3546)
);

BUFx3_ASAP7_75t_L g3547 ( 
.A(n_3496),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3465),
.B(n_3515),
.Y(n_3548)
);

NOR3xp33_ASAP7_75t_L g3549 ( 
.A(n_3482),
.B(n_3370),
.C(n_3381),
.Y(n_3549)
);

INVx2_ASAP7_75t_SL g3550 ( 
.A(n_3496),
.Y(n_3550)
);

OR2x2_ASAP7_75t_L g3551 ( 
.A(n_3503),
.B(n_3399),
.Y(n_3551)
);

A2O1A1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_3497),
.A2(n_3437),
.B(n_3409),
.C(n_3432),
.Y(n_3552)
);

AND3x4_ASAP7_75t_L g3553 ( 
.A(n_3520),
.B(n_3445),
.C(n_3458),
.Y(n_3553)
);

NAND3xp33_ASAP7_75t_L g3554 ( 
.A(n_3522),
.B(n_3435),
.C(n_3418),
.Y(n_3554)
);

AOI211xp5_ASAP7_75t_L g3555 ( 
.A1(n_3466),
.A2(n_3395),
.B(n_3411),
.C(n_3461),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3485),
.B(n_3391),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3471),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3473),
.B(n_3436),
.Y(n_3558)
);

NOR2xp67_ASAP7_75t_L g3559 ( 
.A(n_3525),
.B(n_3451),
.Y(n_3559)
);

NOR2xp67_ASAP7_75t_L g3560 ( 
.A(n_3484),
.B(n_3460),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3480),
.B(n_3441),
.Y(n_3561)
);

NAND2x1p5_ASAP7_75t_L g3562 ( 
.A(n_3478),
.B(n_3440),
.Y(n_3562)
);

XNOR2xp5_ASAP7_75t_L g3563 ( 
.A(n_3546),
.B(n_3518),
.Y(n_3563)
);

INVx5_ASAP7_75t_L g3564 ( 
.A(n_3550),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3535),
.Y(n_3565)
);

OR2x2_ASAP7_75t_L g3566 ( 
.A(n_3551),
.B(n_3507),
.Y(n_3566)
);

NAND3x1_ASAP7_75t_L g3567 ( 
.A(n_3541),
.B(n_3506),
.C(n_3513),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3547),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3531),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3532),
.Y(n_3570)
);

OAI22xp5_ASAP7_75t_L g3571 ( 
.A1(n_3538),
.A2(n_3487),
.B1(n_3501),
.B2(n_3512),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3533),
.Y(n_3572)
);

NAND4xp75_ASAP7_75t_L g3573 ( 
.A(n_3543),
.B(n_3529),
.C(n_3540),
.D(n_3495),
.Y(n_3573)
);

O2A1O1Ixp33_ASAP7_75t_L g3574 ( 
.A1(n_3537),
.A2(n_3477),
.B(n_3504),
.C(n_3474),
.Y(n_3574)
);

AO22x2_ASAP7_75t_L g3575 ( 
.A1(n_3534),
.A2(n_3508),
.B1(n_3470),
.B2(n_3510),
.Y(n_3575)
);

HB1xp67_ASAP7_75t_L g3576 ( 
.A(n_3559),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3548),
.B(n_3511),
.Y(n_3577)
);

XNOR2xp5_ASAP7_75t_L g3578 ( 
.A(n_3553),
.B(n_3475),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3526),
.Y(n_3579)
);

INVx4_ASAP7_75t_L g3580 ( 
.A(n_3562),
.Y(n_3580)
);

AND3x4_ASAP7_75t_L g3581 ( 
.A(n_3528),
.B(n_3494),
.C(n_3517),
.Y(n_3581)
);

BUFx12f_ASAP7_75t_L g3582 ( 
.A(n_3530),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3557),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3564),
.Y(n_3584)
);

HB1xp67_ASAP7_75t_L g3585 ( 
.A(n_3564),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3569),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3581),
.A2(n_3536),
.B1(n_3554),
.B2(n_3552),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3576),
.Y(n_3588)
);

INVx1_ASAP7_75t_SL g3589 ( 
.A(n_3577),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3580),
.Y(n_3590)
);

AOI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3571),
.A2(n_3544),
.B1(n_3549),
.B2(n_3542),
.Y(n_3591)
);

OR2x6_ASAP7_75t_L g3592 ( 
.A(n_3570),
.B(n_3556),
.Y(n_3592)
);

AND3x1_ASAP7_75t_L g3593 ( 
.A(n_3574),
.B(n_3555),
.C(n_3558),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3573),
.A2(n_3545),
.B1(n_3527),
.B2(n_3539),
.Y(n_3594)
);

NOR3xp33_ASAP7_75t_L g3595 ( 
.A(n_3587),
.B(n_3568),
.C(n_3579),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3593),
.A2(n_3561),
.B(n_3575),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3584),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3585),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3592),
.A2(n_3563),
.B(n_3578),
.Y(n_3599)
);

OAI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_3591),
.A2(n_3567),
.B1(n_3582),
.B2(n_3521),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3588),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3586),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_L g3603 ( 
.A1(n_3590),
.A2(n_3572),
.B1(n_3565),
.B2(n_3560),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3589),
.B(n_3486),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3592),
.Y(n_3605)
);

NAND3xp33_ASAP7_75t_L g3606 ( 
.A(n_3596),
.B(n_3594),
.C(n_3583),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3597),
.Y(n_3607)
);

OAI22xp5_ASAP7_75t_L g3608 ( 
.A1(n_3605),
.A2(n_3489),
.B1(n_3566),
.B2(n_3500),
.Y(n_3608)
);

XNOR2x1_ASAP7_75t_L g3609 ( 
.A(n_3600),
.B(n_3604),
.Y(n_3609)
);

OAI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_3603),
.A2(n_3488),
.B1(n_3493),
.B2(n_3417),
.Y(n_3610)
);

OAI331xp33_ASAP7_75t_L g3611 ( 
.A1(n_3598),
.A2(n_3519),
.A3(n_3403),
.B1(n_3427),
.B2(n_3428),
.B3(n_3499),
.C1(n_3509),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3607),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3608),
.B(n_3599),
.Y(n_3613)
);

AOI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3611),
.A2(n_3595),
.B1(n_3601),
.B2(n_3523),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3614),
.A2(n_3606),
.B1(n_3609),
.B2(n_3610),
.Y(n_3615)
);

NAND2xp33_ASAP7_75t_L g3616 ( 
.A(n_3613),
.B(n_3602),
.Y(n_3616)
);

OR2x6_ASAP7_75t_L g3617 ( 
.A(n_3615),
.B(n_3612),
.Y(n_3617)
);

AOI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3617),
.A2(n_3616),
.B1(n_3472),
.B2(n_814),
.Y(n_3618)
);


endmodule