module fake_jpeg_26607_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_18),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_30),
.Y(n_89)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_25),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_24),
.C(n_20),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_51),
.C(n_35),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_39),
.B1(n_21),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_42),
.B(n_39),
.C(n_24),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_72),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_80),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_36),
.B(n_41),
.C(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_35),
.B1(n_55),
.B2(n_45),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_25),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_27),
.B1(n_31),
.B2(n_18),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_88),
.Y(n_99)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_32),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_41),
.B1(n_27),
.B2(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_32),
.B1(n_23),
.B2(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_16),
.B(n_30),
.C(n_4),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_15),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_46),
.B1(n_58),
.B2(n_30),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_46),
.B1(n_16),
.B2(n_30),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_15),
.C(n_14),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_12),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_5),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_76),
.B1(n_67),
.B2(n_66),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_137),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_91),
.B(n_89),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_104),
.B(n_9),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_71),
.B(n_65),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_143),
.B(n_139),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_7),
.B1(n_9),
.B2(n_136),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_113),
.B(n_110),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_111),
.B(n_108),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_138),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_94),
.B1(n_93),
.B2(n_83),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_104),
.B1(n_69),
.B2(n_11),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_83),
.Y(n_137)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_66),
.A3(n_79),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_144),
.B(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_96),
.A2(n_69),
.B1(n_75),
.B2(n_11),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_150),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_109),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_148),
.B(n_153),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_121),
.B1(n_120),
.B2(n_107),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_122),
.B1(n_134),
.B2(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_103),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_163),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_157),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_123),
.B(n_124),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_174),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_153),
.B(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_179),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_171),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_165),
.B1(n_164),
.B2(n_159),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_127),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_161),
.C(n_126),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_133),
.B(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_157),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_193),
.B(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_125),
.B1(n_166),
.B2(n_162),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_161),
.B1(n_149),
.B2(n_158),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_170),
.B(n_177),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_202),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_204),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_126),
.C(n_180),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_183),
.Y(n_208)
);

XOR2x2_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_173),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_129),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_182),
.C(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_211),
.C(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_215),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_184),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_185),
.C(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_191),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_198),
.B1(n_200),
.B2(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_200),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_213),
.B(n_194),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_214),
.C(n_187),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_218),
.A3(n_129),
.B1(n_133),
.B2(n_138),
.C1(n_142),
.C2(n_9),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_138),
.B(n_7),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_223),
.Y(n_226)
);


endmodule