module real_aes_9863_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_1499;
wire n_700;
wire n_399;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_1779;
wire n_473;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_1772;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1323;
wire n_1280;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1142 ( .A(n_0), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_1), .A2(n_152), .B1(n_363), .B2(n_374), .C(n_381), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_1), .A2(n_325), .B1(n_505), .B2(n_508), .C(n_512), .Y(n_504) );
OA22x2_ASAP7_75t_L g1333 ( .A1(n_2), .A2(n_1334), .B1(n_1385), .B2(n_1386), .Y(n_1333) );
INVxp67_ASAP7_75t_SL g1386 ( .A(n_2), .Y(n_1386) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_3), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_4), .Y(n_1029) );
INVx1_ASAP7_75t_L g1517 ( .A(n_5), .Y(n_1517) );
OAI221xp5_ASAP7_75t_L g1130 ( .A1(n_6), .A2(n_293), .B1(n_407), .B2(n_567), .C(n_965), .Y(n_1130) );
OAI22xp33_ASAP7_75t_SL g1152 ( .A1(n_6), .A2(n_293), .B1(n_828), .B2(n_830), .Y(n_1152) );
INVxp33_ASAP7_75t_L g1126 ( .A(n_7), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1147 ( .A1(n_7), .A2(n_82), .B1(n_535), .B2(n_824), .C(n_1148), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_8), .A2(n_79), .B1(n_824), .B2(n_1017), .C(n_1019), .Y(n_1016) );
INVx1_ASAP7_75t_L g1036 ( .A(n_8), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_9), .A2(n_141), .B1(n_902), .B2(n_904), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_9), .A2(n_49), .B1(n_820), .B2(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g1140 ( .A(n_10), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_11), .A2(n_245), .B1(n_713), .B2(n_715), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g773 ( .A(n_11), .Y(n_773) );
INVx1_ASAP7_75t_L g1188 ( .A(n_12), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1237 ( .A1(n_13), .A2(n_54), .B1(n_1238), .B2(n_1240), .Y(n_1237) );
INVx1_ASAP7_75t_L g1262 ( .A(n_13), .Y(n_1262) );
XNOR2x2_ASAP7_75t_L g894 ( .A(n_14), .B(n_895), .Y(n_894) );
AO221x2_ASAP7_75t_L g1515 ( .A1(n_14), .A2(n_242), .B1(n_1479), .B2(n_1514), .C(n_1516), .Y(n_1515) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_15), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_16), .A2(n_49), .B1(n_907), .B2(n_908), .Y(n_906) );
AOI21xp33_ASAP7_75t_L g936 ( .A1(n_16), .A2(n_531), .B(n_937), .Y(n_936) );
CKINVDCx16_ASAP7_75t_R g1537 ( .A(n_17), .Y(n_1537) );
OAI22xp5_ASAP7_75t_L g1336 ( .A1(n_18), .A2(n_218), .B1(n_1193), .B2(n_1337), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_18), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1441 ( .A(n_19), .Y(n_1441) );
INVxp67_ASAP7_75t_L g572 ( .A(n_20), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_20), .A2(n_51), .B1(n_614), .B2(n_615), .C(n_616), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_21), .A2(n_271), .B1(n_843), .B2(n_1173), .Y(n_1177) );
INVxp67_ASAP7_75t_SL g1213 ( .A(n_21), .Y(n_1213) );
OAI221xp5_ASAP7_75t_L g1738 ( .A1(n_22), .A2(n_58), .B1(n_1739), .B2(n_1740), .C(n_1741), .Y(n_1738) );
INVx1_ASAP7_75t_L g1765 ( .A(n_22), .Y(n_1765) );
INVx1_ASAP7_75t_L g924 ( .A(n_23), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_23), .A2(n_276), .B1(n_934), .B2(n_937), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_24), .A2(n_318), .B1(n_859), .B2(n_1220), .C(n_1222), .Y(n_1219) );
INVx1_ASAP7_75t_L g1250 ( .A(n_24), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_25), .A2(n_312), .B1(n_667), .B2(n_1070), .Y(n_1287) );
INVxp67_ASAP7_75t_SL g1327 ( .A(n_25), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_26), .A2(n_327), .B1(n_609), .B2(n_668), .Y(n_711) );
INVx1_ASAP7_75t_L g745 ( .A(n_26), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_27), .A2(n_110), .B1(n_567), .B2(n_568), .C(n_569), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_27), .A2(n_110), .B1(n_609), .B2(n_610), .Y(n_608) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_28), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_28), .A2(n_305), .B1(n_505), .B2(n_616), .C(n_814), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_29), .A2(n_208), .B1(n_615), .B2(n_616), .C(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1048 ( .A(n_29), .Y(n_1048) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_30), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g1170 ( .A1(n_31), .A2(n_550), .B(n_1171), .C(n_1180), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g1207 ( .A1(n_31), .A2(n_173), .B1(n_908), .B2(n_1208), .C(n_1210), .Y(n_1207) );
INVx1_ASAP7_75t_L g1753 ( .A(n_32), .Y(n_1753) );
INVx1_ASAP7_75t_L g335 ( .A(n_33), .Y(n_335) );
INVx1_ASAP7_75t_L g724 ( .A(n_34), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_34), .A2(n_289), .B1(n_763), .B2(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g632 ( .A(n_35), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_35), .A2(n_164), .B1(n_671), .B2(n_673), .C(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g1389 ( .A(n_36), .Y(n_1389) );
OAI221xp5_ASAP7_75t_L g1341 ( .A1(n_37), .A2(n_59), .B1(n_396), .B2(n_406), .C(n_965), .Y(n_1341) );
OAI222xp33_ASAP7_75t_L g1368 ( .A1(n_37), .A2(n_59), .B1(n_203), .B2(n_487), .C1(n_492), .C2(n_861), .Y(n_1368) );
AOI21xp33_ASAP7_75t_L g1448 ( .A1(n_38), .A2(n_687), .B(n_1449), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1469 ( .A1(n_38), .A2(n_73), .B1(n_365), .B2(n_423), .C(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1292 ( .A(n_39), .Y(n_1292) );
OAI221xp5_ASAP7_75t_L g1310 ( .A1(n_39), .A2(n_272), .B1(n_363), .B2(n_1311), .C(n_1312), .Y(n_1310) );
AOI22xp33_ASAP7_75t_SL g1172 ( .A1(n_40), .A2(n_89), .B1(n_619), .B2(n_1173), .Y(n_1172) );
AOI22xp33_ASAP7_75t_SL g1195 ( .A1(n_40), .A2(n_159), .B1(n_758), .B2(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g735 ( .A(n_41), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_41), .A2(n_298), .B1(n_758), .B2(n_760), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_42), .A2(n_179), .B1(n_603), .B2(n_619), .C(n_1179), .Y(n_1178) );
OAI21xp33_ASAP7_75t_SL g1192 ( .A1(n_42), .A2(n_1193), .B(n_1194), .Y(n_1192) );
OAI222xp33_ASAP7_75t_L g853 ( .A1(n_43), .A2(n_156), .B1(n_251), .B2(n_854), .C1(n_856), .C2(n_858), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g888 ( .A1(n_43), .A2(n_156), .B1(n_889), .B2(n_891), .C(n_892), .Y(n_888) );
CKINVDCx16_ASAP7_75t_R g1278 ( .A(n_44), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_45), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g1234 ( .A(n_46), .Y(n_1234) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_47), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_47), .A2(n_192), .B1(n_606), .B2(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_48), .A2(n_97), .B1(n_396), .B2(n_405), .C(n_410), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g486 ( .A1(n_48), .A2(n_97), .B1(n_487), .B2(n_492), .C(n_497), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g1350 ( .A(n_50), .Y(n_1350) );
INVxp33_ASAP7_75t_L g583 ( .A(n_51), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g1398 ( .A1(n_52), .A2(n_80), .B1(n_505), .B2(n_616), .C(n_713), .Y(n_1398) );
INVxp67_ASAP7_75t_L g1426 ( .A(n_52), .Y(n_1426) );
INVxp67_ASAP7_75t_L g953 ( .A(n_53), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1543 ( .A1(n_53), .A2(n_299), .B1(n_1479), .B2(n_1514), .Y(n_1543) );
INVx1_ASAP7_75t_L g1264 ( .A(n_54), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_55), .A2(n_186), .B1(n_534), .B2(n_1159), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_55), .A2(n_186), .B1(n_763), .B2(n_1196), .Y(n_1319) );
OAI221xp5_ASAP7_75t_L g1442 ( .A1(n_56), .A2(n_128), .B1(n_1228), .B2(n_1443), .C(n_1444), .Y(n_1442) );
INVx1_ASAP7_75t_L g1473 ( .A(n_56), .Y(n_1473) );
INVxp67_ASAP7_75t_L g977 ( .A(n_57), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_57), .A2(n_86), .B1(n_823), .B2(n_1002), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1762 ( .A1(n_58), .A2(n_187), .B1(n_880), .B2(n_1763), .C(n_1764), .Y(n_1762) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_60), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g1348 ( .A(n_61), .Y(n_1348) );
AOI21xp33_ASAP7_75t_L g1076 ( .A1(n_62), .A2(n_603), .B(n_720), .Y(n_1076) );
INVxp33_ASAP7_75t_L g1098 ( .A(n_62), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_63), .A2(n_193), .B1(n_830), .B2(n_997), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_63), .A2(n_193), .B1(n_406), .B2(n_569), .C(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1402 ( .A(n_64), .Y(n_1402) );
INVx1_ASAP7_75t_L g982 ( .A(n_65), .Y(n_982) );
AOI22x1_ASAP7_75t_L g1167 ( .A1(n_66), .A2(n_1168), .B1(n_1214), .B2(n_1215), .Y(n_1167) );
INVxp67_ASAP7_75t_L g1214 ( .A(n_66), .Y(n_1214) );
XNOR2x2_ASAP7_75t_L g1216 ( .A(n_67), .B(n_1217), .Y(n_1216) );
INVxp33_ASAP7_75t_L g1125 ( .A(n_68), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_68), .A2(n_254), .B1(n_726), .B2(n_1151), .Y(n_1150) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_69), .Y(n_1068) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_70), .Y(n_921) );
INVxp33_ASAP7_75t_L g565 ( .A(n_71), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_71), .A2(n_328), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_72), .A2(n_160), .B1(n_423), .B2(n_911), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_72), .A2(n_160), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1447 ( .A1(n_73), .A2(n_211), .B1(n_693), .B2(n_934), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g1751 ( .A1(n_74), .A2(n_161), .B1(n_715), .B2(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1772 ( .A(n_74), .Y(n_1772) );
INVxp33_ASAP7_75t_SL g1307 ( .A(n_75), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_75), .A2(n_310), .B1(n_1196), .B2(n_1321), .Y(n_1323) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_76), .A2(n_144), .B1(n_396), .B2(n_568), .C(n_635), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_76), .A2(n_144), .B1(n_667), .B2(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g831 ( .A(n_77), .Y(n_831) );
INVx1_ASAP7_75t_L g371 ( .A(n_78), .Y(n_371) );
OR2x2_ASAP7_75t_L g403 ( .A(n_78), .B(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g416 ( .A(n_78), .Y(n_416) );
BUFx2_ASAP7_75t_L g464 ( .A(n_78), .Y(n_464) );
INVx1_ASAP7_75t_L g1038 ( .A(n_79), .Y(n_1038) );
INVxp33_ASAP7_75t_SL g1424 ( .A(n_80), .Y(n_1424) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_81), .A2(n_95), .B1(n_902), .B2(n_904), .Y(n_912) );
INVx1_ASAP7_75t_L g946 ( .A(n_81), .Y(n_946) );
INVxp33_ASAP7_75t_L g1128 ( .A(n_82), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_83), .Y(n_1065) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_84), .A2(n_206), .B1(n_1080), .B2(n_1082), .C(n_1085), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_84), .Y(n_1108) );
AOI221xp5_ASAP7_75t_SL g1747 ( .A1(n_85), .A2(n_92), .B1(n_535), .B2(n_603), .C(n_840), .Y(n_1747) );
INVx1_ASAP7_75t_L g1760 ( .A(n_85), .Y(n_1760) );
INVxp33_ASAP7_75t_L g968 ( .A(n_86), .Y(n_968) );
INVx1_ASAP7_75t_L g1743 ( .A(n_87), .Y(n_1743) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_88), .A2(n_623), .B1(n_699), .B2(n_700), .Y(n_622) );
INVx1_ASAP7_75t_L g699 ( .A(n_88), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_89), .A2(n_103), .B1(n_764), .B2(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g440 ( .A(n_90), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g1780 ( .A1(n_91), .A2(n_1735), .B1(n_1781), .B2(n_1782), .Y(n_1780) );
CKINVDCx5p33_ASAP7_75t_R g1782 ( .A(n_91), .Y(n_1782) );
INVx1_ASAP7_75t_L g1759 ( .A(n_92), .Y(n_1759) );
XOR2x2_ASAP7_75t_L g1434 ( .A(n_93), .B(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1409 ( .A(n_94), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_95), .B(n_545), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_96), .A2(n_203), .B1(n_461), .B2(n_1339), .Y(n_1338) );
CKINVDCx5p33_ASAP7_75t_R g1379 ( .A(n_96), .Y(n_1379) );
CKINVDCx16_ASAP7_75t_R g1539 ( .A(n_98), .Y(n_1539) );
INVx1_ASAP7_75t_L g989 ( .A(n_99), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_100), .Y(n_476) );
INVxp67_ASAP7_75t_L g963 ( .A(n_101), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_101), .A2(n_134), .B1(n_715), .B2(n_857), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_102), .A2(n_237), .B1(n_607), .B2(n_937), .Y(n_1456) );
OAI211xp5_ASAP7_75t_L g1458 ( .A1(n_102), .A2(n_1459), .B(n_1460), .C(n_1462), .Y(n_1458) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_103), .A2(n_159), .B1(n_505), .B2(n_726), .C(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1005 ( .A(n_104), .Y(n_1005) );
OAI22xp33_ASAP7_75t_SL g1241 ( .A1(n_105), .A2(n_140), .B1(n_717), .B2(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1265 ( .A(n_105), .Y(n_1265) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_106), .Y(n_1015) );
INVx1_ASAP7_75t_L g1139 ( .A(n_107), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1750 ( .A1(n_108), .A2(n_168), .B1(n_505), .B2(n_614), .C(n_616), .Y(n_1750) );
AOI221xp5_ASAP7_75t_L g1767 ( .A1(n_108), .A2(n_161), .B1(n_1768), .B2(n_1769), .C(n_1771), .Y(n_1767) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_109), .B(n_557), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g1513 ( .A1(n_111), .A2(n_295), .B1(n_1479), .B2(n_1514), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_112), .Y(n_1230) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_113), .Y(n_659) );
OAI222xp33_ASAP7_75t_L g860 ( .A1(n_114), .A2(n_177), .B1(n_307), .B2(n_830), .C1(n_861), .C2(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g873 ( .A(n_114), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_115), .A2(n_282), .B1(n_531), .B2(n_726), .C(n_729), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_115), .A2(n_198), .B1(n_658), .B2(n_758), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g1439 ( .A1(n_116), .A2(n_286), .B1(n_500), .B2(n_1228), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1468 ( .A1(n_116), .A2(n_166), .B1(n_752), .B2(n_766), .Y(n_1468) );
INVxp67_ASAP7_75t_L g962 ( .A(n_117), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_117), .A2(n_174), .B1(n_602), .B2(n_603), .C(n_720), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g1457 ( .A1(n_118), .A2(n_823), .B(n_824), .Y(n_1457) );
INVx1_ASAP7_75t_L g1463 ( .A(n_118), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1438 ( .A1(n_119), .A2(n_166), .B1(n_1238), .B2(n_1242), .Y(n_1438) );
AOI22xp5_ASAP7_75t_L g1467 ( .A1(n_119), .A2(n_286), .B1(n_392), .B2(n_907), .Y(n_1467) );
AOI22xp5_ASAP7_75t_L g1553 ( .A1(n_120), .A2(n_125), .B1(n_1508), .B2(n_1511), .Y(n_1553) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_121), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_122), .A2(n_154), .B1(n_407), .B2(n_567), .C(n_569), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_122), .A2(n_154), .B1(n_828), .B2(n_830), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_123), .A2(n_278), .B1(n_614), .B2(n_1176), .C(n_1302), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_123), .A2(n_278), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
XNOR2xp5_ASAP7_75t_L g1120 ( .A(n_124), .B(n_1121), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_124), .A2(n_306), .B1(n_1491), .B2(n_1555), .Y(n_1554) );
CKINVDCx5p33_ASAP7_75t_R g1446 ( .A(n_126), .Y(n_1446) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_127), .A2(n_163), .B1(n_396), .B2(n_406), .C(n_965), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_127), .A2(n_163), .B1(n_610), .B2(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1461 ( .A(n_128), .Y(n_1461) );
INVx1_ASAP7_75t_L g1745 ( .A(n_129), .Y(n_1745) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_130), .A2(n_277), .B1(n_531), .B2(n_615), .C(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g887 ( .A(n_130), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g1353 ( .A(n_131), .Y(n_1353) );
INVx1_ASAP7_75t_L g359 ( .A(n_132), .Y(n_359) );
AO221x2_ASAP7_75t_L g1490 ( .A1(n_132), .A2(n_191), .B1(n_1479), .B2(n_1491), .C(n_1493), .Y(n_1490) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_133), .Y(n_663) );
INVxp67_ASAP7_75t_L g958 ( .A(n_134), .Y(n_958) );
INVx1_ASAP7_75t_L g588 ( .A(n_135), .Y(n_588) );
INVxp33_ASAP7_75t_SL g1306 ( .A(n_136), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_136), .A2(n_262), .B1(n_763), .B2(n_1322), .Y(n_1324) );
INVx1_ASAP7_75t_L g1483 ( .A(n_137), .Y(n_1483) );
INVx1_ASAP7_75t_L g1637 ( .A(n_138), .Y(n_1637) );
AOI22xp5_ASAP7_75t_L g1542 ( .A1(n_139), .A2(n_316), .B1(n_1508), .B2(n_1511), .Y(n_1542) );
INVx1_ASAP7_75t_L g1259 ( .A(n_140), .Y(n_1259) );
INVx1_ASAP7_75t_L g930 ( .A(n_141), .Y(n_930) );
INVx1_ASAP7_75t_L g443 ( .A(n_142), .Y(n_443) );
INVxp67_ASAP7_75t_L g1137 ( .A(n_143), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_143), .A2(n_182), .B1(n_818), .B2(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g592 ( .A(n_145), .Y(n_592) );
INVx1_ASAP7_75t_L g1481 ( .A(n_146), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1502 ( .A(n_146), .B(n_1499), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1748 ( .A1(n_147), .A2(n_221), .B1(n_673), .B2(n_1378), .Y(n_1748) );
OAI221xp5_ASAP7_75t_L g1756 ( .A1(n_147), .A2(n_221), .B1(n_422), .B2(n_1757), .C(n_1758), .Y(n_1756) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_148), .A2(n_198), .B1(n_508), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_148), .A2(n_282), .B1(n_752), .B2(n_754), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_149), .A2(n_682), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g772 ( .A(n_149), .Y(n_772) );
INVx1_ASAP7_75t_L g1143 ( .A(n_150), .Y(n_1143) );
INVx2_ASAP7_75t_L g347 ( .A(n_151), .Y(n_347) );
INVx1_ASAP7_75t_L g499 ( .A(n_152), .Y(n_499) );
BUFx3_ASAP7_75t_L g473 ( .A(n_153), .Y(n_473) );
INVx1_ASAP7_75t_L g503 ( .A(n_153), .Y(n_503) );
INVx1_ASAP7_75t_L g1181 ( .A(n_155), .Y(n_1181) );
INVx1_ASAP7_75t_L g1494 ( .A(n_157), .Y(n_1494) );
INVx1_ASAP7_75t_L g638 ( .A(n_158), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_158), .A2(n_264), .B1(n_536), .B2(n_692), .Y(n_691) );
INVxp33_ASAP7_75t_L g785 ( .A(n_162), .Y(n_785) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_162), .A2(n_202), .B1(n_615), .B2(n_823), .C(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g627 ( .A(n_164), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_165), .Y(n_1229) );
CKINVDCx5p33_ASAP7_75t_R g1413 ( .A(n_167), .Y(n_1413) );
INVx1_ASAP7_75t_L g1773 ( .A(n_168), .Y(n_1773) );
INVxp67_ASAP7_75t_L g418 ( .A(n_169), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_169), .A2(n_297), .B1(n_534), .B2(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g1635 ( .A(n_170), .Y(n_1635) );
OAI221xp5_ASAP7_75t_SL g1069 ( .A1(n_171), .A2(n_313), .B1(n_828), .B2(n_1070), .C(n_1072), .Y(n_1069) );
OAI221xp5_ASAP7_75t_L g1101 ( .A1(n_171), .A2(n_313), .B1(n_396), .B2(n_407), .C(n_635), .Y(n_1101) );
INVx1_ASAP7_75t_L g388 ( .A(n_172), .Y(n_388) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_173), .Y(n_1182) );
INVxp67_ASAP7_75t_L g959 ( .A(n_174), .Y(n_959) );
INVx1_ASAP7_75t_L g1744 ( .A(n_175), .Y(n_1744) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_176), .Y(n_1351) );
INVx1_ASAP7_75t_L g867 ( .A(n_177), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_178), .A2(n_269), .B1(n_732), .B2(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g872 ( .A(n_178), .Y(n_872) );
INVxp33_ASAP7_75t_SL g1204 ( .A(n_179), .Y(n_1204) );
INVx1_ASAP7_75t_L g1500 ( .A(n_180), .Y(n_1500) );
INVxp67_ASAP7_75t_L g581 ( .A(n_181), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_181), .A2(n_236), .B1(n_606), .B2(n_619), .Y(n_618) );
INVxp33_ASAP7_75t_L g1133 ( .A(n_182), .Y(n_1133) );
INVx1_ASAP7_75t_L g1091 ( .A(n_183), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1410 ( .A1(n_184), .A2(n_284), .B1(n_505), .B2(n_508), .C(n_682), .Y(n_1410) );
INVxp33_ASAP7_75t_SL g1419 ( .A(n_184), .Y(n_1419) );
INVx1_ASAP7_75t_L g468 ( .A(n_185), .Y(n_468) );
INVx1_ASAP7_75t_L g516 ( .A(n_185), .Y(n_516) );
INVx1_ASAP7_75t_L g1742 ( .A(n_187), .Y(n_1742) );
INVxp33_ASAP7_75t_SL g782 ( .A(n_188), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_188), .A2(n_194), .B1(n_614), .B2(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1526 ( .A(n_189), .Y(n_1526) );
INVx1_ASAP7_75t_L g1404 ( .A(n_190), .Y(n_1404) );
OAI221xp5_ASAP7_75t_L g1420 ( .A1(n_190), .A2(n_223), .B1(n_567), .B2(n_568), .C(n_635), .Y(n_1420) );
INVx1_ASAP7_75t_L g800 ( .A(n_192), .Y(n_800) );
INVxp33_ASAP7_75t_SL g786 ( .A(n_194), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_195), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_196), .A2(n_288), .B1(n_687), .B2(n_1021), .C(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1269 ( .A(n_196), .Y(n_1269) );
INVx1_ASAP7_75t_L g585 ( .A(n_197), .Y(n_585) );
INVx1_ASAP7_75t_L g775 ( .A(n_199), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g839 ( .A1(n_200), .A2(n_283), .B1(n_535), .B2(n_603), .C(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g870 ( .A(n_200), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g1507 ( .A1(n_201), .A2(n_265), .B1(n_1508), .B2(n_1511), .Y(n_1507) );
INVxp33_ASAP7_75t_L g783 ( .A(n_202), .Y(n_783) );
INVx1_ASAP7_75t_L g596 ( .A(n_204), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_205), .Y(n_898) );
INVx1_ASAP7_75t_L g1106 ( .A(n_206), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_207), .A2(n_213), .B1(n_726), .B2(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1034 ( .A(n_207), .Y(n_1034) );
INVx1_ASAP7_75t_L g1050 ( .A(n_208), .Y(n_1050) );
INVxp67_ASAP7_75t_L g974 ( .A(n_209), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_209), .A2(n_222), .B1(n_524), .B2(n_690), .C(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_210), .A2(n_274), .B1(n_859), .B2(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1105 ( .A(n_210), .Y(n_1105) );
INVx1_ASAP7_75t_L g1471 ( .A(n_211), .Y(n_1471) );
INVxp67_ASAP7_75t_L g1136 ( .A(n_212), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_212), .A2(n_322), .B1(n_505), .B2(n_616), .C(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1039 ( .A(n_213), .Y(n_1039) );
XNOR2xp5_ASAP7_75t_L g1006 ( .A(n_214), .B(n_1007), .Y(n_1006) );
CKINVDCx16_ASAP7_75t_R g1522 ( .A(n_215), .Y(n_1522) );
OAI211xp5_ASAP7_75t_SL g1183 ( .A1(n_216), .A2(n_1184), .B(n_1185), .C(n_1190), .Y(n_1183) );
INVx1_ASAP7_75t_L g1211 ( .A(n_216), .Y(n_1211) );
INVx1_ASAP7_75t_L g925 ( .A(n_217), .Y(n_925) );
OAI211xp5_ASAP7_75t_L g944 ( .A1(n_217), .A2(n_861), .B(n_945), .C(n_950), .Y(n_944) );
CKINVDCx5p33_ASAP7_75t_R g1376 ( .A(n_218), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1354 ( .A(n_219), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_220), .A2(n_267), .B1(n_1088), .B2(n_1173), .Y(n_1399) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_220), .Y(n_1423) );
INVxp33_ASAP7_75t_L g971 ( .A(n_222), .Y(n_971) );
INVx1_ASAP7_75t_L g1405 ( .A(n_223), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_224), .A2(n_233), .B1(n_524), .B2(n_607), .Y(n_1075) );
INVxp33_ASAP7_75t_L g1099 ( .A(n_224), .Y(n_1099) );
INVx1_ASAP7_75t_L g646 ( .A(n_225), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_225), .A2(n_241), .B1(n_687), .B2(n_689), .C(n_690), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_226), .Y(n_598) );
XNOR2x1_ASAP7_75t_L g835 ( .A(n_227), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g1401 ( .A(n_228), .Y(n_1401) );
INVx1_ASAP7_75t_L g441 ( .A(n_229), .Y(n_441) );
BUFx3_ASAP7_75t_L g475 ( .A(n_230), .Y(n_475) );
INVx1_ASAP7_75t_L g483 ( .A(n_230), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_231), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g1347 ( .A(n_232), .Y(n_1347) );
INVxp33_ASAP7_75t_L g1095 ( .A(n_233), .Y(n_1095) );
INVx1_ASAP7_75t_L g1117 ( .A(n_234), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_235), .Y(n_343) );
AND2x2_ASAP7_75t_L g372 ( .A(n_235), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_235), .B(n_303), .Y(n_404) );
INVx1_ASAP7_75t_L g455 ( .A(n_235), .Y(n_455) );
INVxp67_ASAP7_75t_L g576 ( .A(n_236), .Y(n_576) );
INVx1_ASAP7_75t_L g1464 ( .A(n_237), .Y(n_1464) );
AOI21xp5_ASAP7_75t_L g1293 ( .A1(n_238), .A2(n_1294), .B(n_1297), .Y(n_1293) );
INVx1_ASAP7_75t_L g1314 ( .A(n_238), .Y(n_1314) );
OAI332xp33_ASAP7_75t_L g1342 ( .A1(n_239), .A2(n_413), .A3(n_451), .B1(n_1343), .B2(n_1346), .B3(n_1349), .C1(n_1352), .C2(n_1355), .Y(n_1342) );
INVx1_ASAP7_75t_L g1383 ( .A(n_239), .Y(n_1383) );
INVx1_ASAP7_75t_L g1641 ( .A(n_240), .Y(n_1641) );
INVx1_ASAP7_75t_L g641 ( .A(n_241), .Y(n_641) );
INVx1_ASAP7_75t_L g1527 ( .A(n_243), .Y(n_1527) );
INVx2_ASAP7_75t_L g470 ( .A(n_244), .Y(n_470) );
OR2x2_ASAP7_75t_L g485 ( .A(n_244), .B(n_468), .Y(n_485) );
INVx1_ASAP7_75t_L g769 ( .A(n_245), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g1345 ( .A(n_246), .Y(n_1345) );
INVx1_ASAP7_75t_L g1639 ( .A(n_247), .Y(n_1639) );
INVx1_ASAP7_75t_L g980 ( .A(n_248), .Y(n_980) );
INVx1_ASAP7_75t_L g1412 ( .A(n_249), .Y(n_1412) );
INVxp67_ASAP7_75t_L g425 ( .A(n_250), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_250), .A2(n_296), .B1(n_523), .B2(n_525), .C(n_530), .Y(n_522) );
INVx1_ASAP7_75t_L g893 ( .A(n_251), .Y(n_893) );
CKINVDCx16_ASAP7_75t_R g1524 ( .A(n_252), .Y(n_1524) );
AOI222xp33_ASAP7_75t_L g1732 ( .A1(n_252), .A2(n_1733), .B1(n_1775), .B2(n_1779), .C1(n_1783), .C2(n_1787), .Y(n_1732) );
INVx1_ASAP7_75t_L g802 ( .A(n_253), .Y(n_802) );
INVxp33_ASAP7_75t_SL g1129 ( .A(n_254), .Y(n_1129) );
INVx1_ASAP7_75t_L g736 ( .A(n_255), .Y(n_736) );
INVxp67_ASAP7_75t_SL g1186 ( .A(n_256), .Y(n_1186) );
OAI211xp5_ASAP7_75t_SL g1200 ( .A1(n_256), .A2(n_433), .B(n_969), .C(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1397 ( .A(n_257), .Y(n_1397) );
INVx1_ASAP7_75t_L g1078 ( .A(n_258), .Y(n_1078) );
INVx1_ASAP7_75t_L g1532 ( .A(n_259), .Y(n_1532) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_260), .A2(n_280), .B1(n_606), .B2(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g885 ( .A(n_260), .Y(n_885) );
INVx1_ASAP7_75t_L g446 ( .A(n_261), .Y(n_446) );
INVxp67_ASAP7_75t_SL g1300 ( .A(n_262), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_263), .A2(n_272), .B1(n_614), .B2(n_1159), .C(n_1289), .Y(n_1288) );
INVxp33_ASAP7_75t_L g1313 ( .A(n_263), .Y(n_1313) );
INVx1_ASAP7_75t_L g650 ( .A(n_264), .Y(n_650) );
INVx1_ASAP7_75t_L g1407 ( .A(n_266), .Y(n_1407) );
INVxp67_ASAP7_75t_L g1428 ( .A(n_267), .Y(n_1428) );
INVx1_ASAP7_75t_L g916 ( .A(n_268), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_268), .A2(n_514), .B(n_693), .Y(n_942) );
INVx1_ASAP7_75t_L g869 ( .A(n_269), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_270), .Y(n_631) );
INVxp33_ASAP7_75t_L g1205 ( .A(n_271), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1223 ( .A(n_273), .Y(n_1223) );
INVx1_ASAP7_75t_L g1111 ( .A(n_274), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_275), .Y(n_653) );
INVx1_ASAP7_75t_L g920 ( .A(n_276), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_277), .A2(n_280), .B1(n_880), .B2(n_882), .C(n_884), .Y(n_879) );
INVx1_ASAP7_75t_L g1518 ( .A(n_279), .Y(n_1518) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_281), .A2(n_315), .B1(n_619), .B2(n_826), .Y(n_1026) );
INVx1_ASAP7_75t_L g1052 ( .A(n_281), .Y(n_1052) );
INVx1_ASAP7_75t_L g878 ( .A(n_283), .Y(n_878) );
INVxp33_ASAP7_75t_SL g1417 ( .A(n_284), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_285), .Y(n_852) );
INVx1_ASAP7_75t_L g988 ( .A(n_287), .Y(n_988) );
INVx1_ASAP7_75t_L g1271 ( .A(n_288), .Y(n_1271) );
INVx1_ASAP7_75t_L g734 ( .A(n_289), .Y(n_734) );
INVx1_ASAP7_75t_L g1073 ( .A(n_290), .Y(n_1073) );
INVx1_ASAP7_75t_L g777 ( .A(n_291), .Y(n_777) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
AND3x2_ASAP7_75t_L g1482 ( .A(n_292), .B(n_335), .C(n_1483), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1497 ( .A(n_292), .B(n_335), .Y(n_1497) );
INVx2_ASAP7_75t_L g348 ( .A(n_294), .Y(n_348) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_296), .Y(n_432) );
INVxp33_ASAP7_75t_SL g421 ( .A(n_297), .Y(n_421) );
INVx1_ASAP7_75t_L g710 ( .A(n_298), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g1344 ( .A(n_300), .Y(n_1344) );
INVx1_ASAP7_75t_L g805 ( .A(n_301), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_302), .Y(n_1246) );
INVx1_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
INVx2_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g1245 ( .A(n_304), .Y(n_1245) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_305), .Y(n_799) );
INVx1_ASAP7_75t_L g866 ( .A(n_307), .Y(n_866) );
INVxp33_ASAP7_75t_L g564 ( .A(n_308), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_308), .A2(n_309), .B1(n_535), .B2(n_602), .C(n_603), .Y(n_601) );
INVxp33_ASAP7_75t_L g562 ( .A(n_309), .Y(n_562) );
INVxp67_ASAP7_75t_SL g1284 ( .A(n_310), .Y(n_1284) );
INVx1_ASAP7_75t_L g803 ( .A(n_311), .Y(n_803) );
INVxp67_ASAP7_75t_SL g1326 ( .A(n_312), .Y(n_1326) );
INVx1_ASAP7_75t_L g1533 ( .A(n_314), .Y(n_1533) );
INVx1_ASAP7_75t_L g1045 ( .A(n_315), .Y(n_1045) );
INVx1_ASAP7_75t_L g1189 ( .A(n_317), .Y(n_1189) );
INVx1_ASAP7_75t_L g1256 ( .A(n_318), .Y(n_1256) );
INVx1_ASAP7_75t_L g1161 ( .A(n_319), .Y(n_1161) );
CKINVDCx5p33_ASAP7_75t_R g1281 ( .A(n_320), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_321), .Y(n_1013) );
INVxp33_ASAP7_75t_L g1134 ( .A(n_322), .Y(n_1134) );
INVx1_ASAP7_75t_L g1090 ( .A(n_323), .Y(n_1090) );
INVx1_ASAP7_75t_L g806 ( .A(n_324), .Y(n_806) );
INVxp33_ASAP7_75t_SL g382 ( .A(n_325), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_326), .Y(n_718) );
INVx1_ASAP7_75t_L g741 ( .A(n_327), .Y(n_741) );
INVxp33_ASAP7_75t_L g561 ( .A(n_328), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_351), .B(n_1475), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_338), .Y(n_332) );
AND2x4_ASAP7_75t_L g1778 ( .A(n_333), .B(n_339), .Y(n_1778) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_SL g1786 ( .A(n_334), .Y(n_1786) );
NAND2xp5_ASAP7_75t_L g1793 ( .A(n_334), .B(n_336), .Y(n_1793) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_336), .B(n_1786), .Y(n_1785) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_344), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g750 ( .A(n_342), .B(n_350), .Y(n_750) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g414 ( .A(n_343), .B(n_415), .Y(n_414) );
OR2x6_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g420 ( .A(n_345), .Y(n_420) );
OR2x2_ASAP7_75t_L g461 ( .A(n_345), .B(n_403), .Y(n_461) );
INVx2_ASAP7_75t_SL g580 ( .A(n_345), .Y(n_580) );
INVx2_ASAP7_75t_SL g591 ( .A(n_345), .Y(n_591) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_345), .Y(n_652) );
BUFx2_ASAP7_75t_L g886 ( .A(n_345), .Y(n_886) );
OAI22xp33_ASAP7_75t_L g892 ( .A1(n_345), .A2(n_435), .B1(n_852), .B2(n_893), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_345), .A2(n_435), .B1(n_1446), .B2(n_1471), .Y(n_1470) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_L g367 ( .A(n_347), .Y(n_367) );
INVx1_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
AND2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_348), .Y(n_387) );
AND2x4_ASAP7_75t_L g394 ( .A(n_347), .B(n_380), .Y(n_394) );
INVx1_ASAP7_75t_L g438 ( .A(n_347), .Y(n_438) );
INVx1_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
INVx2_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
INVx1_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_348), .B(n_367), .Y(n_431) );
INVx1_ASAP7_75t_L g437 ( .A(n_348), .Y(n_437) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_1057), .B2(n_1058), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_701), .B2(n_1056), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
XNOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_555), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
XNOR2x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_456), .Y(n_360) );
NOR3xp33_ASAP7_75t_SL g361 ( .A(n_362), .B(n_395), .C(n_411), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_364), .A2(n_384), .B1(n_564), .B2(n_565), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_364), .A2(n_384), .B1(n_1038), .B2(n_1039), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_364), .A2(n_384), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_370), .Y(n_364) );
AND2x2_ASAP7_75t_L g633 ( .A(n_365), .B(n_370), .Y(n_633) );
AND2x2_ASAP7_75t_L g774 ( .A(n_365), .B(n_370), .Y(n_774) );
AND2x2_ASAP7_75t_L g919 ( .A(n_365), .B(n_370), .Y(n_919) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_365), .B(n_370), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1209 ( .A(n_365), .Y(n_1209) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g758 ( .A(n_366), .Y(n_758) );
INVx1_ASAP7_75t_L g881 ( .A(n_366), .Y(n_881) );
INVx1_ASAP7_75t_L g890 ( .A(n_366), .Y(n_890) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_366), .Y(n_907) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_366), .Y(n_911) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g409 ( .A(n_367), .Y(n_409) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x6_ASAP7_75t_L g376 ( .A(n_370), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g384 ( .A(n_370), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g391 ( .A(n_370), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g876 ( .A(n_370), .B(n_877), .Y(n_876) );
AND2x2_ASAP7_75t_L g923 ( .A(n_370), .B(n_587), .Y(n_923) );
AND2x2_ASAP7_75t_L g960 ( .A(n_370), .B(n_766), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1755 ( .A1(n_370), .A2(n_767), .B1(n_1756), .B2(n_1762), .Y(n_1755) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g452 ( .A(n_371), .Y(n_452) );
INVx1_ASAP7_75t_L g415 ( .A(n_373), .Y(n_415) );
INVx1_ASAP7_75t_L g454 ( .A(n_373), .Y(n_454) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_375), .A2(n_628), .B1(n_1313), .B2(n_1314), .Y(n_1312) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_376), .A2(n_391), .B1(n_561), .B2(n_562), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_376), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_376), .A2(n_718), .B1(n_769), .B2(n_770), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_376), .A2(n_770), .B1(n_782), .B2(n_783), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_376), .A2(n_774), .B1(n_869), .B2(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_376), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_376), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_376), .A2(n_1073), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_376), .A2(n_1096), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
INVx1_ASAP7_75t_SL g1193 ( .A(n_376), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_376), .A2(n_391), .B1(n_1229), .B2(n_1269), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_376), .A2(n_390), .B1(n_1409), .B2(n_1417), .Y(n_1416) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_377), .B(n_402), .Y(n_410) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_377), .Y(n_1198) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g747 ( .A(n_378), .Y(n_747) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_378), .Y(n_756) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_378), .Y(n_766) );
INVx1_ASAP7_75t_L g905 ( .A(n_378), .Y(n_905) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B1(n_388), .B2(n_389), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g1247 ( .A1(n_383), .A2(n_1230), .B(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1311 ( .A(n_383), .Y(n_1311) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_384), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_384), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_384), .A2(n_774), .B1(n_785), .B2(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_384), .B(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_384), .A2(n_1098), .B1(n_1099), .B2(n_1100), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_384), .A2(n_1100), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_384), .A2(n_1100), .B1(n_1407), .B2(n_1419), .Y(n_1418) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g764 ( .A(n_386), .Y(n_764) );
INVx2_ASAP7_75t_SL g877 ( .A(n_386), .Y(n_877) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_387), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g497 ( .A1(n_388), .A2(n_498), .B1(n_499), .B2(n_500), .C(n_504), .Y(n_497) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g628 ( .A(n_391), .Y(n_628) );
BUFx2_ASAP7_75t_L g770 ( .A(n_391), .Y(n_770) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_391), .Y(n_1035) );
BUFx2_ASAP7_75t_L g1096 ( .A(n_391), .Y(n_1096) );
BUFx3_ASAP7_75t_L g658 ( .A(n_392), .Y(n_658) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g587 ( .A(n_393), .Y(n_587) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_393), .Y(n_909) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
INVx1_ASAP7_75t_L g986 ( .A(n_394), .Y(n_986) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g567 ( .A(n_397), .Y(n_567) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_398), .Y(n_1041) );
NAND2x1_ASAP7_75t_SL g398 ( .A(n_399), .B(n_402), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_399), .A2(n_408), .B1(n_1188), .B2(n_1189), .Y(n_1201) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_401), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_402), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g739 ( .A(n_402), .B(n_740), .Y(n_739) );
AND2x4_ASAP7_75t_L g742 ( .A(n_402), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g746 ( .A(n_402), .B(n_747), .Y(n_746) );
AOI32xp33_ASAP7_75t_L g1194 ( .A1(n_402), .A2(n_1195), .A3(n_1197), .B1(n_1199), .B2(n_1200), .Y(n_1194) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx4f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_407), .Y(n_568) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g569 ( .A(n_410), .Y(n_569) );
BUFx2_ASAP7_75t_L g635 ( .A(n_410), .Y(n_635) );
BUFx3_ASAP7_75t_L g965 ( .A(n_410), .Y(n_965) );
OAI33xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_417), .A3(n_424), .B1(n_439), .B2(n_442), .B3(n_447), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI33xp33_ASAP7_75t_L g570 ( .A1(n_413), .A2(n_449), .A3(n_571), .B1(n_578), .B2(n_584), .B3(n_589), .Y(n_570) );
OAI33xp33_ASAP7_75t_L g636 ( .A1(n_413), .A2(n_449), .A3(n_637), .B1(n_642), .B2(n_651), .B3(n_656), .Y(n_636) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_413), .Y(n_789) );
OAI33xp33_ASAP7_75t_L g966 ( .A1(n_413), .A2(n_967), .A3(n_973), .B1(n_979), .B2(n_987), .B3(n_990), .Y(n_966) );
OAI33xp33_ASAP7_75t_L g1042 ( .A1(n_413), .A2(n_449), .A3(n_1043), .B1(n_1049), .B2(n_1054), .B3(n_1055), .Y(n_1042) );
OAI33xp33_ASAP7_75t_L g1102 ( .A1(n_413), .A2(n_449), .A3(n_1103), .B1(n_1107), .B2(n_1112), .B3(n_1114), .Y(n_1102) );
OAI33xp33_ASAP7_75t_L g1248 ( .A1(n_413), .A2(n_1249), .A3(n_1255), .B1(n_1257), .B2(n_1263), .B3(n_1266), .Y(n_1248) );
OAI33xp33_ASAP7_75t_L g1421 ( .A1(n_413), .A2(n_1266), .A3(n_1422), .B1(n_1425), .B2(n_1429), .B3(n_1430), .Y(n_1421) );
OR2x6_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
BUFx2_ASAP7_75t_L g554 ( .A(n_416), .Y(n_554) );
INVx2_ASAP7_75t_L g698 ( .A(n_416), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_421), .B2(n_422), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g442 ( .A1(n_419), .A2(n_443), .B1(n_444), .B2(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g1104 ( .A(n_420), .Y(n_1104) );
INVx2_ASAP7_75t_L g1251 ( .A(n_420), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_422), .A2(n_426), .B1(n_440), .B2(n_441), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_422), .A2(n_796), .B1(n_1136), .B2(n_1137), .Y(n_1135) );
INVx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx4_ASAP7_75t_L g577 ( .A(n_423), .Y(n_577) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_423), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1770 ( .A(n_423), .Y(n_1770) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_432), .B2(n_433), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_426), .A2(n_1426), .B1(n_1427), .B2(n_1428), .Y(n_1425) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_426), .A2(n_1402), .B1(n_1412), .B2(n_1427), .Y(n_1429) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_428), .A2(n_1068), .B1(n_1091), .B2(n_1113), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_428), .A2(n_1113), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_428), .A2(n_577), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g981 ( .A(n_429), .Y(n_981) );
INVx2_ASAP7_75t_SL g1258 ( .A(n_429), .Y(n_1258) );
INVx2_ASAP7_75t_L g1757 ( .A(n_429), .Y(n_1757) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g575 ( .A(n_430), .Y(n_575) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g645 ( .A(n_431), .Y(n_645) );
INVx1_ASAP7_75t_L g798 ( .A(n_431), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_433), .A2(n_791), .B1(n_805), .B2(n_806), .Y(n_804) );
OAI22xp5_ASAP7_75t_SL g987 ( .A1(n_433), .A2(n_579), .B1(n_988), .B2(n_989), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_433), .A2(n_1012), .B1(n_1028), .B2(n_1044), .Y(n_1055) );
OAI22xp5_ASAP7_75t_SL g1352 ( .A1(n_433), .A2(n_652), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g582 ( .A(n_434), .Y(n_582) );
INVx2_ASAP7_75t_L g1212 ( .A(n_434), .Y(n_1212) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g445 ( .A(n_435), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_435), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_884) );
BUFx3_ASAP7_75t_L g1432 ( .A(n_435), .Y(n_1432) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g595 ( .A(n_437), .B(n_438), .Y(n_595) );
INVx1_ASAP7_75t_L g744 ( .A(n_438), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_440), .A2(n_479), .B(n_486), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_441), .A2(n_443), .B1(n_544), .B2(n_549), .Y(n_543) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_445), .A2(n_1251), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_446), .A2(n_518), .B1(n_522), .B2(n_533), .C(n_538), .Y(n_517) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI33xp33_ASAP7_75t_L g1316 ( .A1(n_448), .A2(n_1317), .A3(n_1319), .B1(n_1320), .B2(n_1323), .B3(n_1324), .Y(n_1316) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI33xp33_ASAP7_75t_L g788 ( .A1(n_449), .A2(n_789), .A3(n_790), .B1(n_795), .B2(n_801), .B3(n_804), .Y(n_788) );
OAI33xp33_ASAP7_75t_L g1131 ( .A1(n_449), .A2(n_789), .A3(n_1132), .B1(n_1135), .B2(n_1138), .B3(n_1141), .Y(n_1131) );
CKINVDCx8_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
INVx5_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx6_ASAP7_75t_L g767 ( .A(n_451), .Y(n_767) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx2_ASAP7_75t_L g914 ( .A(n_453), .Y(n_914) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_476), .B(n_477), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI21xp33_ASAP7_75t_SL g597 ( .A1(n_459), .A2(n_598), .B(n_599), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_459), .A2(n_707), .B1(n_708), .B2(n_736), .Y(n_706) );
AOI21xp33_ASAP7_75t_SL g1064 ( .A1(n_459), .A2(n_1065), .B(n_1066), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_459), .A2(n_1392), .B1(n_1395), .B2(n_1413), .Y(n_1391) );
INVx5_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g662 ( .A(n_460), .Y(n_662) );
INVx1_ASAP7_75t_L g832 ( .A(n_460), .Y(n_832) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_460), .Y(n_1004) );
INVx2_ASAP7_75t_L g1030 ( .A(n_460), .Y(n_1030) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx2_ASAP7_75t_L g874 ( .A(n_461), .Y(n_874) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_L g861 ( .A(n_465), .Y(n_861) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_471), .Y(n_465) );
AND2x4_ASAP7_75t_L g488 ( .A(n_466), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_466), .Y(n_493) );
AND2x4_ASAP7_75t_L g611 ( .A(n_466), .B(n_495), .Y(n_611) );
AND2x2_ASAP7_75t_L g669 ( .A(n_466), .B(n_495), .Y(n_669) );
AND2x4_ASAP7_75t_L g829 ( .A(n_466), .B(n_489), .Y(n_829) );
BUFx2_ASAP7_75t_L g850 ( .A(n_466), .Y(n_850) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_466), .B(n_495), .Y(n_1071) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g515 ( .A(n_469), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g532 ( .A(n_470), .B(n_516), .Y(n_532) );
INVx6_ASAP7_75t_L g511 ( .A(n_471), .Y(n_511) );
BUFx2_ASAP7_75t_L g823 ( .A(n_471), .Y(n_823) );
INVx2_ASAP7_75t_L g1018 ( .A(n_471), .Y(n_1018) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g496 ( .A(n_472), .Y(n_496) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g482 ( .A(n_473), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g507 ( .A(n_473), .B(n_475), .Y(n_507) );
INVx1_ASAP7_75t_L g491 ( .A(n_474), .Y(n_491) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_L g502 ( .A(n_475), .B(n_503), .Y(n_502) );
AOI31xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_517), .A3(n_543), .B(n_552), .Y(n_477) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_480), .A2(n_585), .B1(n_601), .B2(n_604), .C(n_608), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_480), .A2(n_655), .B(n_666), .C(n_670), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_480), .A2(n_544), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g1067 ( .A1(n_480), .A2(n_1068), .B(n_1069), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_480), .A2(n_544), .B1(n_1139), .B2(n_1142), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_480), .A2(n_544), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
INVx1_ASAP7_75t_L g1286 ( .A(n_480), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_480), .B(n_1412), .Y(n_1411) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_484), .Y(n_480) );
INVx2_ASAP7_75t_SL g498 ( .A(n_481), .Y(n_498) );
INVx1_ASAP7_75t_L g672 ( .A(n_481), .Y(n_672) );
BUFx3_ASAP7_75t_L g1378 ( .A(n_481), .Y(n_1378) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_482), .Y(n_524) );
BUFx2_ASAP7_75t_L g614 ( .A(n_482), .Y(n_614) );
INVx2_ASAP7_75t_SL g688 ( .A(n_482), .Y(n_688) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_482), .Y(n_728) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_482), .Y(n_814) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_482), .Y(n_845) );
BUFx2_ASAP7_75t_L g857 ( .A(n_482), .Y(n_857) );
BUFx3_ASAP7_75t_L g937 ( .A(n_482), .Y(n_937) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_482), .Y(n_1157) );
INVx1_ASAP7_75t_L g548 ( .A(n_483), .Y(n_548) );
AND2x4_ASAP7_75t_L g521 ( .A(n_484), .B(n_506), .Y(n_521) );
AND2x2_ASAP7_75t_L g813 ( .A(n_484), .B(n_814), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_484), .A2(n_544), .B1(n_852), .B2(n_853), .C(n_860), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_484), .A2(n_602), .B(n_946), .C(n_947), .Y(n_945) );
OAI21xp33_ASAP7_75t_L g1236 ( .A1(n_484), .A2(n_1237), .B(n_1241), .Y(n_1236) );
OAI21xp5_ASAP7_75t_L g1437 ( .A1(n_484), .A2(n_1438), .B(n_1439), .Y(n_1437) );
AOI222xp33_ASAP7_75t_L g1737 ( .A1(n_484), .A2(n_488), .B1(n_1071), .B2(n_1738), .C1(n_1744), .C2(n_1745), .Y(n_1737) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g545 ( .A(n_485), .B(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g550 ( .A(n_485), .B(n_551), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_SL g1357 ( .A1(n_485), .A2(n_1358), .B(n_1362), .C(n_1367), .Y(n_1357) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g609 ( .A(n_488), .Y(n_609) );
INVx1_ASAP7_75t_L g667 ( .A(n_488), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g1185 ( .A1(n_488), .A2(n_669), .B1(n_1186), .B2(n_1187), .C1(n_1188), .C2(n_1189), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_488), .A2(n_1071), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
INVxp67_ASAP7_75t_L g1443 ( .A(n_489), .Y(n_1443) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_SL g541 ( .A(n_493), .Y(n_541) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g1444 ( .A(n_495), .Y(n_1444) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g605 ( .A(n_498), .Y(n_605) );
INVx1_ASAP7_75t_L g732 ( .A(n_500), .Y(n_732) );
INVx1_ASAP7_75t_L g1159 ( .A(n_500), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_500), .A2(n_1376), .B1(n_1377), .B2(n_1379), .Y(n_1375) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g537 ( .A(n_501), .Y(n_537) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_501), .Y(n_859) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_501), .Y(n_1002) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g551 ( .A(n_502), .Y(n_551) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
INVx1_ASAP7_75t_L g674 ( .A(n_502), .Y(n_674) );
INVx1_ASAP7_75t_L g1361 ( .A(n_502), .Y(n_1361) );
INVx1_ASAP7_75t_L g547 ( .A(n_503), .Y(n_547) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx4f_ASAP7_75t_L g602 ( .A(n_506), .Y(n_602) );
INVx2_ASAP7_75t_SL g841 ( .A(n_506), .Y(n_841) );
AND2x4_ASAP7_75t_L g849 ( .A(n_506), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g1149 ( .A(n_506), .Y(n_1149) );
BUFx6f_ASAP7_75t_L g1366 ( .A(n_506), .Y(n_1366) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_507), .Y(n_529) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_510), .Y(n_535) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_511), .Y(n_620) );
INVx1_ASAP7_75t_L g693 ( .A(n_511), .Y(n_693) );
INVx2_ASAP7_75t_L g720 ( .A(n_511), .Y(n_720) );
INVx2_ASAP7_75t_SL g820 ( .A(n_511), .Y(n_820) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_511), .Y(n_848) );
INVx1_ASAP7_75t_L g1752 ( .A(n_511), .Y(n_1752) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g1227 ( .A1(n_513), .A2(n_679), .B1(n_1228), .B2(n_1229), .C(n_1230), .Y(n_1227) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_515), .Y(n_603) );
INVx2_ASAP7_75t_L g682 ( .A(n_515), .Y(n_682) );
INVx1_ASAP7_75t_L g824 ( .A(n_515), .Y(n_824) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_520), .A2(n_540), .B1(n_596), .B2(n_613), .C(n_618), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_520), .A2(n_540), .B1(n_1078), .B2(n_1079), .C(n_1087), .Y(n_1077) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g685 ( .A(n_521), .Y(n_685) );
INVx2_ASAP7_75t_SL g723 ( .A(n_521), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_521), .A2(n_849), .B1(n_989), .B2(n_999), .C(n_1001), .Y(n_998) );
INVx1_ASAP7_75t_L g1155 ( .A(n_521), .Y(n_1155) );
INVx1_ASAP7_75t_L g1184 ( .A(n_521), .Y(n_1184) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g714 ( .A(n_524), .Y(n_714) );
BUFx3_ASAP7_75t_L g843 ( .A(n_524), .Y(n_843) );
INVx1_ASAP7_75t_L g948 ( .A(n_524), .Y(n_948) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g689 ( .A(n_526), .Y(n_689) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_529), .Y(n_542) );
BUFx6f_ASAP7_75t_L g1000 ( .A(n_529), .Y(n_1000) );
INVx1_ASAP7_75t_L g1084 ( .A(n_529), .Y(n_1084) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g1086 ( .A(n_531), .Y(n_1086) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g617 ( .A(n_532), .Y(n_617) );
INVx1_ASAP7_75t_L g690 ( .A(n_532), .Y(n_690) );
INVx2_ASAP7_75t_L g1451 ( .A(n_532), .Y(n_1451) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_540), .A2(n_660), .B1(n_684), .B2(n_686), .C(n_691), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_540), .A2(n_722), .B1(n_724), .B2(n_725), .C(n_731), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_540), .A2(n_722), .B1(n_806), .B2(n_816), .C(n_817), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_540), .A2(n_1143), .B1(n_1154), .B2(n_1156), .C(n_1158), .Y(n_1153) );
INVx1_ASAP7_75t_L g1190 ( .A(n_540), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_540), .Y(n_1304) );
INVx1_ASAP7_75t_L g1367 ( .A(n_540), .Y(n_1367) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_540), .A2(n_1154), .B1(n_1397), .B2(n_1398), .C(n_1399), .Y(n_1396) );
AOI21xp33_ASAP7_75t_L g1746 ( .A1(n_540), .A2(n_1747), .B(n_1748), .Y(n_1746) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_542), .Y(n_615) );
INVx1_ASAP7_75t_L g730 ( .A(n_542), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g1741 ( .A1(n_542), .A2(n_814), .B1(n_1742), .B2(n_1743), .Y(n_1741) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_544), .A2(n_549), .B1(n_588), .B2(n_592), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_544), .A2(n_549), .B1(n_653), .B2(n_659), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_544), .A2(n_802), .B1(n_805), .B2(n_811), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g1003 ( .A1(n_544), .A2(n_549), .B1(n_982), .B2(n_988), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_544), .A2(n_813), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_544), .A2(n_549), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_544), .A2(n_549), .B1(n_1306), .B2(n_1307), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_544), .A2(n_549), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
INVx6_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g680 ( .A(n_546), .Y(n_680) );
INVx2_ASAP7_75t_L g1239 ( .A(n_546), .Y(n_1239) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g678 ( .A(n_547), .B(n_548), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_549), .A2(n_710), .B(n_711), .C(n_712), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_549), .A2(n_803), .B1(n_822), .B2(n_825), .C(n_827), .Y(n_821) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_549), .A2(n_1015), .B1(n_1016), .B2(n_1020), .C(n_1022), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_549), .A2(n_1140), .B1(n_1147), .B2(n_1150), .C(n_1152), .Y(n_1146) );
INVx4_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g826 ( .A(n_551), .Y(n_826) );
INVx2_ASAP7_75t_L g935 ( .A(n_551), .Y(n_935) );
AOI31xp33_ASAP7_75t_L g599 ( .A1(n_552), .A2(n_600), .A3(n_612), .B(n_621), .Y(n_599) );
INVx5_ASAP7_75t_L g808 ( .A(n_552), .Y(n_808) );
BUFx8_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g1009 ( .A(n_553), .Y(n_1009) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g707 ( .A(n_554), .Y(n_707) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_622), .Y(n_555) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_597), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_566), .C(n_570), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_576), .B2(n_577), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_573), .A2(n_585), .B1(n_586), .B2(n_588), .Y(n_584) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g1051 ( .A(n_574), .Y(n_1051) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g654 ( .A(n_575), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_577), .A2(n_796), .B1(n_799), .B2(n_800), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_577), .A2(n_654), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx2_ASAP7_75t_L g1196 ( .A(n_577), .Y(n_1196) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_578) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_579), .Y(n_1431) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g1422 ( .A1(n_582), .A2(n_1251), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
INVx2_ASAP7_75t_L g891 ( .A(n_586), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_586), .A2(n_643), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g649 ( .A(n_587), .Y(n_649) );
INVx2_ASAP7_75t_L g761 ( .A(n_587), .Y(n_761) );
INVx2_ASAP7_75t_L g883 ( .A(n_587), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B1(n_593), .B2(n_596), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_590), .A2(n_638), .B1(n_639), .B2(n_641), .Y(n_637) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g790 ( .A1(n_593), .A2(n_791), .B1(n_793), .B2(n_794), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_593), .A2(n_1078), .B1(n_1090), .B2(n_1115), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1132 ( .A1(n_593), .A2(n_791), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g1141 ( .A1(n_593), .A2(n_791), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
BUFx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g640 ( .A(n_594), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g1764 ( .A1(n_594), .A2(n_652), .B1(n_1743), .B2(n_1765), .Y(n_1764) );
OAI22xp5_ASAP7_75t_L g1771 ( .A1(n_594), .A2(n_652), .B1(n_1772), .B2(n_1773), .Y(n_1771) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g972 ( .A(n_595), .Y(n_972) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_595), .Y(n_1047) );
INVx2_ASAP7_75t_L g1254 ( .A(n_595), .Y(n_1254) );
INVx1_ASAP7_75t_L g1371 ( .A(n_606), .Y(n_1371) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g1021 ( .A(n_607), .Y(n_1021) );
INVx1_ASAP7_75t_L g1174 ( .A(n_607), .Y(n_1174) );
INVx1_ASAP7_75t_L g1240 ( .A(n_607), .Y(n_1240) );
INVx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g830 ( .A(n_611), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_611), .A2(n_829), .B1(n_898), .B2(n_899), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_611), .A2(n_1244), .B1(n_1245), .B2(n_1246), .Y(n_1243) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_615), .Y(n_1302) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g1176 ( .A(n_617), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_617), .A2(n_1295), .B1(n_1344), .B2(n_1348), .C(n_1373), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_619), .A2(n_1351), .B1(n_1353), .B2(n_1359), .Y(n_1358) );
INVx4_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g1233 ( .A(n_620), .Y(n_1233) );
INVx1_ASAP7_75t_L g700 ( .A(n_623), .Y(n_700) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_661), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_634), .C(n_636), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_630), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_628), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_629), .A2(n_631), .B1(n_676), .B2(n_679), .C(n_681), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_639), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_647), .B2(n_650), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g1763 ( .A(n_649), .Y(n_1763) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_651) );
INVx1_ASAP7_75t_L g792 ( .A(n_652), .Y(n_792) );
INVx1_ASAP7_75t_L g1116 ( .A(n_652), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B(n_664), .Y(n_661) );
AOI31xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_683), .A3(n_694), .B(n_695), .Y(n_664) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g1408 ( .A(n_673), .Y(n_1408) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g715 ( .A(n_674), .Y(n_715) );
INVx1_ASAP7_75t_L g1151 ( .A(n_674), .Y(n_1151) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_676), .A2(n_727), .B1(n_1223), .B2(n_1224), .C(n_1225), .Y(n_1222) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g717 ( .A(n_677), .Y(n_717) );
BUFx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g855 ( .A(n_678), .Y(n_855) );
BUFx4f_ASAP7_75t_L g932 ( .A(n_678), .Y(n_932) );
INVx2_ASAP7_75t_L g940 ( .A(n_678), .Y(n_940) );
INVx1_ASAP7_75t_L g1296 ( .A(n_678), .Y(n_1296) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g1297 ( .A(n_682), .Y(n_1297) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g1025 ( .A(n_688), .Y(n_1025) );
INVx1_ASAP7_75t_L g1225 ( .A(n_690), .Y(n_1225) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g1221 ( .A(n_693), .Y(n_1221) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_696), .A2(n_992), .B1(n_1004), .B2(n_1005), .Y(n_991) );
OAI31xp33_ASAP7_75t_L g1356 ( .A1(n_696), .A2(n_1357), .A3(n_1368), .B(n_1369), .Y(n_1356) );
CKINVDCx8_ASAP7_75t_R g696 ( .A(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g749 ( .A(n_698), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g913 ( .A(n_698), .B(n_914), .Y(n_913) );
AND2x4_ASAP7_75t_L g1199 ( .A(n_698), .B(n_750), .Y(n_1199) );
INVx2_ASAP7_75t_L g1394 ( .A(n_698), .Y(n_1394) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_702), .Y(n_1056) );
XNOR2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_833), .Y(n_702) );
XOR2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_776), .Y(n_703) );
XNOR2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_775), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_737), .Y(n_705) );
INVx2_ASAP7_75t_L g863 ( .A(n_707), .Y(n_863) );
OAI31xp33_ASAP7_75t_L g926 ( .A1(n_707), .A2(n_927), .A3(n_928), .B(n_944), .Y(n_926) );
OAI31xp33_ASAP7_75t_SL g1218 ( .A1(n_707), .A2(n_1219), .A3(n_1226), .B(n_1231), .Y(n_1218) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_709), .B(n_721), .C(n_733), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_718), .B(n_719), .Y(n_716) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_720), .Y(n_1088) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1027 ( .A(n_723), .Y(n_1027) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
BUFx3_ASAP7_75t_L g1374 ( .A(n_728), .Y(n_1374) );
A2O1A1Ixp33_ASAP7_75t_SL g1232 ( .A1(n_729), .A2(n_1233), .B(n_1234), .C(n_1235), .Y(n_1232) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND4x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_748), .C(n_768), .D(n_771), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_741), .B1(n_742), .B2(n_745), .C(n_746), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_739), .A2(n_742), .B1(n_746), .B2(n_866), .C(n_867), .Y(n_865) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_739), .A2(n_742), .B1(n_746), .B2(n_898), .C(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g1276 ( .A(n_739), .Y(n_1276) );
AOI221xp5_ASAP7_75t_L g1325 ( .A1(n_739), .A2(n_742), .B1(n_746), .B2(n_1326), .C(n_1327), .Y(n_1325) );
AOI21xp5_ASAP7_75t_L g1472 ( .A1(n_739), .A2(n_746), .B(n_1473), .Y(n_1472) );
AOI221xp5_ASAP7_75t_L g1774 ( .A1(n_739), .A2(n_742), .B1(n_746), .B2(n_1744), .C(n_1745), .Y(n_1774) );
INVx1_ASAP7_75t_L g1274 ( .A(n_742), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1460 ( .A1(n_742), .A2(n_874), .B1(n_1441), .B2(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g1272 ( .A1(n_746), .A2(n_1245), .B1(n_1246), .B2(n_1273), .C(n_1275), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_747), .Y(n_1322) );
AOI33xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .A3(n_757), .B1(n_759), .B2(n_762), .B3(n_767), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_749), .A2(n_767), .B1(n_876), .B2(n_878), .C1(n_879), .C2(n_888), .Y(n_875) );
AOI33xp33_ASAP7_75t_L g900 ( .A1(n_749), .A2(n_901), .A3(n_906), .B1(n_910), .B2(n_912), .B3(n_913), .Y(n_900) );
AOI322xp5_ASAP7_75t_L g1466 ( .A1(n_749), .A2(n_767), .A3(n_960), .B1(n_1453), .B2(n_1467), .C1(n_1468), .C2(n_1469), .Y(n_1466) );
AOI22xp5_ASAP7_75t_L g1766 ( .A1(n_749), .A2(n_874), .B1(n_1753), .B2(n_1767), .Y(n_1766) );
AOI22xp5_ASAP7_75t_L g1758 ( .A1(n_752), .A2(n_1759), .B1(n_1760), .B2(n_1761), .Y(n_1758) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g903 ( .A(n_753), .Y(n_903) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g1761 ( .A(n_755), .Y(n_1761) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g1321 ( .A(n_758), .Y(n_1321) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_761), .A2(n_1013), .B1(n_1015), .B2(n_1051), .Y(n_1054) );
BUFx3_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g990 ( .A(n_767), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_767), .A2(n_770), .B1(n_1207), .B2(n_1213), .Y(n_1206) );
INVx2_ASAP7_75t_L g1266 ( .A(n_767), .Y(n_1266) );
XNOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_807), .Y(n_778) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_787), .C(n_788), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_797), .A2(n_1108), .B1(n_1109), .B2(n_1111), .Y(n_1107) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g976 ( .A(n_798), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_809), .B1(n_831), .B2(n_832), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_808), .A2(n_1030), .B1(n_1145), .B2(n_1161), .Y(n_1144) );
OAI21xp33_ASAP7_75t_L g1169 ( .A1(n_808), .A2(n_1170), .B(n_1183), .Y(n_1169) );
INVx1_ASAP7_75t_SL g1308 ( .A(n_808), .Y(n_1308) );
NAND3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_815), .C(n_821), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g993 ( .A1(n_813), .A2(n_980), .B1(n_994), .B2(n_995), .C(n_996), .Y(n_993) );
INVx1_ASAP7_75t_L g1081 ( .A(n_814), .Y(n_1081) );
INVx1_ASAP7_75t_L g1242 ( .A(n_814), .Y(n_1242) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g1384 ( .A(n_824), .Y(n_1384) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_SL g862 ( .A(n_829), .Y(n_862) );
INVx4_ASAP7_75t_L g997 ( .A(n_829), .Y(n_997) );
AOI21xp5_ASAP7_75t_L g1280 ( .A1(n_832), .A2(n_1281), .B(n_1282), .Y(n_1280) );
XOR2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_951), .Y(n_833) );
XNOR2x1_ASAP7_75t_L g834 ( .A(n_835), .B(n_894), .Y(n_834) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_837), .B(n_864), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_851), .B(n_863), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_842), .B1(n_844), .B2(n_846), .C(n_849), .Y(n_838) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1019 ( .A(n_841), .Y(n_1019) );
INVx1_ASAP7_75t_L g1179 ( .A(n_841), .Y(n_1179) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g943 ( .A(n_849), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_849), .A2(n_1024), .B1(n_1026), .B2(n_1027), .C(n_1028), .Y(n_1023) );
BUFx3_ASAP7_75t_L g1235 ( .A(n_850), .Y(n_1235) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g1187 ( .A(n_861), .Y(n_1187) );
AOI31xp33_ASAP7_75t_L g1066 ( .A1(n_863), .A2(n_1067), .A3(n_1077), .B(n_1089), .Y(n_1066) );
NAND4xp25_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .C(n_871), .D(n_875), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_874), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g1270 ( .A1(n_874), .A2(n_1100), .B1(n_1234), .B2(n_1271), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_876), .A2(n_919), .B1(n_962), .B2(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g1355 ( .A(n_876), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1462 ( .A1(n_876), .A2(n_923), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1053 ( .A(n_882), .Y(n_1053) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_883), .Y(n_1113) );
INVx2_ASAP7_75t_SL g970 ( .A(n_886), .Y(n_970) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g1768 ( .A(n_890), .Y(n_1768) );
INVx1_ASAP7_75t_L g978 ( .A(n_891), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_917), .C(n_926), .Y(n_895) );
AND3x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .C(n_915), .Y(n_896) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_909), .A2(n_975), .B1(n_1224), .B2(n_1256), .Y(n_1255) );
INVx3_ASAP7_75t_L g1261 ( .A(n_909), .Y(n_1261) );
AND2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_922), .Y(n_917) );
INVx1_ASAP7_75t_L g1337 ( .A(n_919), .Y(n_1337) );
INVx1_ASAP7_75t_L g1459 ( .A(n_919), .Y(n_1459) );
OAI211xp5_ASAP7_75t_L g938 ( .A1(n_921), .A2(n_939), .B(n_941), .C(n_942), .Y(n_938) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_923), .A2(n_958), .B1(n_959), .B2(n_960), .Y(n_957) );
INVx2_ASAP7_75t_L g1339 ( .A(n_923), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_938), .C(n_943), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_931), .B(n_933), .C(n_936), .Y(n_929) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g1074 ( .A(n_932), .Y(n_1074) );
INVx2_ASAP7_75t_SL g1228 ( .A(n_932), .Y(n_1228) );
INVx1_ASAP7_75t_L g1740 ( .A(n_934), .Y(n_1740) );
BUFx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g949 ( .A(n_935), .Y(n_949) );
INVx2_ASAP7_75t_SL g1364 ( .A(n_937), .Y(n_1364) );
OAI211xp5_ASAP7_75t_L g1445 ( .A1(n_939), .A2(n_1446), .B(n_1447), .C(n_1448), .Y(n_1445) );
BUFx3_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g1455 ( .A(n_940), .Y(n_1455) );
XNOR2xp5_ASAP7_75t_L g951 ( .A(n_952), .B(n_1006), .Y(n_951) );
XNOR2x1_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .Y(n_952) );
AND2x2_ASAP7_75t_L g954 ( .A(n_955), .B(n_991), .Y(n_954) );
NOR3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_964), .C(n_966), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_957), .B(n_961), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B1(n_971), .B2(n_972), .Y(n_967) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_970), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_974), .A2(n_975), .B1(n_977), .B2(n_978), .Y(n_973) );
BUFx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
OAI22xp5_ASAP7_75t_SL g979 ( .A1(n_980), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_979) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND3xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_998), .C(n_1003), .Y(n_992) );
INVx1_ASAP7_75t_L g1244 ( .A(n_997), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1031), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1029), .B2(n_1030), .Y(n_1008) );
NAND3xp33_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1014), .C(n_1023), .Y(n_1010) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
NOR3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1040), .C(n_1042), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1037), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B1(n_1046), .B2(n_1048), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_1046), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
INVx2_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1051), .B1(n_1052), .B2(n_1053), .Y(n_1049) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
XNOR2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1329), .Y(n_1058) );
XOR2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1163), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1118), .B1(n_1119), .B2(n_1162), .Y(n_1060) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1061), .Y(n_1162) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
XNOR2x1_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1117), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1092), .Y(n_1063) );
INVx3_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
OAI211xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B(n_1075), .C(n_1076), .Y(n_1072) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NOR3xp33_ASAP7_75t_SL g1092 ( .A(n_1093), .B(n_1101), .C(n_1102), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1097), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_1104), .A2(n_1181), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1144), .Y(n_1121) );
NOR3xp33_ASAP7_75t_SL g1122 ( .A(n_1123), .B(n_1130), .C(n_1131), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1127), .Y(n_1123) );
NAND3xp33_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1153), .C(n_1160), .Y(n_1145) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
AOI22xp5_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1166), .B1(n_1277), .B2(n_1328), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
XNOR2xp5_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1216), .Y(n_1166) );
INVx2_ASAP7_75t_SL g1215 ( .A(n_1168), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1191), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1175), .B1(n_1177), .B2(n_1178), .Y(n_1171) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g1299 ( .A(n_1184), .Y(n_1299) );
AOI22xp5_ASAP7_75t_L g1749 ( .A1(n_1187), .A2(n_1750), .B1(n_1751), .B2(n_1753), .Y(n_1749) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1202), .Y(n_1191) );
INVx2_ASAP7_75t_L g1318 ( .A(n_1199), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1206), .Y(n_1202) );
INVx3_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_1212), .A2(n_1251), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
NAND4xp25_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1247), .C(n_1267), .D(n_1272), .Y(n_1217) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_1223), .A2(n_1250), .B1(n_1251), .B2(n_1252), .Y(n_1249) );
NAND3xp33_ASAP7_75t_SL g1231 ( .A(n_1232), .B(n_1236), .C(n_1243), .Y(n_1231) );
A2O1A1Ixp33_ASAP7_75t_L g1440 ( .A1(n_1233), .A2(n_1235), .B(n_1441), .C(n_1442), .Y(n_1440) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1291 ( .A(n_1239), .Y(n_1291) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1239), .Y(n_1382) );
INVx2_ASAP7_75t_L g1739 ( .A(n_1239), .Y(n_1739) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1259), .B1(n_1260), .B2(n_1262), .Y(n_1257) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1261), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1270), .Y(n_1267) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx2_ASAP7_75t_SL g1328 ( .A(n_1277), .Y(n_1328) );
XNOR2x1_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1279), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1309), .Y(n_1279) );
AOI31xp33_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1298), .A3(n_1305), .B(n_1308), .Y(n_1282) );
AOI211xp5_ASAP7_75t_SL g1283 ( .A1(n_1284), .A2(n_1285), .B(n_1287), .C(n_1288), .Y(n_1283) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
OAI21xp5_ASAP7_75t_SL g1289 ( .A1(n_1290), .A2(n_1292), .B(n_1293), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_1290), .A2(n_1345), .B1(n_1347), .B2(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
OAI221xp5_ASAP7_75t_L g1380 ( .A1(n_1295), .A2(n_1381), .B1(n_1382), .B2(n_1383), .C(n_1384), .Y(n_1380) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1301), .B2(n_1303), .C(n_1304), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1315), .Y(n_1309) );
NAND2xp5_ASAP7_75t_SL g1315 ( .A(n_1316), .B(n_1325), .Y(n_1315) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
XNOR2xp5_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1387), .Y(n_1330) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx2_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1334), .Y(n_1385) );
NAND3xp33_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1340), .C(n_1356), .Y(n_1334) );
NOR2xp33_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1338), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_1350), .A2(n_1354), .B1(n_1363), .B2(n_1365), .Y(n_1362) );
BUFx2_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
BUFx2_ASAP7_75t_SL g1365 ( .A(n_1366), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_1370), .A2(n_1372), .B1(n_1375), .B2(n_1380), .Y(n_1369) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
OAI221xp5_ASAP7_75t_L g1406 ( .A1(n_1377), .A2(n_1407), .B1(n_1408), .B2(n_1409), .C(n_1410), .Y(n_1406) );
INVxp67_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_1388), .A2(n_1433), .B1(n_1434), .B2(n_1474), .Y(n_1387) );
INVx1_ASAP7_75t_SL g1474 ( .A(n_1388), .Y(n_1474) );
XNOR2x1_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1390), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1414), .Y(n_1390) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
AOI31xp33_ASAP7_75t_SL g1736 ( .A1(n_1393), .A2(n_1737), .A3(n_1746), .B(n_1749), .Y(n_1736) );
INVx2_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
AOI211xp5_ASAP7_75t_L g1435 ( .A1(n_1394), .A2(n_1436), .B(n_1458), .C(n_1465), .Y(n_1435) );
NAND5xp2_ASAP7_75t_SL g1395 ( .A(n_1396), .B(n_1400), .C(n_1403), .D(n_1406), .E(n_1411), .Y(n_1395) );
OAI22xp33_ASAP7_75t_L g1430 ( .A1(n_1397), .A2(n_1401), .B1(n_1431), .B2(n_1432), .Y(n_1430) );
NOR3xp33_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1420), .C(n_1421), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1418), .Y(n_1415) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
NAND4xp25_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1440), .C(n_1445), .D(n_1452), .Y(n_1436) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
OAI211xp5_ASAP7_75t_L g1452 ( .A1(n_1453), .A2(n_1454), .B(n_1456), .C(n_1457), .Y(n_1452) );
INVx2_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1466), .B(n_1472), .Y(n_1465) );
OAI21xp5_ASAP7_75t_SL g1475 ( .A1(n_1476), .A2(n_1484), .B(n_1732), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx2_ASAP7_75t_L g1555 ( .A(n_1478), .Y(n_1555) );
OAI22xp5_ASAP7_75t_L g1634 ( .A1(n_1478), .A2(n_1635), .B1(n_1636), .B2(n_1637), .Y(n_1634) );
INVx2_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_SL g1523 ( .A(n_1479), .Y(n_1523) );
AND2x4_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1482), .Y(n_1479) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1480), .Y(n_1492) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1481), .B(n_1499), .Y(n_1498) );
AND2x4_ASAP7_75t_L g1491 ( .A(n_1482), .B(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1482), .B(n_1492), .Y(n_1514) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1483), .Y(n_1499) );
NOR3xp33_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1643), .C(n_1689), .Y(n_1484) );
AOI21xp5_ASAP7_75t_L g1485 ( .A1(n_1486), .A2(n_1594), .B(n_1633), .Y(n_1485) );
AOI221xp5_ASAP7_75t_L g1486 ( .A1(n_1487), .A2(n_1528), .B1(n_1544), .B2(n_1550), .C(n_1557), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g1487 ( .A(n_1488), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1503), .Y(n_1488) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1489), .Y(n_1615) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1489), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1662 ( .A(n_1489), .B(n_1646), .Y(n_1662) );
HB1xp67_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx2_ASAP7_75t_SL g1548 ( .A(n_1490), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1490), .B(n_1541), .Y(n_1592) );
OR2x2_ASAP7_75t_L g1599 ( .A(n_1490), .B(n_1541), .Y(n_1599) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1491), .Y(n_1538) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1491), .Y(n_1636) );
HB1xp67_ASAP7_75t_L g1790 ( .A(n_1492), .Y(n_1790) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_1494), .A2(n_1495), .B1(n_1500), .B2(n_1501), .Y(n_1493) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_1495), .A2(n_1501), .B1(n_1526), .B2(n_1527), .Y(n_1525) );
OAI22xp33_ASAP7_75t_L g1531 ( .A1(n_1495), .A2(n_1532), .B1(n_1533), .B2(n_1534), .Y(n_1531) );
BUFx3_ASAP7_75t_L g1640 ( .A(n_1495), .Y(n_1640) );
BUFx6f_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_1496), .A2(n_1501), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
OR2x2_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1498), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_1497), .B(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1497), .Y(n_1510) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1498), .Y(n_1509) );
HB1xp67_ASAP7_75t_L g1792 ( .A(n_1499), .Y(n_1792) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1501), .Y(n_1535) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1502), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1504), .B(n_1519), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1504), .B(n_1551), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1504), .B(n_1584), .Y(n_1629) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
NOR2xp33_ASAP7_75t_L g1576 ( .A(n_1505), .B(n_1561), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1505), .B(n_1519), .Y(n_1665) );
OR2x2_ASAP7_75t_L g1714 ( .A(n_1505), .B(n_1552), .Y(n_1714) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1515), .Y(n_1505) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1506), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1506), .B(n_1519), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1506), .B(n_1582), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1506), .B(n_1515), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1513), .Y(n_1506) );
AND2x4_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1510), .Y(n_1508) );
AND2x4_ASAP7_75t_L g1511 ( .A(n_1510), .B(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1514), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1515), .B(n_1551), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1515), .B(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1515), .Y(n_1582) );
NOR2xp33_ASAP7_75t_L g1695 ( .A(n_1515), .B(n_1556), .Y(n_1695) );
CKINVDCx6p67_ASAP7_75t_R g1556 ( .A(n_1519), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1519), .B(n_1576), .Y(n_1575) );
OAI331xp33_ASAP7_75t_L g1595 ( .A1(n_1519), .A2(n_1582), .A3(n_1596), .B1(n_1600), .B2(n_1603), .B3(n_1605), .C1(n_1607), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1519), .B(n_1581), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1648 ( .A(n_1519), .B(n_1563), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1519), .B(n_1564), .Y(n_1678) );
OR2x2_ASAP7_75t_L g1685 ( .A(n_1519), .B(n_1564), .Y(n_1685) );
OR2x6_ASAP7_75t_SL g1519 ( .A(n_1520), .B(n_1525), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1522), .B1(n_1523), .B2(n_1524), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1536 ( .A1(n_1523), .A2(n_1537), .B1(n_1538), .B2(n_1539), .Y(n_1536) );
XNOR2x1_ASAP7_75t_L g1734 ( .A(n_1524), .B(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1528), .Y(n_1618) );
A2O1A1Ixp33_ASAP7_75t_SL g1721 ( .A1(n_1528), .A2(n_1704), .B(n_1722), .C(n_1723), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1540), .Y(n_1528) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1529), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1529), .B(n_1571), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1609 ( .A(n_1529), .B(n_1541), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1529), .B(n_1541), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1529), .B(n_1592), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1529), .B(n_1548), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1680 ( .A(n_1529), .B(n_1633), .Y(n_1680) );
INVx3_ASAP7_75t_L g1709 ( .A(n_1529), .Y(n_1709) );
INVx3_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1530), .B(n_1541), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1530), .B(n_1552), .Y(n_1606) );
OR2x2_ASAP7_75t_L g1730 ( .A(n_1530), .B(n_1599), .Y(n_1730) );
OR2x2_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1536), .Y(n_1530) );
HB1xp67_ASAP7_75t_L g1642 ( .A(n_1534), .Y(n_1642) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
OAI211xp5_ASAP7_75t_SL g1557 ( .A1(n_1540), .A2(n_1558), .B(n_1565), .C(n_1587), .Y(n_1557) );
AOI22xp33_ASAP7_75t_SL g1698 ( .A1(n_1540), .A2(n_1664), .B1(n_1699), .B2(n_1703), .Y(n_1698) );
O2A1O1Ixp33_ASAP7_75t_L g1703 ( .A1(n_1540), .A2(n_1561), .B(n_1592), .C(n_1648), .Y(n_1703) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
OR2x2_ASAP7_75t_L g1547 ( .A(n_1541), .B(n_1548), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1541), .B(n_1548), .Y(n_1604) );
OAI22xp5_ASAP7_75t_L g1649 ( .A1(n_1541), .A2(n_1585), .B1(n_1650), .B2(n_1652), .Y(n_1649) );
AND2x4_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1543), .Y(n_1541) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1549), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_1546), .B(n_1647), .Y(n_1720) );
INVx2_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1711 ( .A(n_1547), .B(n_1647), .Y(n_1711) );
INVx2_ASAP7_75t_SL g1571 ( .A(n_1548), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1549), .B(n_1589), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1551), .B(n_1563), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1673 ( .A(n_1551), .B(n_1622), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1556), .Y(n_1551) );
INVx4_ASAP7_75t_L g1561 ( .A(n_1552), .Y(n_1561) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1552), .Y(n_1568) );
NOR2xp33_ASAP7_75t_L g1584 ( .A(n_1552), .B(n_1556), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1552), .B(n_1622), .Y(n_1654) );
OR2x2_ASAP7_75t_L g1664 ( .A(n_1552), .B(n_1665), .Y(n_1664) );
AOI322xp5_ASAP7_75t_L g1668 ( .A1(n_1552), .A2(n_1592), .A3(n_1598), .B1(n_1604), .B2(n_1669), .C1(n_1672), .C2(n_1674), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1552), .B(n_1604), .Y(n_1697) );
AND2x6_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1554), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1556), .B(n_1563), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1556), .B(n_1581), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1556), .B(n_1621), .Y(n_1620) );
NOR2xp33_ASAP7_75t_L g1653 ( .A(n_1556), .B(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1556), .B(n_1582), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1556), .B(n_1582), .Y(n_1725) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1562), .Y(n_1560) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1561), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1561), .B(n_1598), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1561), .B(n_1593), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1561), .B(n_1622), .Y(n_1621) );
NOR2xp33_ASAP7_75t_L g1701 ( .A(n_1561), .B(n_1702), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1562), .B(n_1589), .Y(n_1667) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1563), .Y(n_1602) );
OAI22xp5_ASAP7_75t_SL g1716 ( .A1(n_1564), .A2(n_1717), .B1(n_1718), .B2(n_1720), .Y(n_1716) );
AOI211xp5_ASAP7_75t_L g1565 ( .A1(n_1566), .A2(n_1570), .B(n_1573), .C(n_1577), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1568), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1568), .B(n_1688), .Y(n_1687) );
OAI32xp33_ASAP7_75t_L g1699 ( .A1(n_1568), .A2(n_1592), .A3(n_1648), .B1(n_1700), .B2(n_1701), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1572), .Y(n_1570) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1571), .Y(n_1574) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1571), .Y(n_1589) );
NOR2xp33_ASAP7_75t_L g1676 ( .A(n_1571), .B(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1571), .Y(n_1688) );
OAI22xp5_ASAP7_75t_L g1712 ( .A1(n_1571), .A2(n_1648), .B1(n_1713), .B2(n_1715), .Y(n_1712) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1571), .B(n_1714), .Y(n_1713) );
OAI21xp33_ASAP7_75t_L g1660 ( .A1(n_1572), .A2(n_1661), .B(n_1663), .Y(n_1660) );
NOR2xp33_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1575), .Y(n_1573) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1575), .Y(n_1657) );
AOI21xp33_ASAP7_75t_SL g1577 ( .A1(n_1578), .A2(n_1579), .B(n_1585), .Y(n_1577) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1578), .Y(n_1715) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1579), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1583), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1580), .B(n_1602), .Y(n_1601) );
NOR2xp33_ASAP7_75t_L g1623 ( .A(n_1580), .B(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
NOR3xp33_ASAP7_75t_L g1727 ( .A(n_1582), .B(n_1647), .C(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
OAI21xp5_ASAP7_75t_L g1587 ( .A1(n_1588), .A2(n_1590), .B(n_1593), .Y(n_1587) );
AOI221xp5_ASAP7_75t_SL g1675 ( .A1(n_1588), .A2(n_1676), .B1(n_1679), .B2(n_1681), .C(n_1682), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1593), .Y(n_1671) );
NOR5xp2_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1611), .C(n_1623), .D(n_1626), .E(n_1630), .Y(n_1594) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
A2O1A1Ixp33_ASAP7_75t_L g1731 ( .A1(n_1597), .A2(n_1630), .B(n_1695), .C(n_1709), .Y(n_1731) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
NOR2xp33_ASAP7_75t_L g1630 ( .A(n_1599), .B(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
NOR2x1_ASAP7_75t_R g1659 ( .A(n_1602), .B(n_1647), .Y(n_1659) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1604), .B(n_1628), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_1604), .B(n_1632), .Y(n_1692) );
INVxp67_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1610), .Y(n_1607) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
OAI22xp5_ASAP7_75t_SL g1611 ( .A1(n_1612), .A2(n_1614), .B1(n_1618), .B2(n_1619), .Y(n_1611) );
AOI21xp33_ASAP7_75t_L g1682 ( .A1(n_1612), .A2(n_1680), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1613), .B(n_1724), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1615), .B(n_1673), .Y(n_1717) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1650 ( .A(n_1617), .B(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
AOI21xp33_ASAP7_75t_L g1655 ( .A1(n_1624), .A2(n_1656), .B(n_1658), .Y(n_1655) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1633), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1708 ( .A(n_1633), .B(n_1709), .Y(n_1708) );
CKINVDCx5p33_ASAP7_75t_R g1728 ( .A(n_1633), .Y(n_1728) );
OR2x6_ASAP7_75t_SL g1633 ( .A(n_1634), .B(n_1638), .Y(n_1633) );
OAI22xp5_ASAP7_75t_L g1638 ( .A1(n_1639), .A2(n_1640), .B1(n_1641), .B2(n_1642), .Y(n_1638) );
NAND4xp25_ASAP7_75t_L g1643 ( .A(n_1644), .B(n_1660), .C(n_1668), .D(n_1675), .Y(n_1643) );
AOI211xp5_ASAP7_75t_SL g1644 ( .A1(n_1645), .A2(n_1646), .B(n_1649), .C(n_1655), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1648), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1647), .B(n_1678), .Y(n_1677) );
NOR2x1_ASAP7_75t_L g1724 ( .A(n_1647), .B(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1648), .Y(n_1670) );
OAI31xp33_ASAP7_75t_L g1726 ( .A1(n_1648), .A2(n_1674), .A3(n_1727), .B(n_1729), .Y(n_1726) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1654), .Y(n_1722) );
INVxp67_ASAP7_75t_SL g1656 ( .A(n_1657), .Y(n_1656) );
INVxp33_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
NAND2xp33_ASAP7_75t_L g1663 ( .A(n_1664), .B(n_1666), .Y(n_1663) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1664), .Y(n_1674) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1665), .Y(n_1719) );
INVxp33_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1671), .Y(n_1669) );
NOR2xp33_ASAP7_75t_L g1718 ( .A(n_1672), .B(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
AOI22xp5_ASAP7_75t_L g1706 ( .A1(n_1679), .A2(n_1707), .B1(n_1710), .B2(n_1716), .Y(n_1706) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1686), .Y(n_1683) );
OAI21xp5_ASAP7_75t_SL g1710 ( .A1(n_1684), .A2(n_1711), .B(n_1712), .Y(n_1710) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
NAND5xp2_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1706), .C(n_1721), .D(n_1726), .E(n_1731), .Y(n_1689) );
OAI31xp33_ASAP7_75t_SL g1690 ( .A1(n_1691), .A2(n_1693), .A3(n_1698), .B(n_1704), .Y(n_1690) );
INVxp67_ASAP7_75t_SL g1691 ( .A(n_1692), .Y(n_1691) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1696), .Y(n_1693) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1700), .Y(n_1702) );
CKINVDCx14_ASAP7_75t_R g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1735), .Y(n_1781) );
OR2x2_ASAP7_75t_L g1735 ( .A(n_1736), .B(n_1754), .Y(n_1735) );
NAND3xp33_ASAP7_75t_L g1754 ( .A(n_1755), .B(n_1766), .C(n_1774), .Y(n_1754) );
INVxp67_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
BUFx2_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
INVxp67_ASAP7_75t_SL g1779 ( .A(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
CKINVDCx5p33_ASAP7_75t_R g1784 ( .A(n_1785), .Y(n_1784) );
A2O1A1Ixp33_ASAP7_75t_L g1788 ( .A1(n_1786), .A2(n_1789), .B(n_1791), .C(n_1793), .Y(n_1788) );
HB1xp67_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
endmodule