module real_jpeg_25142_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_82),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_49),
.C(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_7),
.B(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_54),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_10),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_23),
.B1(n_49),
.B2(n_50),
.Y(n_130)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_13),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_99),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_97),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_88),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_17),
.B(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_58),
.B2(n_59),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_22),
.A2(n_28),
.B1(n_62),
.B2(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_26),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_24),
.B(n_63),
.CON(n_62),
.SN(n_62)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_31),
.C(n_34),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_32),
.B(n_62),
.C(n_64),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_31),
.A2(n_32),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_32),
.B(n_104),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_46),
.B2(n_57),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B(n_53),
.Y(n_46)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_52),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_50),
.B1(n_76),
.B2(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_50),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_51),
.A2(n_69),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_54),
.A2(n_123),
.B1(n_130),
.B2(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_73),
.B1(n_86),
.B2(n_87),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_90),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_63),
.B(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B(n_70),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_80),
.B(n_83),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_79),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_79),
.B1(n_95),
.B2(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_85),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.C(n_93),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_93),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_144),
.B(n_148),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_119),
.B(n_143),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_114),
.C(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_127),
.B(n_142),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_125),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_138),
.B(n_141),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);


endmodule