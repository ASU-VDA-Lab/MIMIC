module real_jpeg_6586_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_0),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_0),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_0),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_0),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_0),
.B(n_34),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_1),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_2),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_2),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_2),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_2),
.B(n_235),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_2),
.B(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_3),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_3),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_4),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_5),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_5),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_5),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_5),
.B(n_420),
.Y(n_419)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_6),
.Y(n_152)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_7),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_8),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_8),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_8),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_8),
.B(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_9),
.Y(n_222)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_9),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_9),
.Y(n_308)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_11),
.Y(n_240)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_11),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_12),
.B(n_41),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_12),
.B(n_48),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_12),
.B(n_221),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_12),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_242),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_12),
.B(n_139),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_12),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_12),
.B(n_99),
.Y(n_460)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_14),
.B(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_14),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_14),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_14),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_15),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_15),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_15),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_15),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_15),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_15),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_15),
.B(n_202),
.Y(n_363)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_17),
.B(n_31),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_17),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_17),
.B(n_155),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_17),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_17),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_17),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_17),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_18),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_18),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_18),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_18),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_19),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_19),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_19),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_19),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_19),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_19),
.B(n_221),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_19),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_19),
.B(n_436),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_502),
.B(n_504),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_163),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_162),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_142),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_24),
.B(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_103),
.C(n_114),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_25),
.B(n_488),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_71),
.C(n_85),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_26),
.B(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.C(n_56),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_27),
.B(n_46),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_28),
.B(n_38),
.C(n_45),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_29),
.B(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_31),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_35),
.Y(n_217)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_37),
.Y(n_329)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_43),
.Y(n_324)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_44),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_44),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.C(n_53),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_47),
.B(n_53),
.Y(n_451)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_51),
.B(n_451),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_56),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_63),
.C(n_70),
.Y(n_112)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_60),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_61),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_61),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_64),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_106),
.C(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_88),
.C(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_65),
.A2(n_70),
.B1(n_88),
.B2(n_89),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_69),
.Y(n_282)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_69),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_71),
.A2(n_85),
.B1(n_86),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_71),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_77),
.C(n_80),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_95),
.C(n_100),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_87),
.B(n_478),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_88),
.A2(n_89),
.B1(n_431),
.B2(n_433),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_88),
.B(n_431),
.C(n_434),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_91),
.B(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_478)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_100),
.A2(n_101),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_101),
.B(n_461),
.C(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_103),
.B(n_114),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.C(n_113),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_104),
.B(n_494),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_107),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_124),
.C(n_129),
.Y(n_159)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_108),
.Y(n_295)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_112),
.B(n_113),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_132),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_130),
.B2(n_131),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_131),
.C(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_123),
.B2(n_129),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_125),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_137),
.C(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_157),
.B2(n_158),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

AO21x1_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_483),
.B(n_499),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_466),
.B(n_482),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_440),
.B(n_465),
.Y(n_165)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_397),
.B(n_439),
.Y(n_166)
);

AOI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_356),
.B(n_396),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_275),
.B(n_355),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_260),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_170),
.B(n_260),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_211),
.B2(n_259),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_171),
.B(n_212),
.C(n_243),
.Y(n_395)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_188),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_173),
.B(n_189),
.C(n_210),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.C(n_187),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_174),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_187),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_198),
.B1(n_209),
.B2(n_210),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B(n_197),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_193),
.Y(n_197)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_197),
.B(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_197),
.B(n_361),
.C(n_374),
.Y(n_404)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_199),
.B(n_204),
.C(n_207),
.Y(n_394)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_243),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_224),
.C(n_236),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_218),
.C(n_223),
.Y(n_258)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_222),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_225),
.B1(n_236),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_233),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_226),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_348)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_228),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_231),
.Y(n_383)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_241),
.Y(n_257)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g432 ( 
.A(n_240),
.Y(n_432)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

XOR2x1_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_256),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_244),
.B(n_257),
.C(n_258),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_245),
.B(n_250),
.C(n_254),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_250),
.B1(n_254),
.B2(n_255),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_249),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_253),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.C(n_273),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_261),
.B(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_264),
.B(n_273),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_266),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_267),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_271),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_350),
.B(n_354),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_335),
.B(n_349),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_315),
.B(n_334),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_302),
.B(n_314),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_296),
.B2(n_297),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_293),
.C(n_296),
.Y(n_333)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g411 ( 
.A(n_292),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_301),
.Y(n_319)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_309),
.B(n_313),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_333),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_333),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_319),
.C(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_330),
.C(n_332),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVx11_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_325)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_338),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_345),
.C(n_346),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_352),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_395),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_395),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_376),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_360),
.C(n_376),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_373),
.B2(n_375),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_366),
.C(n_368),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_368),
.B2(n_369),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_379),
.C(n_389),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_389),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_385),
.C(n_386),
.Y(n_427)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_393),
.C(n_394),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_399),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_417),
.C(n_437),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_417),
.B1(n_437),
.B2(n_438),
.Y(n_401)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_405),
.B2(n_416),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_406),
.C(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_415),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_412),
.C(n_415),
.Y(n_457)
);

INVx8_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx6_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_426),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_427),
.C(n_428),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g509 ( 
.A(n_418),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_422),
.CI(n_425),
.CON(n_418),
.SN(n_418)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_422),
.C(n_425),
.Y(n_462)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_434),
.B2(n_435),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_431),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_464),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_464),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_442),
.B(n_444),
.C(n_453),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_453),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_452),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_449),
.C(n_450),
.Y(n_472)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_448),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_456),
.B2(n_463),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_457),
.C(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_456),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_460),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_481),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_481),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_470),
.C(n_479),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_479),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_475),
.C(n_477),
.Y(n_495)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.Y(n_474)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_496),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_500),
.B(n_501),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_489),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.C(n_495),
.Y(n_489)
);

FAx1_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_493),
.CI(n_495),
.CON(n_497),
.SN(n_497)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_498),
.Y(n_500)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_497),
.Y(n_507)
);

INVx13_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx8_ASAP7_75t_L g505 ( 
.A(n_503),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);


endmodule