module real_aes_18436_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_840, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_840;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g114 ( .A(n_0), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_1), .A2(n_4), .B1(n_142), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_2), .A2(n_42), .B1(n_149), .B2(n_185), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_3), .A2(n_24), .B1(n_185), .B2(n_227), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_5), .A2(n_16), .B1(n_139), .B2(n_216), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_6), .A2(n_62), .B1(n_199), .B2(n_229), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_7), .A2(n_17), .B1(n_149), .B2(n_170), .Y(n_620) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_9), .A2(n_473), .B(n_829), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_10), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_11), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_12), .A2(n_18), .B1(n_198), .B2(n_201), .Y(n_197) );
OR2x2_ASAP7_75t_L g110 ( .A(n_13), .B(n_37), .Y(n_110) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_15), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_19), .A2(n_101), .B1(n_139), .B2(n_142), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_20), .A2(n_38), .B1(n_174), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_21), .B(n_140), .Y(n_171) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_22), .A2(n_57), .B(n_158), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_23), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_25), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_26), .B(n_146), .Y(n_540) );
INVx4_ASAP7_75t_R g588 ( .A(n_27), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_28), .A2(n_47), .B1(n_187), .B2(n_188), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_29), .A2(n_54), .B1(n_139), .B2(n_188), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_30), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_31), .B(n_174), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_32), .Y(n_250) );
INVx1_ASAP7_75t_L g519 ( .A(n_33), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_34), .B(n_185), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_SL g531 ( .A1(n_35), .A2(n_145), .B(n_149), .C(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_36), .A2(n_55), .B1(n_149), .B2(n_188), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_39), .A2(n_88), .B1(n_149), .B2(n_226), .Y(n_225) );
XOR2x2_ASAP7_75t_L g822 ( .A(n_40), .B(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_41), .A2(n_45), .B1(n_149), .B2(n_170), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_43), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_44), .A2(n_60), .B1(n_139), .B2(n_148), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_46), .A2(n_74), .B1(n_824), .B2(n_825), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_46), .Y(n_825) );
INVx1_ASAP7_75t_L g543 ( .A(n_48), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_49), .B(n_149), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_50), .Y(n_560) );
INVx2_ASAP7_75t_L g481 ( .A(n_51), .Y(n_481) );
BUFx3_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g467 ( .A(n_52), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_53), .A2(n_118), .B(n_469), .Y(n_117) );
AOI31xp33_ASAP7_75t_L g469 ( .A1(n_53), .A2(n_470), .A3(n_472), .B(n_473), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_56), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_58), .A2(n_89), .B1(n_149), .B2(n_188), .Y(n_621) );
INVx1_ASAP7_75t_L g836 ( .A(n_59), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_61), .A2(n_69), .B1(n_121), .B2(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_63), .A2(n_77), .B1(n_148), .B2(n_187), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_64), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_65), .A2(n_79), .B1(n_149), .B2(n_170), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_66), .A2(n_100), .B1(n_139), .B2(n_201), .Y(n_247) );
AND2x4_ASAP7_75t_L g135 ( .A(n_67), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g158 ( .A(n_68), .Y(n_158) );
INVx1_ASAP7_75t_L g121 ( .A(n_69), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_70), .A2(n_92), .B1(n_187), .B2(n_188), .Y(n_515) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_71), .A2(n_78), .B1(n_213), .B2(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g136 ( .A(n_72), .Y(n_136) );
AND2x2_ASAP7_75t_L g535 ( .A(n_73), .B(n_180), .Y(n_535) );
INVx1_ASAP7_75t_L g824 ( .A(n_74), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_75), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_76), .B(n_229), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_80), .B(n_185), .Y(n_561) );
INVx2_ASAP7_75t_L g146 ( .A(n_81), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_82), .B(n_180), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_83), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_84), .A2(n_99), .B1(n_188), .B2(n_229), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_85), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_86), .B(n_156), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_87), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_90), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_91), .B(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_93), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_94), .B(n_180), .Y(n_557) );
INVx1_ASAP7_75t_L g113 ( .A(n_95), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_95), .B(n_466), .Y(n_465) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_96), .B(n_140), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_97), .A2(n_204), .B(n_229), .C(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g590 ( .A(n_98), .B(n_591), .Y(n_590) );
NAND2xp33_ASAP7_75t_L g565 ( .A(n_102), .B(n_175), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_116), .B(n_835), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx6f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx12f_ASAP7_75t_L g838 ( .A(n_106), .Y(n_838) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g834 ( .A(n_108), .B(n_495), .Y(n_834) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g489 ( .A(n_109), .Y(n_489) );
INVx1_ASAP7_75t_L g468 ( .A(n_110), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g495 ( .A(n_113), .Y(n_495) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_477), .B(n_482), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_462), .Y(n_118) );
INVx1_ASAP7_75t_L g472 ( .A(n_119), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx2_ASAP7_75t_L g496 ( .A(n_123), .Y(n_496) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_365), .Y(n_123) );
NAND4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_289), .C(n_320), .D(n_349), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_256), .Y(n_125) );
OAI322xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_192), .A3(n_221), .B1(n_234), .B2(n_242), .C1(n_251), .C2(n_253), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_128), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_162), .Y(n_128) );
AND2x2_ASAP7_75t_L g286 ( .A(n_129), .B(n_287), .Y(n_286) );
INVx4_ASAP7_75t_L g322 ( .A(n_129), .Y(n_322) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g297 ( .A(n_130), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g300 ( .A(n_130), .B(n_194), .Y(n_300) );
AND2x2_ASAP7_75t_L g317 ( .A(n_130), .B(n_210), .Y(n_317) );
AND2x2_ASAP7_75t_L g415 ( .A(n_130), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g238 ( .A(n_131), .Y(n_238) );
AND2x4_ASAP7_75t_L g421 ( .A(n_131), .B(n_416), .Y(n_421) );
AO31x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .A3(n_153), .B(n_159), .Y(n_131) );
AO31x2_ASAP7_75t_L g245 ( .A1(n_132), .A2(n_205), .A3(n_246), .B(n_249), .Y(n_245) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_133), .A2(n_583), .B(n_586), .Y(n_582) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AO31x2_ASAP7_75t_L g182 ( .A1(n_134), .A2(n_183), .A3(n_189), .B(n_190), .Y(n_182) );
AO31x2_ASAP7_75t_L g195 ( .A1(n_134), .A2(n_196), .A3(n_205), .B(n_207), .Y(n_195) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_134), .A2(n_211), .A3(n_218), .B(n_219), .Y(n_210) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_134), .A2(n_161), .A3(n_619), .B(n_622), .Y(n_618) );
BUFx10_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
BUFx10_ASAP7_75t_L g510 ( .A(n_135), .Y(n_510) );
INVx1_ASAP7_75t_L g534 ( .A(n_135), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B1(n_147), .B2(n_150), .Y(n_137) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_140), .Y(n_578) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g143 ( .A(n_141), .Y(n_143) );
INVx3_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx1_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
INVx1_ASAP7_75t_L g214 ( .A(n_141), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
INVx2_ASAP7_75t_L g227 ( .A(n_141), .Y(n_227) );
INVx1_ASAP7_75t_L g229 ( .A(n_141), .Y(n_229) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_143), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_144), .A2(n_173), .B(n_176), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_144), .A2(n_150), .B1(n_184), .B2(n_186), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_144), .A2(n_197), .B1(n_202), .B2(n_203), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_144), .A2(n_150), .B1(n_212), .B2(n_215), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_144), .A2(n_225), .B1(n_228), .B2(n_230), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_144), .A2(n_203), .B1(n_247), .B2(n_248), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_144), .A2(n_150), .B1(n_266), .B2(n_267), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_144), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_144), .A2(n_230), .B1(n_515), .B2(n_516), .Y(n_514) );
OAI22x1_ASAP7_75t_L g619 ( .A1(n_144), .A2(n_230), .B1(n_620), .B2(n_621), .Y(n_619) );
INVx6_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
O2A1O1Ixp5_ASAP7_75t_L g168 ( .A1(n_145), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_145), .A2(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_145), .B(n_577), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_145), .A2(n_573), .B(n_577), .C(n_580), .Y(n_634) );
BUFx8_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
INVx1_ASAP7_75t_L g530 ( .A(n_146), .Y(n_530) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
INVx1_ASAP7_75t_L g201 ( .A(n_149), .Y(n_201) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g509 ( .A(n_151), .Y(n_509) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g563 ( .A(n_152), .Y(n_563) );
AO31x2_ASAP7_75t_L g264 ( .A1(n_153), .A2(n_231), .A3(n_265), .B(n_268), .Y(n_264) );
AO21x2_ASAP7_75t_L g581 ( .A1(n_153), .A2(n_582), .B(n_590), .Y(n_581) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_SL g207 ( .A(n_155), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_155), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
INVx2_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
OAI21xp33_ASAP7_75t_L g580 ( .A1(n_156), .A2(n_534), .B(n_575), .Y(n_580) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_157), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_161), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g426 ( .A(n_162), .B(n_327), .Y(n_426) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g255 ( .A(n_163), .Y(n_255) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_163), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_181), .Y(n_163) );
AND2x2_ASAP7_75t_L g243 ( .A(n_164), .B(n_182), .Y(n_243) );
INVx1_ASAP7_75t_L g284 ( .A(n_164), .Y(n_284) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_179), .Y(n_164) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_165), .A2(n_167), .B(n_179), .Y(n_279) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_166), .B(n_191), .Y(n_190) );
BUFx3_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_166), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_166), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g547 ( .A(n_166), .B(n_510), .Y(n_547) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_172), .B(n_177), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_170), .A2(n_560), .B(n_561), .C(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g187 ( .A(n_175), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_175), .A2(n_217), .B1(n_588), .B2(n_589), .Y(n_587) );
INVx2_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_SL g231 ( .A(n_178), .Y(n_231) );
INVx2_ASAP7_75t_L g189 ( .A(n_180), .Y(n_189) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_180), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g275 ( .A(n_181), .Y(n_275) );
AND2x2_ASAP7_75t_L g339 ( .A(n_181), .B(n_278), .Y(n_339) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g293 ( .A(n_182), .Y(n_293) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_182), .Y(n_346) );
OR2x2_ASAP7_75t_L g417 ( .A(n_182), .B(n_223), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_185), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g517 ( .A(n_188), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_188), .B(n_542), .Y(n_541) );
AO31x2_ASAP7_75t_L g505 ( .A1(n_189), .A2(n_506), .A3(n_510), .B(n_511), .Y(n_505) );
NAND4xp25_ASAP7_75t_L g295 ( .A(n_192), .B(n_296), .C(n_299), .D(n_301), .Y(n_295) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g433 ( .A(n_193), .B(n_421), .Y(n_433) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_209), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_194), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g287 ( .A(n_194), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g307 ( .A(n_194), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_194), .Y(n_324) );
INVx1_ASAP7_75t_L g332 ( .A(n_194), .Y(n_332) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_194), .Y(n_446) );
INVx4_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_195), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g364 ( .A(n_195), .B(n_264), .Y(n_364) );
AND2x2_ASAP7_75t_L g372 ( .A(n_195), .B(n_210), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_195), .B(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g437 ( .A(n_195), .Y(n_437) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_200), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g230 ( .A(n_204), .Y(n_230) );
AO31x2_ASAP7_75t_L g513 ( .A1(n_205), .A2(n_231), .A3(n_514), .B(n_518), .Y(n_513) );
AOI21x1_ASAP7_75t_L g522 ( .A1(n_205), .A2(n_523), .B(n_535), .Y(n_522) );
BUFx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_206), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_206), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g591 ( .A(n_206), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_206), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
OR2x2_ASAP7_75t_L g302 ( .A(n_210), .B(n_264), .Y(n_302) );
INVx2_ASAP7_75t_L g309 ( .A(n_210), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_210), .B(n_262), .Y(n_333) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_210), .Y(n_420) );
OAI21xp33_ASAP7_75t_SL g539 ( .A1(n_213), .A2(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_218), .A2(n_224), .A3(n_231), .B(n_232), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_221), .B(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g244 ( .A(n_223), .B(n_245), .Y(n_244) );
BUFx2_ASAP7_75t_L g254 ( .A(n_223), .Y(n_254) );
INVx2_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
AND2x4_ASAP7_75t_L g304 ( .A(n_223), .B(n_276), .Y(n_304) );
OR2x2_ASAP7_75t_L g384 ( .A(n_223), .B(n_284), .Y(n_384) );
INVx2_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_227), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_230), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_239), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_236), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g301 ( .A(n_236), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_236), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_237), .B(n_307), .Y(n_315) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
OR2x2_ASAP7_75t_L g353 ( .A(n_238), .B(n_263), .Y(n_353) );
INVx1_ASAP7_75t_L g280 ( .A(n_239), .Y(n_280) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g252 ( .A(n_240), .Y(n_252) );
INVx1_ASAP7_75t_L g288 ( .A(n_241), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
OAI322xp33_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_257), .A3(n_270), .B1(n_273), .B2(n_280), .C1(n_281), .C2(n_285), .Y(n_256) );
AND2x4_ASAP7_75t_L g303 ( .A(n_243), .B(n_304), .Y(n_303) );
AOI211xp5_ASAP7_75t_SL g334 ( .A1(n_243), .A2(n_335), .B(n_336), .C(n_340), .Y(n_334) );
AND2x2_ASAP7_75t_L g354 ( .A(n_243), .B(n_244), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_243), .B(n_271), .Y(n_360) );
AND2x4_ASAP7_75t_SL g282 ( .A(n_244), .B(n_283), .Y(n_282) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_244), .B(n_300), .C(n_328), .Y(n_373) );
AND2x2_ASAP7_75t_L g404 ( .A(n_244), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g271 ( .A(n_245), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
BUFx2_ASAP7_75t_L g344 ( .A(n_245), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_254), .B(n_278), .Y(n_277) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_254), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g337 ( .A(n_254), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_255), .B(n_271), .Y(n_402) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g345 ( .A(n_260), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_264), .Y(n_298) );
AND2x4_ASAP7_75t_L g308 ( .A(n_264), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g395 ( .A(n_264), .Y(n_395) );
INVx2_ASAP7_75t_L g416 ( .A(n_264), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_270), .A2(n_429), .B1(n_431), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g340 ( .A(n_271), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g294 ( .A(n_272), .B(n_278), .Y(n_294) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g313 ( .A(n_274), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x4_ASAP7_75t_L g283 ( .A(n_275), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g405 ( .A(n_275), .Y(n_405) );
INVx2_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
AND2x2_ASAP7_75t_L g319 ( .A(n_276), .B(n_278), .Y(n_319) );
INVx3_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_276), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx2_ASAP7_75t_L g328 ( .A(n_279), .Y(n_328) );
OAI222xp33_ASAP7_75t_L g451 ( .A1(n_281), .A2(n_441), .B1(n_452), .B2(n_455), .C1(n_457), .C2(n_459), .Y(n_451) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g392 ( .A(n_283), .Y(n_392) );
AND2x2_ASAP7_75t_L g456 ( .A(n_283), .B(n_326), .Y(n_456) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_286), .B(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .B1(n_303), .B2(n_305), .C(n_310), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
INVx2_ASAP7_75t_L g440 ( .A(n_292), .Y(n_440) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g341 ( .A(n_293), .Y(n_341) );
AND2x2_ASAP7_75t_L g377 ( .A(n_293), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g343 ( .A(n_294), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g458 ( .A(n_294), .Y(n_458) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g430 ( .A(n_300), .B(n_308), .Y(n_430) );
AND2x2_ASAP7_75t_L g453 ( .A(n_300), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g314 ( .A(n_302), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g449 ( .A(n_302), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_303), .A2(n_357), .B1(n_391), .B2(n_393), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_303), .A2(n_419), .B(n_422), .Y(n_418) );
INVxp67_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx2_ASAP7_75t_SL g439 ( .A(n_304), .Y(n_439) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
OR2x2_ASAP7_75t_L g352 ( .A(n_306), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g450 ( .A(n_306), .B(n_449), .Y(n_450) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g323 ( .A(n_308), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_308), .B(n_332), .Y(n_348) );
INVx2_ASAP7_75t_L g375 ( .A(n_308), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B1(n_316), .B2(n_318), .Y(n_310) );
NOR2xp33_ASAP7_75t_SL g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_312), .A2(n_386), .B1(n_399), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g408 ( .A(n_317), .B(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_325), .B(n_329), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g389 ( .A(n_322), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_322), .B(n_372), .Y(n_400) );
INVx1_ASAP7_75t_L g358 ( .A(n_324), .Y(n_358) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_326), .B(n_339), .Y(n_431) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_327), .A2(n_445), .B(n_447), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_334), .B(n_342), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g388 ( .A(n_333), .Y(n_388) );
INVx1_ASAP7_75t_L g454 ( .A(n_333), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g427 ( .A(n_337), .Y(n_427) );
OR2x2_ASAP7_75t_L g438 ( .A(n_338), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .C(n_347), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_343), .A2(n_404), .B1(n_406), .B2(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_345), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_348), .B(n_352), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_348), .A2(n_411), .B1(n_414), .B2(n_417), .C(n_418), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B(n_355), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g359 ( .A(n_353), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B1(n_361), .B2(n_840), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g442 ( .A(n_364), .B(n_420), .Y(n_442) );
NAND4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_396), .C(n_423), .D(n_443), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_379), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_373), .B2(n_374), .C(n_376), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_369), .A2(n_426), .B1(n_448), .B2(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_372), .B(n_415), .Y(n_414) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_372), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_374), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g381 ( .A(n_378), .B(n_382), .Y(n_381) );
OAI21xp33_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_385), .B(n_390), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g409 ( .A(n_395), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_395), .A2(n_424), .B(n_428), .C(n_434), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_410), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_403), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g457 ( .A(n_405), .B(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx3_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI22xp33_ASAP7_75t_R g434 ( .A1(n_435), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g448 ( .A(n_437), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_451), .Y(n_443) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx5_ASAP7_75t_L g471 ( .A(n_464), .Y(n_471) );
INVx5_ASAP7_75t_L g476 ( .A(n_464), .Y(n_476) );
AND2x6_ASAP7_75t_SL g464 ( .A(n_465), .B(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_468), .B(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx8_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g487 ( .A(n_481), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_481), .B(n_833), .Y(n_832) );
OAI321xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_490), .A3(n_821), .B1(n_826), .B2(n_827), .C(n_828), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_484), .B(n_821), .Y(n_827) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx6_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x6_ASAP7_75t_SL g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g826 ( .A(n_490), .Y(n_826) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_494), .Y(n_497) );
BUFx8_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_713), .Y(n_498) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_500), .B(n_655), .Y(n_499) );
NAND3xp33_ASAP7_75t_SL g500 ( .A(n_501), .B(n_592), .C(n_637), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_548), .B(n_569), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_502), .A2(n_593), .B1(n_612), .B2(n_624), .Y(n_592) );
AOI22x1_ASAP7_75t_L g717 ( .A1(n_502), .A2(n_718), .B1(n_722), .B2(n_723), .Y(n_717) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_520), .Y(n_503) );
OR2x2_ASAP7_75t_L g678 ( .A(n_504), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
OR2x2_ASAP7_75t_L g553 ( .A(n_505), .B(n_513), .Y(n_553) );
AND2x2_ASAP7_75t_L g596 ( .A(n_505), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_SL g604 ( .A(n_505), .Y(n_604) );
BUFx2_ASAP7_75t_L g654 ( .A(n_505), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_509), .A2(n_545), .B(n_546), .Y(n_544) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_509), .A2(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g568 ( .A(n_510), .Y(n_568) );
AND2x2_ASAP7_75t_L g599 ( .A(n_513), .B(n_536), .Y(n_599) );
INVx1_ASAP7_75t_L g606 ( .A(n_513), .Y(n_606) );
INVx1_ASAP7_75t_L g611 ( .A(n_513), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_513), .B(n_604), .Y(n_673) );
INVx1_ASAP7_75t_L g694 ( .A(n_513), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_513), .B(n_597), .Y(n_764) );
INVx1_ASAP7_75t_L g657 ( .A(n_520), .Y(n_657) );
OR2x2_ASAP7_75t_L g709 ( .A(n_520), .B(n_673), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_536), .Y(n_520) );
AND2x2_ASAP7_75t_L g554 ( .A(n_521), .B(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g602 ( .A(n_521), .B(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_521), .B(n_551), .Y(n_685) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_531), .B(n_534), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_527), .B(n_529), .Y(n_524) );
BUFx4f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_530), .B(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g551 ( .A(n_536), .Y(n_551) );
INVx1_ASAP7_75t_L g651 ( .A(n_536), .Y(n_651) );
AND2x2_ASAP7_75t_L g653 ( .A(n_536), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g671 ( .A(n_536), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g693 ( .A(n_536), .B(n_694), .Y(n_693) );
NAND2x1p5_ASAP7_75t_SL g704 ( .A(n_536), .B(n_680), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_536), .B(n_611), .Y(n_794) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_544), .B(n_547), .Y(n_538) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_554), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_549), .A2(n_733), .B1(n_734), .B2(n_736), .Y(n_732) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_550), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_550), .B(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g811 ( .A(n_550), .B(n_669), .Y(n_811) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g610 ( .A(n_551), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_551), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g699 ( .A(n_551), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g650 ( .A(n_552), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g740 ( .A(n_553), .Y(n_740) );
OR2x2_ASAP7_75t_L g814 ( .A(n_553), .B(n_741), .Y(n_814) );
INVx1_ASAP7_75t_L g645 ( .A(n_554), .Y(n_645) );
INVx3_ASAP7_75t_L g649 ( .A(n_555), .Y(n_649) );
BUFx2_ASAP7_75t_L g660 ( .A(n_555), .Y(n_660) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g630 ( .A(n_556), .B(n_581), .Y(n_630) );
INVx2_ASAP7_75t_L g676 ( .A(n_556), .Y(n_676) );
INVx1_ASAP7_75t_L g708 ( .A(n_556), .Y(n_708) );
AND2x2_ASAP7_75t_L g721 ( .A(n_556), .B(n_618), .Y(n_721) );
AND2x2_ASAP7_75t_L g743 ( .A(n_556), .B(n_642), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .B(n_567), .Y(n_558) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g734 ( .A(n_570), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_570), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g759 ( .A(n_570), .B(n_627), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_570), .B(n_761), .Y(n_760) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_581), .Y(n_570) );
INVx2_ASAP7_75t_L g616 ( .A(n_571), .Y(n_616) );
AND2x2_ASAP7_75t_L g643 ( .A(n_571), .B(n_644), .Y(n_643) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_579), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g617 ( .A(n_581), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g636 ( .A(n_581), .Y(n_636) );
INVx2_ASAP7_75t_L g644 ( .A(n_581), .Y(n_644) );
OR2x2_ASAP7_75t_L g664 ( .A(n_581), .B(n_618), .Y(n_664) );
AND2x2_ASAP7_75t_L g675 ( .A(n_581), .B(n_676), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_600), .B2(n_605), .C(n_607), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI32xp33_ASAP7_75t_L g705 ( .A1(n_595), .A2(n_609), .A3(n_706), .B1(n_709), .B2(n_710), .Y(n_705) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g695 ( .A(n_596), .Y(n_695) );
AND2x2_ASAP7_75t_L g731 ( .A(n_596), .B(n_610), .Y(n_731) );
INVx1_ASAP7_75t_L g795 ( .A(n_596), .Y(n_795) );
OR2x2_ASAP7_75t_L g669 ( .A(n_597), .B(n_604), .Y(n_669) );
INVx2_ASAP7_75t_L g680 ( .A(n_597), .Y(n_680) );
BUFx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g819 ( .A(n_599), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_L g806 ( .A(n_602), .Y(n_806) );
INVx1_ASAP7_75t_L g820 ( .A(n_602), .Y(n_820) );
OR2x2_ASAP7_75t_L g700 ( .A(n_603), .B(n_680), .Y(n_700) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_605), .B(n_700), .Y(n_722) );
INVx1_ASAP7_75t_L g753 ( .A(n_605), .Y(n_753) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g787 ( .A(n_606), .Y(n_787) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2x1_ASAP7_75t_L g756 ( .A(n_608), .B(n_757), .Y(n_756) );
OAI21xp5_ASAP7_75t_SL g778 ( .A1(n_609), .A2(n_779), .B(n_784), .Y(n_778) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
AND2x2_ASAP7_75t_L g688 ( .A(n_614), .B(n_630), .Y(n_688) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_614), .Y(n_818) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g720 ( .A(n_615), .Y(n_720) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g702 ( .A(n_616), .B(n_676), .Y(n_702) );
AND2x2_ASAP7_75t_L g773 ( .A(n_616), .B(n_644), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_617), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g701 ( .A(n_617), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g780 ( .A(n_617), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g629 ( .A(n_618), .Y(n_629) );
INVx2_ASAP7_75t_L g642 ( .A(n_618), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_618), .B(n_633), .Y(n_690) );
AND2x2_ASAP7_75t_L g750 ( .A(n_618), .B(n_644), .Y(n_750) );
NAND2xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_631), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g725 ( .A(n_628), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_628), .B(n_708), .Y(n_800) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g632 ( .A(n_629), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g761 ( .A(n_629), .B(n_676), .Y(n_761) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
OR2x2_ASAP7_75t_L g706 ( .A(n_632), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g663 ( .A(n_633), .Y(n_663) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g689 ( .A(n_636), .B(n_690), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_645), .B(n_646), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g652 ( .A(n_640), .B(n_649), .Y(n_652) );
BUFx2_ASAP7_75t_L g670 ( .A(n_640), .Y(n_670) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g681 ( .A(n_641), .Y(n_681) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g696 ( .A(n_643), .B(n_660), .Y(n_696) );
INVx2_ASAP7_75t_L g712 ( .A(n_643), .Y(n_712) );
AND2x2_ASAP7_75t_L g754 ( .A(n_643), .B(n_676), .Y(n_754) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g729 ( .A(n_649), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g776 ( .A(n_650), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g807 ( .A(n_651), .Y(n_807) );
INVx2_ASAP7_75t_L g746 ( .A(n_654), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_665), .C(n_682), .D(n_697), .Y(n_655) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_658), .A2(n_736), .B1(n_752), .B2(n_754), .C(n_755), .Y(n_751) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g733 ( .A(n_662), .Y(n_733) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx2_ASAP7_75t_L g726 ( .A(n_663), .Y(n_726) );
INVx2_ASAP7_75t_L g798 ( .A(n_664), .Y(n_798) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B1(n_671), .B2(n_674), .C1(n_677), .C2(n_681), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g752 ( .A(n_668), .B(n_753), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_668), .A2(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g791 ( .A(n_669), .B(n_735), .Y(n_791) );
OAI21xp33_ASAP7_75t_SL g765 ( .A1(n_670), .A2(n_691), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g684 ( .A(n_673), .B(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_673), .Y(n_736) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g735 ( .A(n_676), .Y(n_735) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g741 ( .A(n_680), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_686), .B1(n_691), .B2(n_696), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_688), .A2(n_698), .B1(n_701), .B2(n_703), .C(n_705), .Y(n_697) );
INVx3_ASAP7_75t_R g812 ( .A(n_689), .Y(n_812) );
INVx1_ASAP7_75t_L g730 ( .A(n_690), .Y(n_730) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_693), .Y(n_747) );
INVx1_ASAP7_75t_L g757 ( .A(n_693), .Y(n_757) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_702), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g775 ( .A(n_702), .Y(n_775) );
AND2x2_ASAP7_75t_L g803 ( .A(n_702), .B(n_750), .Y(n_803) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g797 ( .A(n_707), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_769), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_751), .C(n_765), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_727), .C(n_737), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI21xp33_ASAP7_75t_L g728 ( .A1(n_718), .A2(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g768 ( .A(n_720), .Y(n_768) );
AND2x2_ASAP7_75t_L g809 ( .A(n_720), .B(n_798), .Y(n_809) );
NAND2x1_ASAP7_75t_L g767 ( .A(n_721), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g789 ( .A(n_726), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_732), .Y(n_727) );
INVx1_ASAP7_75t_L g781 ( .A(n_735), .Y(n_781) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_742), .B1(n_744), .B2(n_748), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g777 ( .A(n_741), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_743), .B(n_773), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g816 ( .A(n_749), .Y(n_816) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp33_ASAP7_75t_SL g755 ( .A1(n_756), .A2(n_758), .B1(n_760), .B2(n_762), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_796), .Y(n_769) );
O2A1O1Ixp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_774), .B(n_776), .C(n_778), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OAI21xp33_ASAP7_75t_L g785 ( .A1(n_772), .A2(n_786), .B(n_788), .Y(n_785) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
O2A1O1Ixp5_ASAP7_75t_SL g796 ( .A1(n_776), .A2(n_797), .B(n_799), .C(n_801), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_780), .A2(n_785), .B1(n_790), .B2(n_792), .Y(n_784) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI211xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_804), .B(n_808), .C(n_815), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_812), .B2(n_813), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI21xp5_ASAP7_75t_SL g815 ( .A1(n_816), .A2(n_817), .B(n_819), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_R g835 ( .A(n_836), .B(n_837), .Y(n_835) );
CKINVDCx16_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
endmodule