module real_aes_5671_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_932;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g608 ( .A(n_0), .B(n_307), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_1), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_SL g655 ( .A1(n_2), .A2(n_200), .B(n_656), .C(n_657), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_3), .A2(n_79), .B1(n_149), .B2(n_198), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_4), .A2(n_30), .B1(n_134), .B2(n_138), .Y(n_133) );
INVxp67_ASAP7_75t_L g107 ( .A(n_5), .Y(n_107) );
INVx1_ASAP7_75t_L g547 ( .A(n_5), .Y(n_547) );
INVx1_ASAP7_75t_L g906 ( .A(n_5), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_6), .A2(n_86), .B1(n_214), .B2(n_215), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_7), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_8), .A2(n_66), .B1(n_136), .B2(n_198), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_9), .A2(n_31), .B1(n_174), .B2(n_175), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_10), .Y(n_586) );
INVx2_ASAP7_75t_L g321 ( .A(n_11), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_12), .A2(n_58), .B1(n_149), .B2(n_176), .Y(n_572) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_13), .A2(n_65), .B(n_159), .Y(n_158) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_13), .A2(n_65), .B(n_159), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_14), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_SL g319 ( .A(n_15), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_16), .B(n_259), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_17), .Y(n_632) );
BUFx3_ASAP7_75t_L g116 ( .A(n_18), .Y(n_116) );
BUFx8_ASAP7_75t_SL g944 ( .A(n_18), .Y(n_944) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_19), .A2(n_153), .B(n_273), .C(n_661), .Y(n_660) );
OAI22xp33_ASAP7_75t_SL g611 ( .A1(n_20), .A2(n_47), .B1(n_149), .B2(n_255), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_21), .A2(n_29), .B1(n_151), .B2(n_255), .Y(n_600) );
O2A1O1Ixp5_ASAP7_75t_L g263 ( .A1(n_22), .A2(n_142), .B(n_264), .C(n_267), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_23), .B(n_148), .Y(n_249) );
O2A1O1Ixp5_ASAP7_75t_L g556 ( .A1(n_24), .A2(n_200), .B(n_313), .C(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_26), .B(n_916), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_27), .Y(n_937) );
INVx1_ASAP7_75t_SL g272 ( .A(n_28), .Y(n_272) );
AND2x2_ASAP7_75t_L g118 ( .A(n_32), .B(n_119), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_33), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_34), .B(n_156), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_35), .A2(n_39), .B1(n_147), .B2(n_150), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_36), .A2(n_64), .B1(n_150), .B2(n_197), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_37), .B(n_139), .Y(n_248) );
INVx2_ASAP7_75t_L g190 ( .A(n_38), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_40), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_41), .B(n_184), .Y(n_220) );
OAI22xp33_ASAP7_75t_SL g931 ( .A1(n_42), .A2(n_90), .B1(n_932), .B2(n_933), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_42), .Y(n_932) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_43), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_44), .A2(n_153), .B(n_316), .C(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g295 ( .A(n_45), .Y(n_295) );
INVx2_ASAP7_75t_L g274 ( .A(n_46), .Y(n_274) );
INVx1_ASAP7_75t_L g159 ( .A(n_48), .Y(n_159) );
AND2x4_ASAP7_75t_L g162 ( .A(n_49), .B(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g205 ( .A(n_49), .B(n_163), .Y(n_205) );
INVx2_ASAP7_75t_L g199 ( .A(n_50), .Y(n_199) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_51), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_52), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_53), .Y(n_564) );
INVx2_ASAP7_75t_L g590 ( .A(n_54), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_55), .A2(n_200), .B(n_634), .C(n_635), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_56), .Y(n_619) );
INVx1_ASAP7_75t_SL g268 ( .A(n_57), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_59), .A2(n_75), .B1(n_135), .B2(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_60), .B(n_259), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_61), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_62), .Y(n_623) );
NAND2xp33_ASAP7_75t_R g575 ( .A(n_63), .B(n_166), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_63), .A2(n_99), .B1(n_156), .B2(n_820), .Y(n_819) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_67), .A2(n_134), .B(n_153), .C(n_202), .Y(n_201) );
OR2x6_ASAP7_75t_L g109 ( .A(n_68), .B(n_110), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g281 ( .A(n_69), .Y(n_281) );
INVx1_ASAP7_75t_L g291 ( .A(n_70), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_71), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_72), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_73), .B(n_174), .Y(n_256) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_74), .B(n_313), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_76), .A2(n_194), .B(n_196), .C(n_200), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_76), .A2(n_194), .B(n_196), .C(n_200), .Y(n_232) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_78), .A2(n_89), .B1(n_909), .B2(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_78), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_80), .A2(n_92), .B1(n_179), .B2(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_82), .Y(n_141) );
BUFx5_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
INVx2_ASAP7_75t_L g665 ( .A(n_83), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_84), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g638 ( .A(n_85), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_87), .Y(n_662) );
INVx2_ASAP7_75t_SL g163 ( .A(n_88), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_89), .Y(n_910) );
INVx1_ASAP7_75t_L g933 ( .A(n_90), .Y(n_933) );
INVx1_ASAP7_75t_L g562 ( .A(n_91), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_93), .B(n_166), .Y(n_292) );
INVx1_ASAP7_75t_SL g167 ( .A(n_94), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_95), .B(n_206), .Y(n_277) );
INVx2_ASAP7_75t_L g566 ( .A(n_96), .Y(n_566) );
AND2x2_ASAP7_75t_L g185 ( .A(n_97), .B(n_186), .Y(n_185) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_98), .A2(n_149), .B(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_99), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_99), .B(n_156), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_120), .B(n_920), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_113), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx12f_ASAP7_75t_L g927 ( .A(n_105), .Y(n_927) );
BUFx6f_ASAP7_75t_L g947 ( .A(n_105), .Y(n_947) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x6_ASAP7_75t_L g546 ( .A(n_108), .B(n_547), .Y(n_546) );
INVx8_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g905 ( .A(n_109), .B(n_906), .Y(n_905) );
OR2x6_ASAP7_75t_L g919 ( .A(n_109), .B(n_906), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
CKINVDCx6p67_ASAP7_75t_R g924 ( .A(n_116), .Y(n_924) );
OR2x2_ASAP7_75t_SL g922 ( .A(n_117), .B(n_923), .Y(n_922) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_118), .A2(n_943), .B(n_945), .Y(n_942) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_907), .B1(n_908), .B2(n_911), .C(n_915), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
OAI22x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_543), .B1(n_548), .B2(n_903), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g912 ( .A(n_125), .Y(n_912) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_433), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_359), .C(n_393), .D(n_402), .Y(n_126) );
O2A1O1Ixp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_221), .B(n_237), .C(n_297), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_168), .Y(n_128) );
INVxp67_ASAP7_75t_L g367 ( .A(n_129), .Y(n_367) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g223 ( .A(n_130), .B(n_224), .Y(n_223) );
NAND2x1_ASAP7_75t_L g382 ( .A(n_130), .B(n_236), .Y(n_382) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_130), .B(n_228), .Y(n_391) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g330 ( .A(n_131), .Y(n_330) );
AOI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_145), .B(n_164), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_142), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_134), .B(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g656 ( .A(n_135), .Y(n_656) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g151 ( .A(n_137), .Y(n_151) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
INVx1_ASAP7_75t_L g313 ( .A(n_140), .Y(n_313) );
INVx1_ASAP7_75t_L g560 ( .A(n_140), .Y(n_560) );
INVx1_ASAP7_75t_L g634 ( .A(n_140), .Y(n_634) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx2_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
INVx6_ASAP7_75t_L g255 ( .A(n_141), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_142), .B(n_178), .Y(n_177) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OA22x2_ASAP7_75t_L g599 ( .A1(n_143), .A2(n_600), .B1(n_601), .B2(n_603), .Y(n_599) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
INVxp67_ASAP7_75t_L g217 ( .A(n_144), .Y(n_217) );
INVx4_ASAP7_75t_L g251 ( .A(n_144), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_144), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g603 ( .A(n_144), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_144), .B(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_152), .B(n_154), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx2_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
INVx1_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
INVx2_ASAP7_75t_L g214 ( .A(n_149), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g310 ( .A(n_149), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_149), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_149), .B(n_564), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_149), .A2(n_255), .B1(n_586), .B2(n_587), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_149), .A2(n_255), .B1(n_619), .B2(n_620), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_149), .A2(n_176), .B1(n_622), .B2(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_149), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_151), .A2(n_176), .B1(n_589), .B2(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_151), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_151), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_152), .B(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_153), .A2(n_613), .B(n_614), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_153), .A2(n_162), .B1(n_200), .B2(n_618), .C(n_621), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_160), .Y(n_154) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_155), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g307 ( .A(n_157), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_157), .B(n_162), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g664 ( .A(n_157), .B(n_665), .Y(n_664) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx2_ASAP7_75t_L g245 ( .A(n_158), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_160), .A2(n_247), .B(n_252), .Y(n_246) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_161), .A2(n_243), .B(n_292), .Y(n_296) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g182 ( .A(n_162), .B(n_183), .Y(n_182) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
INVx1_ASAP7_75t_L g276 ( .A(n_162), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_167), .Y(n_164) );
INVx1_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
INVx1_ASAP7_75t_L g820 ( .A(n_165), .Y(n_820) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx3_ASAP7_75t_L g186 ( .A(n_166), .Y(n_186) );
INVx1_ASAP7_75t_L g191 ( .A(n_166), .Y(n_191) );
INVx1_ASAP7_75t_L g567 ( .A(n_166), .Y(n_567) );
INVx1_ASAP7_75t_L g628 ( .A(n_166), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_168), .A2(n_378), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_168), .Y(n_440) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_187), .Y(n_168) );
INVx1_ASAP7_75t_L g350 ( .A(n_169), .Y(n_350) );
AND2x6_ASAP7_75t_SL g365 ( .A(n_169), .B(n_223), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_169), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_169), .B(n_391), .Y(n_390) );
BUFx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_170), .B(n_208), .Y(n_325) );
AND2x2_ASAP7_75t_L g470 ( .A(n_170), .B(n_188), .Y(n_470) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_SL g236 ( .A(n_171), .Y(n_236) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_177), .A3(n_182), .B(n_185), .Y(n_171) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g273 ( .A(n_176), .Y(n_273) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_176), .Y(n_316) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g289 ( .A(n_181), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_183), .B(n_211), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_183), .A2(n_646), .B(n_647), .Y(n_645) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_184), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g583 ( .A(n_186), .Y(n_583) );
INVx1_ASAP7_75t_L g485 ( .A(n_187), .Y(n_485) );
NOR2x1_ASAP7_75t_L g187 ( .A(n_188), .B(n_207), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_188), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g370 ( .A(n_188), .Y(n_370) );
AND2x4_ASAP7_75t_L g396 ( .A(n_188), .B(n_235), .Y(n_396) );
INVx1_ASAP7_75t_L g406 ( .A(n_188), .Y(n_406) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_192), .Y(n_188) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_189), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx1_ASAP7_75t_L g209 ( .A(n_191), .Y(n_209) );
NOR4xp25_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .C(n_204), .D(n_206), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_197), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g271 ( .A(n_197), .Y(n_271) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g286 ( .A(n_198), .Y(n_286) );
INVx2_ASAP7_75t_SL g219 ( .A(n_200), .Y(n_219) );
INVx1_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_200), .B(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_200), .B(n_295), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_200), .A2(n_251), .B1(n_572), .B2(n_573), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_200), .A2(n_251), .B1(n_585), .B2(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g693 ( .A(n_200), .Y(n_693) );
INVxp67_ASAP7_75t_SL g233 ( .A(n_201), .Y(n_233) );
NOR2x1_ASAP7_75t_SL g304 ( .A(n_204), .B(n_305), .Y(n_304) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_204), .B(n_556), .C(n_559), .Y(n_555) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_204), .B(n_307), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_204), .A2(n_250), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_690) );
INVx4_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_205), .B(n_583), .Y(n_598) );
AND2x2_ASAP7_75t_L g627 ( .A(n_205), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g349 ( .A(n_208), .B(n_336), .Y(n_349) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_208), .Y(n_358) );
INVx1_ASAP7_75t_L g525 ( .A(n_208), .Y(n_525) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_220), .Y(n_208) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_209), .A2(n_246), .B(n_258), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_211), .B(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_212), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B1(n_218), .B2(n_219), .Y(n_212) );
OAI21xp5_ASAP7_75t_SL g269 ( .A1(n_216), .A2(n_270), .B(n_275), .Y(n_269) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g226 ( .A(n_220), .Y(n_226) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_227), .Y(n_222) );
AND2x2_ASAP7_75t_L g456 ( .A(n_223), .B(n_375), .Y(n_456) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_223), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_223), .B(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g335 ( .A(n_224), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g427 ( .A(n_224), .Y(n_427) );
AND2x2_ASAP7_75t_L g356 ( .A(n_227), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g379 ( .A(n_227), .B(n_367), .Y(n_379) );
AND2x4_ASAP7_75t_L g542 ( .A(n_227), .B(n_395), .Y(n_542) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_235), .Y(n_227) );
AND2x4_ASAP7_75t_L g376 ( .A(n_228), .B(n_336), .Y(n_376) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_228), .Y(n_522) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_234), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g334 ( .A(n_235), .Y(n_334) );
BUFx2_ASAP7_75t_SL g375 ( .A(n_235), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_235), .B(n_427), .Y(n_507) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_237), .A2(n_376), .B1(n_394), .B2(n_397), .C(n_400), .Y(n_393) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_239), .B(n_260), .Y(n_238) );
INVx2_ASAP7_75t_L g399 ( .A(n_239), .Y(n_399) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g412 ( .A(n_240), .B(n_345), .Y(n_412) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_240), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_240), .B(n_278), .Y(n_454) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g373 ( .A(n_241), .B(n_279), .Y(n_373) );
AND2x2_ASAP7_75t_L g416 ( .A(n_241), .B(n_261), .Y(n_416) );
AND2x2_ASAP7_75t_L g491 ( .A(n_241), .B(n_355), .Y(n_491) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .B(n_258), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_244), .A2(n_555), .B(n_565), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_244), .B(n_690), .Y(n_689) );
BUFx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g259 ( .A(n_245), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_245), .B(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_245), .B(n_638), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_250), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_250), .A2(n_630), .B(n_633), .Y(n_629) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
O2A1O1Ixp5_ASAP7_75t_SL g280 ( .A1(n_251), .A2(n_281), .B(n_282), .C(n_285), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_251), .A2(n_560), .B1(n_561), .B2(n_563), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .B(n_257), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g266 ( .A(n_255), .Y(n_266) );
INVx1_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
INVx2_ASAP7_75t_L g318 ( .A(n_255), .Y(n_318) );
INVx2_ASAP7_75t_SL g602 ( .A(n_255), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_257), .A2(n_309), .B(n_312), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_259), .B(n_276), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_260), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_278), .Y(n_260) );
INVx2_ASAP7_75t_SL g340 ( .A(n_261), .Y(n_340) );
BUFx2_ASAP7_75t_L g519 ( .A(n_261), .Y(n_519) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
INVx3_ASAP7_75t_L g348 ( .A(n_262), .Y(n_348) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_269), .B(n_277), .Y(n_262) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_273), .B2(n_274), .Y(n_270) );
AND2x4_ASAP7_75t_L g302 ( .A(n_278), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g477 ( .A(n_278), .B(n_303), .Y(n_477) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g363 ( .A(n_279), .B(n_347), .Y(n_363) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_287), .B(n_296), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_280), .A2(n_287), .B(n_296), .Y(n_342) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_283), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND3x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .C(n_293), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_322), .B(n_331), .C(n_343), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
AND2x2_ASAP7_75t_L g452 ( .A(n_300), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_300), .B(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g476 ( .A(n_300), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_R g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g421 ( .A(n_301), .Y(n_421) );
INVx2_ASAP7_75t_L g392 ( .A(n_302), .Y(n_392) );
AND2x2_ASAP7_75t_L g398 ( .A(n_302), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_302), .B(n_421), .Y(n_420) );
OAI322xp33_ASAP7_75t_L g448 ( .A1(n_302), .A2(n_378), .A3(n_449), .B1(n_451), .B2(n_455), .C1(n_457), .C2(n_463), .Y(n_448) );
AND2x2_ASAP7_75t_L g536 ( .A(n_302), .B(n_491), .Y(n_536) );
OR2x2_ASAP7_75t_L g341 ( .A(n_303), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx1_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
AND2x2_ASAP7_75t_L g527 ( .A(n_303), .B(n_342), .Y(n_527) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_303), .Y(n_539) );
AO31x2_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_308), .A3(n_314), .B(n_320), .Y(n_303) );
OA21x2_ASAP7_75t_L g616 ( .A1(n_305), .A2(n_617), .B(n_624), .Y(n_616) );
OA21x2_ASAP7_75t_L g717 ( .A1(n_305), .A2(n_617), .B(n_624), .Y(n_717) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g591 ( .A(n_306), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_318), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g426 ( .A(n_329), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g432 ( .A(n_329), .Y(n_432) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_329), .Y(n_531) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g336 ( .A(n_330), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_337), .Y(n_331) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_332), .B(n_365), .C(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g425 ( .A(n_334), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g495 ( .A(n_334), .Y(n_495) );
INVx2_ASAP7_75t_L g395 ( .A(n_335), .Y(n_395) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g541 ( .A(n_339), .B(n_373), .Y(n_541) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g372 ( .A(n_340), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g397 ( .A(n_340), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g447 ( .A(n_340), .B(n_341), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_340), .B(n_495), .C(n_522), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_341), .A2(n_436), .B(n_438), .Y(n_435) );
OAI31xp33_ASAP7_75t_L g439 ( .A1(n_341), .A2(n_440), .A3(n_441), .B(n_442), .Y(n_439) );
AOI32xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_349), .A3(n_350), .B1(n_351), .B2(n_356), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x2_ASAP7_75t_L g409 ( .A(n_345), .B(n_355), .Y(n_409) );
INVx1_ASAP7_75t_L g461 ( .A(n_345), .Y(n_461) );
INVx1_ASAP7_75t_L g473 ( .A(n_345), .Y(n_473) );
AND2x2_ASAP7_75t_L g486 ( .A(n_345), .B(n_373), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_345), .Y(n_490) );
OR2x2_ASAP7_75t_L g493 ( .A(n_345), .B(n_459), .Y(n_493) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
INVx1_ASAP7_75t_L g514 ( .A(n_346), .Y(n_514) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g354 ( .A(n_347), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_348), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_348), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g418 ( .A(n_349), .Y(n_418) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g362 ( .A(n_353), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g513 ( .A(n_353), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g378 ( .A(n_354), .Y(n_378) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_354), .Y(n_441) );
AND2x2_ASAP7_75t_L g411 ( .A(n_355), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g422 ( .A(n_356), .Y(n_422) );
INVx1_ASAP7_75t_L g469 ( .A(n_357), .Y(n_469) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
NOR2x1p5_ASAP7_75t_L g445 ( .A(n_358), .B(n_382), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_358), .B(n_376), .Y(n_497) );
NOR2xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_380), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_371), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_362), .B(n_374), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_363), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g472 ( .A(n_363), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_363), .B(n_421), .Y(n_492) );
INVx1_ASAP7_75t_L g442 ( .A(n_365), .Y(n_442) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_367), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_369), .B(n_459), .Y(n_462) );
INVx1_ASAP7_75t_L g444 ( .A(n_370), .Y(n_444) );
AND2x2_ASAP7_75t_L g450 ( .A(n_370), .B(n_432), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B1(n_377), .B2(n_379), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_372), .A2(n_411), .B(n_413), .Y(n_410) );
INVx2_ASAP7_75t_L g459 ( .A(n_373), .Y(n_459) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_384), .C(n_392), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g484 ( .A(n_382), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g482 ( .A(n_383), .Y(n_482) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_386), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_386), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g480 ( .A(n_390), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_391), .A2(n_482), .B1(n_483), .B2(n_486), .Y(n_481) );
AND2x2_ASAP7_75t_L g505 ( .A(n_391), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_396), .Y(n_413) );
INVx2_ASAP7_75t_SL g419 ( .A(n_396), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_396), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g530 ( .A(n_396), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI211xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B(n_414), .C(n_423), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_407), .B(n_410), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g430 ( .A(n_409), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_412), .A2(n_541), .B(n_542), .Y(n_540) );
OAI22xp33_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_417), .B1(n_420), .B2(n_422), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_416), .B(n_533), .Y(n_532) );
NAND2x1_ASAP7_75t_SL g538 ( .A(n_416), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g500 ( .A(n_426), .Y(n_500) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_430), .B(n_479), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_465), .C(n_508), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_439), .B1(n_443), .B2(n_446), .C(n_448), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_438), .A2(n_499), .B1(n_501), .B2(n_502), .C(n_503), .Y(n_498) );
INVx1_ASAP7_75t_L g510 ( .A(n_443), .Y(n_510) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_445), .Y(n_535) );
INVxp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_456), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .Y(n_457) );
INVx2_ASAP7_75t_SL g501 ( .A(n_458), .Y(n_501) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_487), .C(n_498), .Y(n_465) );
OAI211xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_471), .B(n_474), .C(n_481), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g533 ( .A(n_473), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_478), .B(n_480), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI31xp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_492), .A3(n_493), .B(n_494), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_488), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_495), .Y(n_517) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g511 ( .A(n_505), .Y(n_511) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI211xp5_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_512), .B(n_515), .C(n_528), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_518), .B(n_520), .C(n_526), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI211xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B(n_534), .C(n_540), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g914 ( .A(n_543), .Y(n_914) );
BUFx12f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
CKINVDCx11_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI22x1_ASAP7_75t_L g911 ( .A1(n_548), .A2(n_904), .B1(n_912), .B2(n_913), .Y(n_911) );
AND4x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_762), .C(n_802), .D(n_870), .Y(n_548) );
NAND4xp75_ASAP7_75t_L g934 ( .A(n_549), .B(n_762), .C(n_802), .D(n_870), .Y(n_934) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_700), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_551), .B(n_680), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_576), .B(n_593), .C(n_639), .Y(n_551) );
AND2x2_ASAP7_75t_L g694 ( .A(n_552), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_552), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g748 ( .A(n_552), .Y(n_748) );
AND2x2_ASAP7_75t_L g768 ( .A(n_552), .B(n_641), .Y(n_768) );
AND2x2_ASAP7_75t_L g869 ( .A(n_552), .B(n_850), .Y(n_869) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_568), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_553), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g895 ( .A(n_553), .B(n_834), .Y(n_895) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g667 ( .A(n_554), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g674 ( .A(n_554), .Y(n_674) );
BUFx2_ASAP7_75t_R g734 ( .A(n_554), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_554), .B(n_653), .Y(n_842) );
AND2x2_ASAP7_75t_L g846 ( .A(n_554), .B(n_652), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_SL g578 ( .A(n_568), .Y(n_578) );
INVx1_ASAP7_75t_L g675 ( .A(n_568), .Y(n_675) );
AND2x2_ASAP7_75t_L g757 ( .A(n_568), .B(n_652), .Y(n_757) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g668 ( .A(n_569), .Y(n_668) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_569), .Y(n_684) );
AND2x2_ASAP7_75t_L g772 ( .A(n_569), .B(n_674), .Y(n_772) );
AND2x2_ASAP7_75t_L g843 ( .A(n_569), .B(n_581), .Y(n_843) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
AND2x2_ASAP7_75t_L g818 ( .A(n_570), .B(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_579), .B(n_666), .Y(n_892) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g759 ( .A(n_581), .B(n_653), .Y(n_759) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B(n_591), .Y(n_581) );
INVx1_ASAP7_75t_L g691 ( .A(n_585), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_588), .Y(n_692) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_605), .Y(n_594) );
AND2x4_ASAP7_75t_L g677 ( .A(n_595), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g761 ( .A(n_596), .B(n_730), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_596), .B(n_755), .Y(n_774) );
OR2x2_ASAP7_75t_L g877 ( .A(n_596), .B(n_833), .Y(n_877) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g714 ( .A(n_597), .Y(n_714) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_604), .Y(n_597) );
INVx1_ASAP7_75t_L g646 ( .A(n_599), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_604), .Y(n_647) );
BUFx2_ASAP7_75t_SL g742 ( .A(n_605), .Y(n_742) );
NOR2xp67_ASAP7_75t_L g605 ( .A(n_606), .B(n_615), .Y(n_605) );
INVx1_ASAP7_75t_L g697 ( .A(n_606), .Y(n_697) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g679 ( .A(n_607), .Y(n_679) );
INVx3_ASAP7_75t_L g716 ( .A(n_607), .Y(n_716) );
AND2x2_ASAP7_75t_L g751 ( .A(n_607), .B(n_717), .Y(n_751) );
AND2x2_ASAP7_75t_L g781 ( .A(n_607), .B(n_625), .Y(n_781) );
AND2x4_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_625), .Y(n_615) );
INVx2_ASAP7_75t_L g648 ( .A(n_616), .Y(n_648) );
INVx2_ASAP7_75t_L g699 ( .A(n_616), .Y(n_699) );
INVx1_ASAP7_75t_L g642 ( .A(n_625), .Y(n_642) );
AND2x2_ASAP7_75t_L g698 ( .A(n_625), .B(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g724 ( .A(n_625), .B(n_679), .Y(n_724) );
INVx2_ASAP7_75t_L g730 ( .A(n_625), .Y(n_730) );
AND2x2_ASAP7_75t_L g755 ( .A(n_625), .B(n_716), .Y(n_755) );
BUFx2_ASAP7_75t_L g823 ( .A(n_625), .Y(n_823) );
INVx2_ASAP7_75t_L g834 ( .A(n_625), .Y(n_834) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI21x1_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_637), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_649), .B1(n_669), .B2(n_676), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g736 ( .A(n_644), .B(n_729), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_644), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_SL g829 ( .A(n_644), .Y(n_829) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
OR2x2_ASAP7_75t_L g722 ( .A(n_645), .B(n_717), .Y(n_722) );
AND2x4_ASAP7_75t_L g678 ( .A(n_648), .B(n_679), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_649), .B(n_703), .C(n_707), .Y(n_702) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_666), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g685 ( .A(n_651), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g695 ( .A(n_653), .B(n_687), .Y(n_695) );
INVx1_ASAP7_75t_L g706 ( .A(n_653), .Y(n_706) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_653), .Y(n_710) );
OR2x2_ASAP7_75t_L g739 ( .A(n_653), .B(n_687), .Y(n_739) );
INVx1_ASAP7_75t_L g776 ( .A(n_653), .Y(n_776) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_653), .Y(n_897) );
AO31x2_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_659), .A3(n_663), .B(n_664), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g725 ( .A(n_666), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g737 ( .A(n_667), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g746 ( .A(n_667), .B(n_695), .Y(n_746) );
AND2x4_ASAP7_75t_L g782 ( .A(n_667), .B(n_759), .Y(n_782) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g826 ( .A(n_672), .B(n_710), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_673), .B(n_687), .Y(n_866) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_674), .Y(n_801) );
AND2x2_ASAP7_75t_L g851 ( .A(n_674), .B(n_817), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_676), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g858 ( .A(n_677), .B(n_812), .Y(n_858) );
NAND2x1p5_ASAP7_75t_L g822 ( .A(n_678), .B(n_823), .Y(n_822) );
NAND2x1p5_ASAP7_75t_L g868 ( .A(n_678), .B(n_863), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_678), .B(n_761), .Y(n_881) );
AND2x2_ASAP7_75t_L g744 ( .A(n_679), .B(n_714), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_694), .B(n_696), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
AND2x2_ASAP7_75t_L g704 ( .A(n_683), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_683), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g785 ( .A(n_683), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_683), .B(n_837), .Y(n_836) );
INVx2_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g830 ( .A(n_685), .Y(n_830) );
INVx1_ASAP7_75t_L g901 ( .A(n_686), .Y(n_901) );
AND2x2_ASAP7_75t_L g705 ( .A(n_687), .B(n_706), .Y(n_705) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_687), .Y(n_791) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g817 ( .A(n_689), .B(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_695), .B(n_734), .Y(n_733) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_695), .Y(n_837) );
AOI22xp5_ASAP7_75t_SL g777 ( .A1(n_696), .A2(n_778), .B1(n_779), .B2(n_782), .Y(n_777) );
AND2x4_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_735), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_711), .B(n_718), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g749 ( .A(n_705), .Y(n_749) );
OR2x2_ASAP7_75t_L g815 ( .A(n_706), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g886 ( .A(n_706), .B(n_843), .Y(n_886) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_707), .Y(n_778) );
BUFx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g726 ( .A(n_709), .Y(n_726) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_712), .A2(n_781), .B(n_784), .C(n_787), .Y(n_783) );
OR2x2_ASAP7_75t_L g855 ( .A(n_712), .B(n_724), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_712), .B(n_715), .Y(n_889) );
AND2x2_ASAP7_75t_L g902 ( .A(n_712), .B(n_751), .Y(n_902) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g811 ( .A(n_713), .B(n_715), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_713), .B(n_751), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_713), .B(n_755), .Y(n_873) );
AND2x2_ASAP7_75t_L g878 ( .A(n_713), .B(n_781), .Y(n_878) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g767 ( .A(n_714), .Y(n_767) );
AND2x2_ASAP7_75t_L g884 ( .A(n_714), .B(n_717), .Y(n_884) );
AND2x2_ASAP7_75t_L g792 ( .A(n_715), .B(n_761), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_715), .B(n_823), .Y(n_854) );
AND2x4_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_716), .B(n_834), .Y(n_833) );
AND2x2_ASAP7_75t_L g766 ( .A(n_717), .B(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_719), .A2(n_725), .B1(n_727), .B2(n_731), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
AND2x2_ASAP7_75t_L g728 ( .A(n_721), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_721), .B(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g753 ( .A(n_722), .Y(n_753) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g812 ( .A(n_729), .Y(n_812) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g795 ( .A(n_730), .B(n_744), .Y(n_795) );
AND2x2_ASAP7_75t_L g797 ( .A(n_730), .B(n_751), .Y(n_797) );
INVx1_ASAP7_75t_L g864 ( .A(n_730), .Y(n_864) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_732), .A2(n_869), .B1(n_876), .B2(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g807 ( .A(n_734), .Y(n_807) );
AOI211xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_737), .B(n_740), .C(n_747), .Y(n_735) );
NOR2x1_ASAP7_75t_L g874 ( .A(n_737), .B(n_840), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_738), .B(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_743), .B(n_745), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI332xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .A3(n_750), .B1(n_752), .B2(n_754), .B3(n_756), .C1(n_758), .C2(n_760), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_751), .A2(n_840), .B1(n_844), .B2(n_845), .Y(n_839) );
INVxp67_ASAP7_75t_SL g844 ( .A(n_752), .Y(n_844) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g899 ( .A(n_754), .Y(n_899) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g865 ( .A(n_757), .B(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g900 ( .A(n_757), .B(n_901), .Y(n_900) );
INVx2_ASAP7_75t_SL g786 ( .A(n_759), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_759), .B(n_772), .Y(n_787) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND4x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_777), .C(n_783), .D(n_788), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_768), .B(n_769), .C(n_775), .Y(n_763) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
OAI321xp33_ASAP7_75t_L g890 ( .A1(n_765), .A2(n_831), .A3(n_844), .B1(n_891), .B2(n_893), .C(n_898), .Y(n_890) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_SL g850 ( .A(n_776), .Y(n_850) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_786), .A2(n_794), .B(n_796), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_792), .B(n_793), .C(n_798), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_797), .A2(n_814), .B1(n_821), .B2(n_824), .Y(n_813) );
INVxp67_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_838), .Y(n_802) );
OAI211xp5_ASAP7_75t_SL g803 ( .A1(n_804), .A2(n_808), .B(n_813), .C(n_827), .Y(n_803) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
OR2x2_ASAP7_75t_L g882 ( .A(n_812), .B(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_815), .B(n_889), .Y(n_888) );
OR2x2_ASAP7_75t_L g896 ( .A(n_816), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g857 ( .A(n_817), .Y(n_857) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AOI32xp33_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_830), .A3(n_831), .B1(n_832), .B2(n_835), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND3xp33_ASAP7_75t_SL g838 ( .A(n_839), .B(n_847), .C(n_859), .Y(n_838) );
AND2x4_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g845 ( .A(n_843), .B(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_843), .A2(n_899), .B1(n_900), .B2(n_902), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_852), .B1(n_856), .B2(n_858), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND2x1p5_ASAP7_75t_SL g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .C(n_855), .Y(n_852) );
A2O1A1Ixp33_ASAP7_75t_L g871 ( .A1(n_855), .A2(n_872), .B(n_874), .C(n_875), .Y(n_871) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_865), .B1(n_867), .B2(n_869), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_879), .C(n_890), .Y(n_870) );
BUFx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
A2O1A1Ixp33_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_882), .B(n_885), .C(n_887), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVxp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
NOR2x1_ASAP7_75t_L g894 ( .A(n_895), .B(n_896), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_904), .Y(n_903) );
BUFx8_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
BUFx3_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_925), .B1(n_932), .B2(n_939), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI21x1_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_928), .B(n_936), .Y(n_925) );
BUFx5_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
BUFx2_ASAP7_75t_L g938 ( .A(n_927), .Y(n_938) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OA22x2_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_931), .B1(n_934), .B2(n_935), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx2_ASAP7_75t_L g935 ( .A(n_934), .Y(n_935) );
NOR2xp33_ASAP7_75t_SL g936 ( .A(n_937), .B(n_938), .Y(n_936) );
CKINVDCx11_ASAP7_75t_R g939 ( .A(n_940), .Y(n_939) );
BUFx6f_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
CKINVDCx8_ASAP7_75t_R g941 ( .A(n_942), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx5_ASAP7_75t_SL g946 ( .A(n_947), .Y(n_946) );
endmodule