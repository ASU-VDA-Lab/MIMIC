module fake_netlist_6_2621_n_83 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_83);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_83;

wire n_52;
wire n_46;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_78;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_5),
.Y(n_25)
);

AND2x4_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx6p67_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_3),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_16),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_18),
.Y(n_50)
);

AO21x2_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_38),
.B(n_36),
.Y(n_51)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_25),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_23),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_25),
.B(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_43),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_58),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_28),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_50),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_47),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_45),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_65),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_68),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_62),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_62),
.B(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NAND4xp25_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_24),
.C(n_31),
.D(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_80),
.B(n_37),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_34),
.B1(n_37),
.B2(n_44),
.Y(n_82)
);

OR2x6_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);


endmodule