module fake_ariane_823_n_800 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_800);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_800;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_0),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_37),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_68),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_57),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_17),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_30),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_44),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_65),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_29),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_157),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_78),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_93),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_49),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_45),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_11),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_32),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_56),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_29),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_121),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_39),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_114),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_77),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_59),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_0),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_1),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_213),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_1),
.Y(n_231)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_179),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_181),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_213),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_194),
.B(n_2),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_175),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_162),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_165),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_204),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_2),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_3),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_209),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

AND3x2_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_214),
.C(n_212),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_224),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_235),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_188),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_222),
.A2(n_214),
.B(n_177),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_237),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_245),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_223),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_223),
.B(n_176),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_255),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_256),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_236),
.B(n_178),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_258),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_218),
.B(n_188),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_202),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_248),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_172),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_237),
.B(n_164),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_257),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_242),
.B(n_164),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_242),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_243),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_238),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_307),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_220),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_243),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_220),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_244),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_244),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_278),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_282),
.Y(n_327)
);

BUFx4f_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_263),
.B(n_221),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_231),
.B1(n_253),
.B2(n_254),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_261),
.B1(n_259),
.B2(n_246),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_246),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_274),
.B(n_259),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_267),
.B(n_261),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_207),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_227),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_286),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_279),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_207),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_294),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_285),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_168),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_3),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_169),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_171),
.Y(n_348)
);

OR2x6_ASAP7_75t_L g349 ( 
.A(n_265),
.B(n_4),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_302),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_173),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_270),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_288),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_292),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_283),
.B(n_180),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_283),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_273),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_276),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_281),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_269),
.B(n_4),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_305),
.B(n_286),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_290),
.B(n_182),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_264),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_290),
.A2(n_208),
.B1(n_206),
.B2(n_205),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_305),
.B(n_184),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_281),
.B(n_5),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_298),
.B(n_185),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_281),
.A2(n_203),
.B1(n_200),
.B2(n_199),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_264),
.Y(n_376)
);

NOR3xp33_ASAP7_75t_SL g377 ( 
.A(n_325),
.B(n_276),
.C(n_296),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_264),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_264),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_266),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_314),
.B(n_334),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_317),
.B(n_270),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_317),
.B(n_291),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_266),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_313),
.B(n_266),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_374),
.B(n_291),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_313),
.B(n_266),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_374),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_319),
.B(n_332),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_266),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_275),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_322),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_275),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_275),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_275),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_338),
.B(n_275),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_308),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_373),
.A2(n_308),
.B1(n_296),
.B2(n_192),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_340),
.B(n_308),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g410 ( 
.A(n_338),
.B(n_308),
.C(n_191),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_348),
.B(n_308),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_348),
.B(n_5),
.Y(n_413)
);

AO221x1_ASAP7_75t_L g414 ( 
.A1(n_350),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_340),
.B(n_189),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_346),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

OR2x6_ASAP7_75t_SL g418 ( 
.A(n_325),
.B(n_361),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_347),
.B(n_7),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_335),
.B(n_190),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_331),
.B(n_8),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_312),
.B(n_9),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_361),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_337),
.B(n_11),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_373),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_336),
.Y(n_426)
);

NAND2x1_ASAP7_75t_L g427 ( 
.A(n_323),
.B(n_34),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_341),
.B(n_12),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_369),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_364),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

BUFx8_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_352),
.B(n_15),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_328),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_16),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_369),
.B(n_18),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_326),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_346),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_19),
.Y(n_439)
);

NAND2x1_ASAP7_75t_L g440 ( 
.A(n_323),
.B(n_35),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_343),
.B(n_371),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_346),
.B(n_36),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_324),
.B(n_20),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_324),
.B(n_21),
.Y(n_444)
);

OAI22xp33_ASAP7_75t_L g445 ( 
.A1(n_349),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_423),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_381),
.B(n_357),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_430),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_379),
.A2(n_378),
.B(n_386),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_441),
.A2(n_354),
.B1(n_356),
.B2(n_349),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_442),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_330),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_393),
.B(n_342),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_442),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_413),
.A2(n_328),
.B(n_375),
.C(n_354),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_398),
.B(n_342),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_416),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_SL g465 ( 
.A(n_445),
.B(n_364),
.C(n_367),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_416),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_389),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_342),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_344),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_401),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_358),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_417),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_426),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_431),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_391),
.B(n_356),
.Y(n_481)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_425),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_413),
.B(n_356),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_408),
.A2(n_318),
.B1(n_349),
.B2(n_328),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_365),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_405),
.B(n_365),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_420),
.B(n_379),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_406),
.B(n_359),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_380),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_436),
.B(n_349),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_SL g495 ( 
.A(n_429),
.B(n_318),
.C(n_353),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_388),
.B(n_366),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_418),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_377),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_408),
.B(n_355),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_450),
.B(n_489),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_447),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_454),
.A2(n_419),
.B(n_433),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_459),
.A2(n_419),
.B(n_433),
.Y(n_503)
);

NOR2x1_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_383),
.Y(n_504)
);

O2A1O1Ixp5_ASAP7_75t_L g505 ( 
.A1(n_485),
.A2(n_435),
.B(n_412),
.C(n_409),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_475),
.B(n_439),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_404),
.B(n_399),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_499),
.A2(n_422),
.B(n_424),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_485),
.A2(n_407),
.B(n_428),
.Y(n_509)
);

AO31x2_ASAP7_75t_L g510 ( 
.A1(n_493),
.A2(n_412),
.A3(n_396),
.B(n_406),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_382),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_489),
.A2(n_385),
.B(n_403),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_460),
.B(n_366),
.Y(n_514)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_482),
.A2(n_439),
.B(n_421),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_467),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_490),
.A2(n_457),
.B(n_452),
.Y(n_517)
);

NOR2x1_ASAP7_75t_SL g518 ( 
.A(n_482),
.B(n_484),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_434),
.C(n_438),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_446),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_482),
.A2(n_444),
.B1(n_443),
.B2(n_415),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_468),
.A2(n_396),
.B(n_385),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_470),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_469),
.B(n_366),
.Y(n_525)
);

AO22x2_ASAP7_75t_L g526 ( 
.A1(n_495),
.A2(n_414),
.B1(n_410),
.B2(n_355),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_403),
.Y(n_527)
);

AOI21xp33_ASAP7_75t_L g528 ( 
.A1(n_482),
.A2(n_376),
.B(n_370),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_484),
.B(n_323),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_463),
.A2(n_376),
.B(n_370),
.Y(n_531)
);

NAND3x1_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_22),
.C(n_23),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_456),
.B(n_323),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_490),
.A2(n_376),
.B(n_370),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_484),
.B(n_481),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_452),
.A2(n_376),
.B(n_370),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_484),
.A2(n_376),
.B1(n_370),
.B2(n_323),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_484),
.B(n_24),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_473),
.B(n_25),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_473),
.B(n_26),
.Y(n_540)
);

AO31x2_ASAP7_75t_L g541 ( 
.A1(n_493),
.A2(n_94),
.A3(n_158),
.B(n_153),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_490),
.A2(n_90),
.B(n_151),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g543 ( 
.A(n_452),
.B(n_38),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_518),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_530),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_500),
.A2(n_457),
.B(n_462),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_L g548 ( 
.A(n_502),
.B(n_465),
.C(n_488),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_502),
.B(n_473),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_519),
.A2(n_494),
.B1(n_496),
.B2(n_492),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_503),
.A2(n_457),
.B(n_462),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_513),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_509),
.A2(n_534),
.B(n_517),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_512),
.A2(n_462),
.B(n_483),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_503),
.A2(n_471),
.B(n_455),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

AOI221xp5_ASAP7_75t_L g557 ( 
.A1(n_506),
.A2(n_494),
.B1(n_486),
.B2(n_496),
.C(n_470),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_519),
.A2(n_466),
.B1(n_494),
.B2(n_478),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_501),
.A2(n_466),
.B1(n_478),
.B2(n_458),
.Y(n_559)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_542),
.A2(n_483),
.B(n_476),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_453),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_527),
.A2(n_453),
.B1(n_458),
.B2(n_464),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_525),
.A2(n_453),
.B1(n_458),
.B2(n_448),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_529),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_510),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_505),
.A2(n_455),
.B(n_474),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_515),
.A2(n_496),
.B1(n_472),
.B2(n_479),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_522),
.A2(n_538),
.B(n_523),
.C(n_540),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_524),
.B(n_448),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_522),
.A2(n_458),
.B(n_453),
.C(n_472),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_526),
.A2(n_497),
.B1(n_449),
.B2(n_458),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_524),
.A2(n_477),
.B1(n_474),
.B2(n_479),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_523),
.A2(n_477),
.B(n_476),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_516),
.B(n_480),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_514),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_521),
.B(n_480),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_508),
.A2(n_480),
.B(n_487),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_533),
.A2(n_498),
.B(n_449),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_531),
.A2(n_487),
.B(n_95),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_498),
.B(n_27),
.C(n_28),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_536),
.A2(n_537),
.B(n_543),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_543),
.A2(n_487),
.B(n_92),
.Y(n_584)
);

AOI21xp33_ASAP7_75t_SL g585 ( 
.A1(n_526),
.A2(n_26),
.B(n_27),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_552),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_561),
.Y(n_588)
);

O2A1O1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_585),
.A2(n_504),
.B(n_511),
.C(n_514),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_577),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_552),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_570),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_548),
.A2(n_514),
.B1(n_528),
.B2(n_520),
.Y(n_595)
);

AOI221xp5_ASAP7_75t_L g596 ( 
.A1(n_585),
.A2(n_520),
.B1(n_532),
.B2(n_487),
.C(n_510),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_566),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_545),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_548),
.B(n_28),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_578),
.Y(n_600)
);

BUFx4_ASAP7_75t_R g601 ( 
.A(n_545),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_575),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_576),
.Y(n_603)
);

OAI221xp5_ASAP7_75t_L g604 ( 
.A1(n_582),
.A2(n_487),
.B1(n_541),
.B2(n_510),
.C(n_33),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_549),
.A2(n_541),
.B1(n_31),
.B2(n_32),
.Y(n_605)
);

A2O1A1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_569),
.A2(n_541),
.B(n_31),
.C(n_33),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_545),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_549),
.B(n_30),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_572),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_558),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_580),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_574),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_557),
.B(n_159),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_574),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_581),
.A2(n_51),
.B(n_52),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_566),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_550),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_572),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_559),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_564),
.A2(n_147),
.B1(n_70),
.B2(n_71),
.C(n_73),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_551),
.A2(n_144),
.B(n_75),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_578),
.B(n_143),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_555),
.B(n_69),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_578),
.B(n_76),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_578),
.B(n_79),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_568),
.B(n_80),
.C(n_81),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_561),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_561),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_571),
.A2(n_142),
.B(n_83),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_563),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_555),
.B(n_87),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_573),
.A2(n_141),
.B1(n_97),
.B2(n_98),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_562),
.A2(n_89),
.B1(n_99),
.B2(n_100),
.Y(n_637)
);

NAND4xp25_ASAP7_75t_SL g638 ( 
.A(n_595),
.B(n_544),
.C(n_547),
.D(n_556),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_611),
.B(n_565),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_599),
.A2(n_562),
.B1(n_544),
.B2(n_579),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_586),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_598),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_592),
.Y(n_643)
);

AOI222xp33_ASAP7_75t_L g644 ( 
.A1(n_599),
.A2(n_544),
.B1(n_556),
.B2(n_584),
.C1(n_567),
.C2(n_565),
.Y(n_644)
);

AOI222xp33_ASAP7_75t_L g645 ( 
.A1(n_605),
.A2(n_556),
.B1(n_584),
.B2(n_567),
.C1(n_565),
.C2(n_560),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_594),
.B(n_565),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_620),
.A2(n_562),
.B1(n_579),
.B2(n_560),
.Y(n_647)
);

OAI211xp5_ASAP7_75t_L g648 ( 
.A1(n_606),
.A2(n_596),
.B(n_595),
.C(n_608),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_602),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_603),
.B(n_562),
.Y(n_650)
);

AOI222xp33_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_581),
.B1(n_547),
.B2(n_554),
.C1(n_583),
.C2(n_546),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_590),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_620),
.A2(n_562),
.B1(n_579),
.B2(n_554),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_604),
.A2(n_546),
.B1(n_547),
.B2(n_583),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_622),
.A2(n_553),
.B1(n_102),
.B2(n_106),
.Y(n_655)
);

OAI221xp5_ASAP7_75t_L g656 ( 
.A1(n_606),
.A2(n_553),
.B1(n_108),
.B2(n_110),
.C(n_111),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_SL g657 ( 
.A1(n_609),
.A2(n_601),
.B1(n_630),
.B2(n_613),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_622),
.A2(n_101),
.B1(n_112),
.B2(n_113),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_601),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_619),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_600),
.B(n_124),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_600),
.B(n_125),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_589),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_619),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_664)
);

AOI222xp33_ASAP7_75t_L g665 ( 
.A1(n_636),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.C1(n_140),
.C2(n_623),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_616),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_632),
.B(n_628),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_610),
.A2(n_636),
.B1(n_627),
.B2(n_598),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_627),
.A2(n_598),
.B1(n_607),
.B2(n_590),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_634),
.A2(n_637),
.B1(n_633),
.B2(n_625),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_598),
.B(n_607),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_607),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_591),
.Y(n_673)
);

NAND4xp25_ASAP7_75t_L g674 ( 
.A(n_612),
.B(n_614),
.C(n_632),
.D(n_629),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_626),
.A2(n_635),
.B1(n_617),
.B2(n_621),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_624),
.A2(n_631),
.B(n_588),
.Y(n_676)
);

AOI221xp5_ASAP7_75t_L g677 ( 
.A1(n_621),
.A2(n_591),
.B1(n_607),
.B2(n_597),
.C(n_618),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_666),
.B(n_597),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_656),
.A2(n_615),
.B1(n_618),
.B2(n_588),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_666),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_639),
.B(n_631),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_643),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_674),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_652),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_673),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_675),
.B(n_615),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_675),
.B(n_631),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_646),
.B(n_631),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_651),
.B(n_587),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_650),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_642),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_657),
.A2(n_629),
.B1(n_665),
.B2(n_640),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_671),
.B(n_642),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_677),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_654),
.B(n_644),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_649),
.B(n_667),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_653),
.B(n_647),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_642),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_638),
.B(n_672),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_645),
.B(n_655),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_657),
.A2(n_659),
.B1(n_668),
.B2(n_670),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_676),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_648),
.B(n_669),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_662),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_659),
.B(n_662),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_661),
.Y(n_707)
);

OAI221xp5_ASAP7_75t_L g708 ( 
.A1(n_702),
.A2(n_658),
.B1(n_663),
.B2(n_660),
.C(n_664),
.Y(n_708)
);

OAI31xp33_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_701),
.A3(n_696),
.B(n_704),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_706),
.A2(n_701),
.B1(n_693),
.B2(n_696),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_680),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_701),
.A2(n_696),
.B1(n_698),
.B2(n_704),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_SL g713 ( 
.A1(n_698),
.A2(n_695),
.B1(n_700),
.B2(n_684),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_681),
.B(n_688),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_694),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_681),
.B(n_688),
.Y(n_716)
);

NOR4xp25_ASAP7_75t_SL g717 ( 
.A(n_703),
.B(n_680),
.C(n_695),
.D(n_682),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_705),
.Y(n_718)
);

AOI31xp33_ASAP7_75t_L g719 ( 
.A1(n_706),
.A2(n_684),
.A3(n_700),
.B(n_690),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_705),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_703),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_688),
.B(n_697),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_690),
.A2(n_707),
.B1(n_679),
.B2(n_687),
.Y(n_723)
);

CKINVDCx8_ASAP7_75t_R g724 ( 
.A(n_694),
.Y(n_724)
);

AOI222xp33_ASAP7_75t_SL g725 ( 
.A1(n_682),
.A2(n_707),
.B1(n_683),
.B2(n_685),
.C1(n_686),
.C2(n_699),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_685),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_711),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_722),
.B(n_697),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_722),
.B(n_678),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_726),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_714),
.B(n_690),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_714),
.B(n_716),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_718),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_721),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_719),
.B(n_689),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_726),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_716),
.B(n_689),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_718),
.B(n_691),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_721),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_733),
.B(n_732),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_733),
.B(n_720),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_731),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_736),
.B(n_719),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_732),
.B(n_720),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_729),
.B(n_718),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_741),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_R g748 ( 
.A(n_744),
.B(n_717),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_741),
.B(n_736),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_745),
.B(n_742),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_743),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_751),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_710),
.B1(n_708),
.B2(n_713),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_749),
.B(n_746),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_751),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_747),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_754),
.B(n_750),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_756),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_757),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_756),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_758),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_759),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_760),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_755),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_758),
.B(n_753),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_709),
.C(n_710),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_742),
.Y(n_767)
);

OAI221xp5_ASAP7_75t_SL g768 ( 
.A1(n_765),
.A2(n_709),
.B1(n_712),
.B2(n_708),
.C(n_723),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_761),
.B(n_725),
.C(n_717),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_764),
.A2(n_763),
.B1(n_745),
.B2(n_734),
.Y(n_770)
);

AOI221x1_ASAP7_75t_L g771 ( 
.A1(n_762),
.A2(n_713),
.B1(n_740),
.B2(n_735),
.C(n_728),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_770),
.B(n_729),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_767),
.Y(n_773)
);

NOR2x1_ASAP7_75t_L g774 ( 
.A(n_769),
.B(n_735),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_766),
.B(n_735),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_768),
.A2(n_721),
.B(n_727),
.C(n_728),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_773),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_772),
.B(n_771),
.Y(n_778)
);

AND4x1_ASAP7_75t_L g779 ( 
.A(n_776),
.B(n_739),
.C(n_738),
.D(n_725),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_775),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_774),
.B(n_738),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_778),
.A2(n_727),
.B(n_737),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_777),
.B(n_737),
.Y(n_783)
);

OAI211xp5_ASAP7_75t_L g784 ( 
.A1(n_780),
.A2(n_721),
.B(n_731),
.C(n_720),
.Y(n_784)
);

O2A1O1Ixp5_ASAP7_75t_L g785 ( 
.A1(n_781),
.A2(n_739),
.B(n_730),
.C(n_699),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_779),
.B(n_705),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_783),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_782),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_786),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_785),
.B(n_699),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_784),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_786),
.A2(n_692),
.B1(n_699),
.B2(n_687),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_788),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_793),
.A2(n_789),
.B1(n_792),
.B2(n_787),
.Y(n_794)
);

AO21x2_ASAP7_75t_L g795 ( 
.A1(n_794),
.A2(n_791),
.B(n_790),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_SL g796 ( 
.A1(n_795),
.A2(n_724),
.B1(n_692),
.B2(n_715),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_796),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_797),
.A2(n_692),
.B1(n_715),
.B2(n_687),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_686),
.B1(n_683),
.B2(n_694),
.C(n_678),
.Y(n_799)
);

AOI211xp5_ASAP7_75t_L g800 ( 
.A1(n_799),
.A2(n_694),
.B(n_678),
.C(n_691),
.Y(n_800)
);


endmodule