module real_jpeg_13356_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_4),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_37),
.C(n_40),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_28),
.C(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_4),
.A2(n_21),
.B1(n_66),
.B2(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_18),
.C(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_100),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_81),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_80),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_58),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_13),
.B(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_45),
.C(n_50),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_14)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_16),
.A2(n_33),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_16),
.A2(n_33),
.B1(n_47),
.B2(n_48),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_16),
.A2(n_33),
.B1(n_97),
.B2(n_101),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_16),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_22),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_23),
.Y(n_24)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_18),
.A2(n_19),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_21),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_21),
.B(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_33),
.C(n_43),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_27),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_27),
.B(n_76),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_27)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_28),
.A2(n_32),
.B1(n_66),
.B2(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_33),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_33),
.B(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_33),
.B(n_50),
.C(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_34),
.A2(n_43),
.B1(n_50),
.B2(n_79),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_34),
.A2(n_79),
.B(n_84),
.C(n_86),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_79),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B(n_42),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OA22x2_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_40),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_79),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_50),
.A2(n_79),
.B1(n_94),
.B2(n_112),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_57),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_69),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_90),
.B(n_118),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_114),
.B(n_117),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_102),
.B(n_113),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_110),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);


endmodule