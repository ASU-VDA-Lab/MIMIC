module fake_netlist_6_1064_n_1114 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1114);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1114;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_955;
wire n_284;
wire n_400;
wire n_337;
wire n_739;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_844;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_1060;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_212),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_30),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_30),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_209),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_58),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_56),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_27),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_64),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_48),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_101),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_99),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_24),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_6),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_49),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_45),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_46),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_123),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_67),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_187),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_23),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_98),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_21),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_100),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_118),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_53),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_63),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_62),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_165),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_61),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_130),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_96),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_42),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_91),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_25),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_29),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_10),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_12),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_71),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_129),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_188),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_132),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_102),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_110),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_147),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_18),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_82),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_177),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_84),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_88),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_145),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_190),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_81),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_215),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_213),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_263),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_255),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_214),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_227),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_231),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_218),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_220),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_218),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_217),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_262),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_215),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_224),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_264),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_221),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_246),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_240),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_240),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_225),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_222),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_295),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_236),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_266),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_298),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_329),
.A2(n_276),
.B1(n_267),
.B2(n_279),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_329),
.A2(n_240),
.B1(n_241),
.B2(n_248),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_238),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g353 ( 
.A1(n_332),
.A2(n_248),
.B(n_244),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_244),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_331),
.A2(n_260),
.B1(n_269),
.B2(n_282),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_325),
.B(n_241),
.Y(n_358)
);

OAI22x1_ASAP7_75t_R g359 ( 
.A1(n_294),
.A2(n_284),
.B1(n_283),
.B2(n_278),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_241),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_250),
.B1(n_274),
.B2(n_272),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_306),
.A2(n_269),
.B(n_260),
.Y(n_371)
);

OAI21x1_ASAP7_75t_L g372 ( 
.A1(n_321),
.A2(n_226),
.B(n_223),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_312),
.B(n_228),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_292),
.B(n_275),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_302),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_302),
.B(n_229),
.Y(n_383)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_303),
.B(n_232),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_303),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_233),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_339),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_336),
.A2(n_252),
.B1(n_268),
.B2(n_265),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_378),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_343),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_378),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_343),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_377),
.B(n_323),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_378),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_343),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_377),
.B(n_323),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_378),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_359),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_377),
.B(n_294),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_389),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_389),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_389),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_354),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_354),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_385),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_362),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_362),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_336),
.B(n_373),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_383),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_R g424 ( 
.A(n_382),
.B(n_234),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_387),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_358),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_336),
.B(n_237),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_381),
.B(n_239),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_380),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_386),
.B(n_259),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_379),
.B(n_242),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_258),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_367),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_341),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_R g438 ( 
.A(n_379),
.B(n_245),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_R g439 ( 
.A(n_388),
.B(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_341),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_349),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_357),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_379),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_388),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_351),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_336),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_353),
.A2(n_32),
.B(n_31),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_337),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_363),
.B(n_33),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_355),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_R g455 ( 
.A(n_365),
.B(n_211),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_337),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_384),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_346),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_363),
.B(n_34),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_358),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_337),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_365),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_335),
.B(n_36),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_335),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_347),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_413),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_442),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_409),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_347),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_423),
.A2(n_372),
.B1(n_347),
.B2(n_352),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_425),
.B(n_372),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_335),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_352),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_440),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_340),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_452),
.B(n_363),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_370),
.B1(n_369),
.B2(n_368),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_352),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_458),
.B(n_368),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_446),
.B(n_370),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_448),
.B(n_370),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_396),
.B(n_369),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_434),
.B(n_340),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_459),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_340),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_356),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_403),
.B(n_344),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_403),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_400),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_408),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_399),
.B(n_402),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_408),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_429),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_344),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_449),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_449),
.B(n_344),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_457),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_455),
.B(n_348),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_453),
.B(n_360),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_360),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_451),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_455),
.B(n_356),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_390),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_391),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_438),
.B(n_346),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_431),
.B(n_356),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_346),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_346),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_461),
.B(n_346),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_411),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_414),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_444),
.A2(n_371),
.B1(n_1),
.B2(n_2),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_428),
.B(n_371),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_416),
.B(n_418),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_398),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_401),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_424),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_417),
.B(n_0),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_490),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_498),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_501),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_534),
.B(n_432),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_475),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_477),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_465),
.B(n_404),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_484),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_501),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_470),
.B(n_371),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_479),
.A2(n_439),
.B1(n_407),
.B2(n_353),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_472),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_468),
.B(n_37),
.Y(n_565)
);

BUFx6f_ASAP7_75t_SL g566 ( 
.A(n_545),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_490),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_491),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_492),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_38),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_517),
.Y(n_574)
);

AO22x2_ASAP7_75t_L g575 ( 
.A1(n_529),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_531),
.B(n_3),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_547),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_533),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_533),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_476),
.B(n_527),
.Y(n_581)
);

AO22x2_ASAP7_75t_L g582 ( 
.A1(n_474),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_467),
.B(n_39),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_467),
.B(n_40),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_473),
.B(n_7),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_489),
.B(n_41),
.Y(n_589)
);

NAND2x1p5_ASAP7_75t_L g590 ( 
.A(n_490),
.B(n_476),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_510),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_504),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_541),
.A2(n_522),
.B1(n_543),
.B2(n_495),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_493),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_514),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_485),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_516),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_512),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_512),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_543),
.B(n_43),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_523),
.B(n_8),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_482),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

OAI221xp5_ASAP7_75t_L g606 ( 
.A1(n_536),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_521),
.B(n_44),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_538),
.B(n_47),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_548),
.B(n_9),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_544),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_11),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_546),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_505),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_520),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_553),
.B(n_598),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_550),
.Y(n_619)
);

AOI21x1_ASAP7_75t_L g620 ( 
.A1(n_594),
.A2(n_535),
.B(n_530),
.Y(n_620)
);

AO21x1_ASAP7_75t_L g621 ( 
.A1(n_587),
.A2(n_478),
.B(n_565),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_581),
.A2(n_519),
.B(n_497),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_556),
.A2(n_548),
.B1(n_468),
.B2(n_486),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_560),
.A2(n_480),
.B(n_519),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_559),
.B(n_468),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_599),
.A2(n_497),
.B(n_481),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_616),
.A2(n_502),
.B(n_481),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_597),
.A2(n_502),
.B(n_526),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_572),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_552),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_562),
.B(n_563),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_607),
.A2(n_526),
.B(n_525),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_589),
.A2(n_468),
.B1(n_494),
.B2(n_539),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_600),
.A2(n_525),
.B(n_524),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_601),
.A2(n_524),
.B(n_496),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_605),
.A2(n_488),
.B(n_482),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_568),
.B(n_554),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_615),
.B(n_542),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_566),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_551),
.A2(n_499),
.B(n_518),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_612),
.B(n_545),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_613),
.A2(n_537),
.B(n_532),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_564),
.B(n_466),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_583),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_551),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_561),
.A2(n_603),
.B(n_576),
.C(n_570),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_L g647 ( 
.A1(n_611),
.A2(n_549),
.B(n_487),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_SL g648 ( 
.A(n_592),
.B(n_499),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_589),
.B(n_545),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_590),
.A2(n_593),
.B(n_592),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_566),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_573),
.B(n_540),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_550),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_593),
.A2(n_528),
.B(n_499),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_550),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_583),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_571),
.B(n_542),
.Y(n_657)
);

NOR2x1p5_ASAP7_75t_SL g658 ( 
.A(n_558),
.B(n_499),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_573),
.A2(n_569),
.B(n_609),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_609),
.A2(n_528),
.B1(n_518),
.B2(n_124),
.Y(n_660)
);

BUFx8_ASAP7_75t_L g661 ( 
.A(n_579),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_610),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_580),
.B(n_14),
.C(n_15),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_591),
.A2(n_518),
.B(n_17),
.C(n_18),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_SL g665 ( 
.A1(n_606),
.A2(n_518),
.B(n_127),
.C(n_128),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_555),
.A2(n_126),
.B(n_208),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_614),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_557),
.A2(n_574),
.B(n_577),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_567),
.B(n_16),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_567),
.B(n_584),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_588),
.A2(n_122),
.B(n_202),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_596),
.A2(n_121),
.B(n_201),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_567),
.Y(n_673)
);

O2A1O1Ixp5_ASAP7_75t_L g674 ( 
.A1(n_585),
.A2(n_608),
.B(n_602),
.C(n_586),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_16),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_575),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_624),
.A2(n_604),
.B(n_608),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_645),
.Y(n_678)
);

NOR2xp67_ASAP7_75t_SL g679 ( 
.A(n_667),
.B(n_614),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_617),
.B(n_582),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_618),
.B(n_608),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_644),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_632),
.A2(n_608),
.B(n_578),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_622),
.A2(n_575),
.B(n_578),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_647),
.B(n_582),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_619),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_659),
.A2(n_17),
.B(n_19),
.C(n_20),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_661),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_621),
.A2(n_131),
.B(n_200),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_649),
.B(n_50),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_656),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_SL g692 ( 
.A1(n_672),
.A2(n_120),
.B(n_199),
.C(n_197),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_619),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_619),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_646),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_643),
.B(n_22),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_641),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_652),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_663),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_637),
.B(n_51),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_629),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_626),
.A2(n_52),
.B(n_54),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_657),
.B(n_55),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_653),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_630),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_631),
.B(n_57),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_661),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_SL g708 ( 
.A(n_633),
.B(n_623),
.C(n_662),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_638),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_639),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_670),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_675),
.A2(n_665),
.B(n_664),
.C(n_669),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_673),
.B(n_66),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_676),
.B(n_68),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_651),
.B(n_69),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_653),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_660),
.B(n_70),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_653),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_655),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_625),
.B(n_72),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_655),
.B(n_73),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_634),
.A2(n_74),
.B(n_75),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_627),
.A2(n_76),
.B(n_77),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_642),
.B(n_78),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_628),
.A2(n_79),
.B(n_80),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_640),
.A2(n_83),
.B(n_85),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_636),
.B(n_86),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_668),
.B(n_87),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_650),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_672),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_635),
.B(n_654),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_666),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_620),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_716),
.Y(n_734)
);

BUFx2_ASAP7_75t_SL g735 ( 
.A(n_688),
.Y(n_735)
);

BUFx6f_ASAP7_75t_SL g736 ( 
.A(n_693),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_710),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_701),
.Y(n_738)
);

BUFx2_ASAP7_75t_SL g739 ( 
.A(n_686),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_693),
.Y(n_740)
);

BUFx12f_ASAP7_75t_L g741 ( 
.A(n_707),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_693),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_704),
.Y(n_743)
);

BUFx5_ASAP7_75t_L g744 ( 
.A(n_728),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_704),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_681),
.B(n_648),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_730),
.B(n_658),
.Y(n_747)
);

BUFx5_ASAP7_75t_L g748 ( 
.A(n_678),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_704),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_686),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_691),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_718),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_711),
.B(n_671),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_719),
.Y(n_754)
);

BUFx8_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_719),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_682),
.B(n_674),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_705),
.Y(n_758)
);

INVx5_ASAP7_75t_L g759 ( 
.A(n_719),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_721),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_700),
.B(n_97),
.Y(n_761)
);

BUFx12f_ASAP7_75t_L g762 ( 
.A(n_690),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_694),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_714),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_694),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_713),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_690),
.B(n_103),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_703),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_684),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_729),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_715),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_680),
.B(n_104),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_724),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_679),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_687),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_685),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_698),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_698),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_677),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_683),
.B(n_105),
.Y(n_783)
);

BUFx12f_ASAP7_75t_L g784 ( 
.A(n_697),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_695),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_720),
.B(n_107),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_706),
.B(n_108),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_699),
.B(n_111),
.Y(n_788)
);

BUFx4f_ASAP7_75t_L g789 ( 
.A(n_717),
.Y(n_789)
);

BUFx12f_ASAP7_75t_L g790 ( 
.A(n_699),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_712),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_708),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_733),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_725),
.Y(n_794)
);

AO31x2_ASAP7_75t_L g795 ( 
.A1(n_769),
.A2(n_732),
.A3(n_689),
.B(n_726),
.Y(n_795)
);

NAND2x1p5_ASAP7_75t_L g796 ( 
.A(n_789),
.B(n_722),
.Y(n_796)
);

CKINVDCx16_ASAP7_75t_R g797 ( 
.A(n_737),
.Y(n_797)
);

OAI21x1_ASAP7_75t_L g798 ( 
.A1(n_794),
.A2(n_702),
.B(n_723),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_751),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_789),
.B(n_692),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_774),
.A2(n_116),
.B(n_117),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_766),
.B(n_760),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_776),
.B(n_119),
.Y(n_803)
);

OAI21x1_ASAP7_75t_SL g804 ( 
.A1(n_778),
.A2(n_133),
.B(n_134),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_742),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_785),
.A2(n_135),
.B(n_136),
.Y(n_806)
);

AO31x2_ASAP7_75t_L g807 ( 
.A1(n_793),
.A2(n_137),
.A3(n_138),
.B(n_139),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_738),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_763),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_736),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_787),
.A2(n_140),
.B(n_141),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_771),
.B(n_143),
.Y(n_812)
);

NAND2x1p5_ASAP7_75t_L g813 ( 
.A(n_783),
.B(n_773),
.Y(n_813)
);

AOI221xp5_ASAP7_75t_L g814 ( 
.A1(n_779),
.A2(n_144),
.B1(n_146),
.B2(n_148),
.C(n_149),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_780),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_758),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_764),
.B(n_153),
.Y(n_817)
);

AOI221xp5_ASAP7_75t_L g818 ( 
.A1(n_788),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.C(n_157),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_774),
.A2(n_158),
.B(n_159),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_746),
.B(n_161),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_765),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_SL g822 ( 
.A(n_768),
.B(n_163),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_768),
.B(n_164),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_746),
.B(n_166),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_747),
.B(n_167),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_757),
.A2(n_168),
.B(n_170),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_752),
.Y(n_828)
);

BUFx4_ASAP7_75t_SL g829 ( 
.A(n_756),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_748),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_790),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_752),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_762),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_755),
.B(n_174),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_757),
.A2(n_753),
.B(n_747),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_753),
.A2(n_175),
.B(n_176),
.Y(n_836)
);

INVx6_ASAP7_75t_SL g837 ( 
.A(n_767),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_748),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_787),
.A2(n_178),
.B(n_180),
.C(n_181),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_748),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_743),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_770),
.B(n_182),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_786),
.A2(n_792),
.B(n_754),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_786),
.A2(n_184),
.B(n_185),
.Y(n_844)
);

OA21x2_ASAP7_75t_L g845 ( 
.A1(n_782),
.A2(n_186),
.B(n_189),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_792),
.A2(n_191),
.B(n_192),
.Y(n_846)
);

OA21x2_ASAP7_75t_L g847 ( 
.A1(n_782),
.A2(n_193),
.B(n_194),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_832),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_828),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_799),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_813),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_838),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_813),
.Y(n_853)
);

OA21x2_ASAP7_75t_L g854 ( 
.A1(n_835),
.A2(n_783),
.B(n_772),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_808),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_827),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_800),
.A2(n_761),
.B(n_767),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_810),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_828),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_819),
.A2(n_791),
.B(n_748),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_830),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_840),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_816),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_811),
.A2(n_784),
.B1(n_777),
.B2(n_781),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_811),
.A2(n_772),
.B1(n_773),
.B2(n_755),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_802),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_843),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_809),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_798),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_809),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_797),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_845),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_796),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_845),
.B(n_773),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_812),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_847),
.Y(n_878)
);

BUFx4f_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_818),
.A2(n_744),
.B1(n_775),
.B2(n_735),
.Y(n_880)
);

OAI22xp33_ASAP7_75t_R g881 ( 
.A1(n_834),
.A2(n_734),
.B1(n_775),
.B2(n_741),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_826),
.A2(n_754),
.B(n_744),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_807),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_817),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_810),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_817),
.Y(n_887)
);

AOI21xp33_ASAP7_75t_L g888 ( 
.A1(n_806),
.A2(n_734),
.B(n_763),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_801),
.A2(n_744),
.B(n_745),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_842),
.Y(n_890)
);

BUFx2_ASAP7_75t_SL g891 ( 
.A(n_886),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_864),
.B(n_806),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_855),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_855),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_855),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_856),
.B(n_795),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_849),
.B(n_820),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_856),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_859),
.B(n_824),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_852),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_873),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_856),
.B(n_795),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_852),
.B(n_795),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_SL g904 ( 
.A(n_866),
.B(n_833),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_R g905 ( 
.A(n_854),
.B(n_805),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_858),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_850),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_853),
.B(n_841),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_852),
.B(n_825),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_858),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_871),
.A2(n_819),
.B(n_804),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_L g912 ( 
.A(n_890),
.B(n_818),
.C(n_814),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_850),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_874),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_848),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_879),
.A2(n_814),
.B(n_822),
.C(n_839),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_880),
.A2(n_837),
.B1(n_796),
.B2(n_815),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_861),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_863),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_861),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_877),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_915),
.B(n_868),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_898),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_898),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_893),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_900),
.B(n_869),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_900),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_894),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_900),
.B(n_848),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_894),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_914),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_905),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_903),
.B(n_879),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_897),
.B(n_890),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_893),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_895),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_918),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_895),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_918),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_920),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_920),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_907),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_907),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_903),
.B(n_879),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_942),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_942),
.Y(n_946)
);

AND4x1_ASAP7_75t_L g947 ( 
.A(n_933),
.B(n_916),
.C(n_912),
.D(n_881),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_932),
.A2(n_896),
.B(n_902),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_931),
.Y(n_949)
);

OAI22xp33_ASAP7_75t_SL g950 ( 
.A1(n_934),
.A2(n_921),
.B1(n_910),
.B2(n_879),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_937),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_933),
.A2(n_892),
.B(n_888),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_938),
.A2(n_874),
.B(n_878),
.Y(n_953)
);

AOI221xp5_ASAP7_75t_L g954 ( 
.A1(n_922),
.A2(n_892),
.B1(n_904),
.B2(n_899),
.C(n_885),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_927),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_937),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_942),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_944),
.B(n_922),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_943),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_927),
.Y(n_960)
);

OAI31xp33_ASAP7_75t_L g961 ( 
.A1(n_950),
.A2(n_917),
.A3(n_944),
.B(n_906),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_949),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_949),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_958),
.B(n_929),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_953),
.Y(n_965)
);

OAI31xp33_ASAP7_75t_L g966 ( 
.A1(n_952),
.A2(n_906),
.A3(n_901),
.B(n_831),
.Y(n_966)
);

NOR2x1_ASAP7_75t_SL g967 ( 
.A(n_958),
.B(n_891),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_954),
.A2(n_921),
.B1(n_891),
.B2(n_875),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_960),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_955),
.B(n_927),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_953),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_962),
.B(n_948),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_962),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_963),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_963),
.B(n_948),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_964),
.B(n_947),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_965),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_964),
.B(n_908),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_976),
.A2(n_961),
.B(n_968),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_973),
.B(n_969),
.Y(n_980)
);

OAI31xp33_ASAP7_75t_L g981 ( 
.A1(n_972),
.A2(n_966),
.A3(n_881),
.B(n_969),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_974),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_978),
.B(n_967),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_974),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_975),
.B(n_970),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_983),
.B(n_970),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_984),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_980),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_SL g989 ( 
.A1(n_979),
.A2(n_877),
.B1(n_948),
.B2(n_875),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_985),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_985),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_981),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_981),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_984),
.B(n_948),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_980),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_980),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_987),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_987),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_991),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_990),
.B(n_986),
.Y(n_1000)
);

AND2x4_ASAP7_75t_SL g1001 ( 
.A(n_988),
.B(n_886),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_970),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_996),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_993),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_993),
.B(n_977),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_1004),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_999),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1004),
.A2(n_992),
.B1(n_989),
.B2(n_994),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_997),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_998),
.B(n_977),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1000),
.A2(n_908),
.B1(n_960),
.B2(n_877),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_1002),
.B(n_960),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1001),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1003),
.B(n_960),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_1013),
.B(n_1005),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1014),
.B(n_1005),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1006),
.B(n_960),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1012),
.B(n_955),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_1007),
.B(n_955),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_1008),
.B(n_908),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1010),
.B(n_951),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1011),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1016),
.B(n_951),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1018),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1017),
.B(n_965),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1020),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_1020),
.B(n_971),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1021),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1023),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1019),
.Y(n_1032)
);

NAND2x1_ASAP7_75t_SL g1033 ( 
.A(n_1016),
.B(n_971),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1028),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1033),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1031),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_1027),
.B(n_842),
.C(n_823),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1030),
.B(n_956),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1031),
.Y(n_1039)
);

OAI211xp5_ASAP7_75t_L g1040 ( 
.A1(n_1025),
.A2(n_829),
.B(n_750),
.C(n_749),
.Y(n_1040)
);

AOI21xp33_ASAP7_75t_SL g1041 ( 
.A1(n_1032),
.A2(n_844),
.B(n_196),
.Y(n_1041)
);

AOI211xp5_ASAP7_75t_L g1042 ( 
.A1(n_1040),
.A2(n_1026),
.B(n_1024),
.C(n_1029),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1034),
.A2(n_945),
.B(n_957),
.C(n_956),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_SL g1044 ( 
.A1(n_1036),
.A2(n_803),
.B(n_736),
.C(n_745),
.Y(n_1044)
);

AOI211xp5_ASAP7_75t_SL g1045 ( 
.A1(n_1039),
.A2(n_803),
.B(n_885),
.C(n_887),
.Y(n_1045)
);

AOI211xp5_ASAP7_75t_L g1046 ( 
.A1(n_1038),
.A2(n_846),
.B(n_887),
.C(n_876),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1035),
.Y(n_1047)
);

AOI211xp5_ASAP7_75t_SL g1048 ( 
.A1(n_1037),
.A2(n_957),
.B(n_945),
.C(n_946),
.Y(n_1048)
);

AOI211xp5_ASAP7_75t_L g1049 ( 
.A1(n_1047),
.A2(n_1041),
.B(n_926),
.C(n_959),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_1042),
.A2(n_750),
.B1(n_740),
.B2(n_749),
.Y(n_1050)
);

AOI221xp5_ASAP7_75t_L g1051 ( 
.A1(n_1043),
.A2(n_763),
.B1(n_926),
.B2(n_927),
.C(n_929),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_1046),
.A2(n_953),
.B(n_739),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_1048),
.C(n_1045),
.Y(n_1053)
);

AOI211xp5_ASAP7_75t_L g1054 ( 
.A1(n_1047),
.A2(n_876),
.B(n_878),
.C(n_851),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1047),
.B(n_923),
.Y(n_1055)
);

OAI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1047),
.A2(n_860),
.B1(n_857),
.B2(n_740),
.C(n_749),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1042),
.A2(n_884),
.B(n_865),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1047),
.B(n_759),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_SL g1059 ( 
.A1(n_1058),
.A2(n_1055),
.B(n_1052),
.C(n_1049),
.Y(n_1059)
);

AOI211xp5_ASAP7_75t_L g1060 ( 
.A1(n_1050),
.A2(n_851),
.B(n_889),
.C(n_853),
.Y(n_1060)
);

AOI221x1_ASAP7_75t_L g1061 ( 
.A1(n_1053),
.A2(n_930),
.B1(n_928),
.B2(n_936),
.C(n_938),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_L g1062 ( 
.A(n_1054),
.B(n_759),
.C(n_749),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1057),
.A2(n_860),
.B(n_889),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_1056),
.B(n_1051),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1049),
.A2(n_837),
.B1(n_943),
.B2(n_940),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1058),
.A2(n_884),
.B(n_943),
.C(n_853),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_L g1067 ( 
.A(n_1058),
.B(n_940),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1053),
.B(n_925),
.Y(n_1068)
);

OR3x1_ASAP7_75t_L g1069 ( 
.A(n_1059),
.B(n_936),
.C(n_930),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_877),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1060),
.B(n_1067),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_SL g1072 ( 
.A(n_1064),
.B(n_740),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_1062),
.B(n_195),
.Y(n_1073)
);

OAI211xp5_ASAP7_75t_L g1074 ( 
.A1(n_1061),
.A2(n_740),
.B(n_759),
.C(n_857),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1066),
.B(n_923),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1065),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1063),
.A2(n_884),
.B(n_759),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_L g1078 ( 
.A(n_1068),
.B(n_884),
.C(n_882),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1068),
.Y(n_1079)
);

XNOR2x1_ASAP7_75t_L g1080 ( 
.A(n_1064),
.B(n_210),
.Y(n_1080)
);

AOI322xp5_ASAP7_75t_L g1081 ( 
.A1(n_1068),
.A2(n_928),
.A3(n_937),
.B1(n_940),
.B2(n_941),
.C1(n_939),
.C2(n_872),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1069),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1080),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1070),
.B(n_872),
.Y(n_1084)
);

CKINVDCx6p67_ASAP7_75t_R g1085 ( 
.A(n_1079),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_1076),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1072),
.A2(n_851),
.B1(n_870),
.B2(n_854),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1073),
.B(n_851),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1071),
.Y(n_1089)
);

AND3x1_ASAP7_75t_L g1090 ( 
.A(n_1077),
.B(n_940),
.C(n_937),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1089),
.A2(n_1075),
.B(n_1078),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1086),
.A2(n_1074),
.B1(n_1081),
.B2(n_935),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_1082),
.B(n_941),
.C(n_939),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_SL g1094 ( 
.A(n_1083),
.B(n_851),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1088),
.A2(n_870),
.B1(n_923),
.B2(n_935),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1085),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1084),
.Y(n_1097)
);

OAI22x1_ASAP7_75t_L g1098 ( 
.A1(n_1090),
.A2(n_925),
.B1(n_935),
.B2(n_938),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_1096),
.B(n_1087),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_925),
.B1(n_851),
.B2(n_924),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1094),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_1099),
.Y(n_1102)
);

AOI22x1_ASAP7_75t_L g1103 ( 
.A1(n_1102),
.A2(n_1101),
.B1(n_1091),
.B2(n_1095),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1103),
.B(n_1092),
.Y(n_1104)
);

BUFx2_ASAP7_75t_SL g1105 ( 
.A(n_1104),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1104),
.A2(n_1093),
.B1(n_1100),
.B2(n_1098),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1105),
.Y(n_1107)
);

OAI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1106),
.A2(n_924),
.B1(n_919),
.B2(n_913),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1107),
.A2(n_909),
.B1(n_883),
.B2(n_919),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1108),
.A2(n_911),
.B1(n_865),
.B2(n_883),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_1109),
.B(n_882),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_1110),
.B(n_909),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_1111),
.B1(n_911),
.B2(n_862),
.Y(n_1113)
);

AOI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_913),
.B(n_863),
.C(n_867),
.Y(n_1114)
);


endmodule