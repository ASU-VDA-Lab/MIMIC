module fake_ariane_2543_n_1824 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1824);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1824;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVxp33_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_32),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_8),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_2),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_44),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_60),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_66),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_35),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_56),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_35),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_147),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_26),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_83),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_36),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_19),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_11),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_43),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_150),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_117),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_63),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_13),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_91),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_55),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_113),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_103),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_72),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_45),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_1),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_82),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_30),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_60),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_89),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_132),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_25),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_143),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

INVxp33_ASAP7_75t_SL g248 ( 
.A(n_59),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_138),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_87),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_119),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_118),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_21),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_152),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_168),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_141),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_107),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_39),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_5),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_59),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_71),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_11),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_136),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_123),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_170),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_64),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_131),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_26),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_81),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_22),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_32),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_122),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_40),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_57),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_84),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_69),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_129),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_21),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_13),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_31),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_55),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_9),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_20),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_135),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_58),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_171),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_18),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_41),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_14),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_102),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_112),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_65),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_104),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_172),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_42),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_124),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_56),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_142),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_3),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_19),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_94),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_51),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_57),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_130),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_47),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_79),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_0),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_47),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_24),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_16),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_25),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_28),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_111),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_48),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_144),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_151),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_38),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_126),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_101),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_125),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_49),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_30),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_99),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_109),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_54),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_108),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_9),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_1),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_8),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_52),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_33),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_53),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_200),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_291),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_282),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_253),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_215),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_200),
.B(n_0),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_284),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_193),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_282),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_246),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_232),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_253),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_249),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_252),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_176),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_257),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_189),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_294),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_176),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_3),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_199),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_258),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_274),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_192),
.B(n_4),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_248),
.B(n_4),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_244),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_280),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_258),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_199),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_201),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_189),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_258),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_239),
.B(n_6),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_262),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_266),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_280),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_202),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_206),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_193),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_178),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_193),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_202),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_224),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_308),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_280),
.B(n_6),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_179),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_201),
.B(n_7),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_192),
.B(n_7),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_193),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_224),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_233),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_311),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_233),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_316),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_181),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_237),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_237),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_204),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_193),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_182),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_204),
.B(n_207),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_242),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_207),
.B(n_10),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_184),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_185),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_242),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_314),
.B(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_279),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_187),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_314),
.B(n_14),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_306),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_190),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_279),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_196),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_288),
.B(n_297),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_208),
.B(n_15),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_288),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_203),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_297),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_205),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_320),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_328),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_330),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_333),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_362),
.B(n_333),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_347),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_388),
.B(n_208),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_216),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_R g452 ( 
.A(n_344),
.B(n_209),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_366),
.B(n_338),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_352),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_380),
.B(n_174),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_344),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_394),
.B(n_338),
.C(n_191),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_368),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_385),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_351),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_348),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_387),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_377),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_405),
.B(n_303),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_410),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_369),
.B(n_177),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_369),
.B(n_375),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_384),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_392),
.B(n_303),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_398),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_345),
.B(n_216),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_409),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_422),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_354),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_426),
.B(n_330),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_415),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_346),
.B(n_306),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_429),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_424),
.B(n_217),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_430),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_431),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_371),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_364),
.B(n_306),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_357),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_395),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_428),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_385),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_435),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_458),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_477),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_374),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_484),
.B(n_350),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_477),
.B(n_353),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_462),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_375),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_444),
.B(n_365),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_435),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_477),
.B(n_367),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_462),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_477),
.B(n_358),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_458),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_484),
.A2(n_372),
.B1(n_414),
.B2(n_417),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_475),
.B(n_379),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_217),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_462),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_495),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_475),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_462),
.Y(n_539)
);

CKINVDCx11_ASAP7_75t_R g540 ( 
.A(n_468),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_492),
.B(n_379),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_492),
.B(n_484),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_495),
.B(n_507),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_469),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_506),
.B(n_358),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_469),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_435),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_506),
.B(n_360),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_435),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_475),
.B(n_360),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_469),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_438),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_475),
.B(n_407),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_484),
.B(n_356),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_495),
.B(n_383),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_475),
.B(n_407),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_478),
.B(n_411),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_460),
.B(n_373),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_506),
.B(n_411),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_450),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_484),
.B(n_177),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_468),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_478),
.B(n_412),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_450),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_433),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_468),
.B(n_416),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_461),
.A2(n_432),
.B1(n_340),
.B2(n_425),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_461),
.A2(n_425),
.B1(n_421),
.B2(n_419),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_433),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_438),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_475),
.B(n_416),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_508),
.B(n_219),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_454),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_475),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_474),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_463),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

AOI22x1_ASAP7_75t_L g594 ( 
.A1(n_504),
.A2(n_427),
.B1(n_421),
.B2(n_419),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_454),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_454),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_470),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_459),
.Y(n_599)
);

XNOR2x2_ASAP7_75t_L g600 ( 
.A(n_457),
.B(n_349),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_476),
.B(n_427),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_459),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_219),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_508),
.B(n_223),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_459),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_470),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_470),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_450),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_433),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_473),
.B(n_223),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_507),
.B(n_418),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_SL g613 ( 
.A(n_463),
.B(n_213),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_471),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_450),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_467),
.B(n_218),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_508),
.B(n_226),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_444),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_504),
.B(n_180),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_444),
.A2(n_194),
.B1(n_210),
.B2(n_222),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_479),
.B(n_355),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_479),
.B(n_508),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_467),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_493),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_433),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_498),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_444),
.A2(n_275),
.B1(n_281),
.B2(n_283),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_466),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_472),
.B(n_381),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_494),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_498),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_507),
.B(n_228),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_466),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_471),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_466),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_507),
.B(n_229),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_471),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_230),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_444),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_473),
.B(n_226),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_471),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_437),
.B(n_453),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_434),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_444),
.A2(n_275),
.B1(n_281),
.B2(n_278),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_510),
.B(n_437),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_473),
.A2(n_287),
.B1(n_276),
.B2(n_270),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_473),
.B(n_227),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_494),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_494),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_494),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_434),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_494),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_451),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_450),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_645),
.B(n_436),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_515),
.B(n_472),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_656),
.B(n_485),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_517),
.B(n_485),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_587),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_645),
.B(n_436),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_543),
.B(n_508),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_543),
.B(n_498),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_543),
.B(n_510),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_597),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_515),
.B(n_496),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_597),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_588),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_598),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_645),
.B(n_510),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_632),
.B(n_496),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_524),
.Y(n_675)
);

O2A1O1Ixp5_ASAP7_75t_L g676 ( 
.A1(n_623),
.A2(n_503),
.B(n_473),
.C(n_501),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_645),
.B(n_436),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_598),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_517),
.A2(n_488),
.B1(n_473),
.B2(n_509),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_599),
.Y(n_680)
);

BUFx5_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_543),
.B(n_501),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_537),
.B(n_619),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_632),
.B(n_503),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_SL g685 ( 
.A1(n_567),
.A2(n_391),
.B1(n_401),
.B2(n_399),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_537),
.B(n_544),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_544),
.B(n_503),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_606),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_625),
.Y(n_689)
);

AND2x6_ASAP7_75t_SL g690 ( 
.A(n_622),
.B(n_437),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_625),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_517),
.A2(n_488),
.B1(n_505),
.B2(n_509),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_606),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_607),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_628),
.B(n_503),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_565),
.B(n_574),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_538),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_633),
.B(n_503),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_542),
.B(n_361),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_538),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_599),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_538),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_607),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_648),
.B(n_493),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_602),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_602),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_648),
.B(n_529),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_605),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_638),
.B(n_493),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_514),
.B(n_363),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_538),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_524),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_632),
.B(n_436),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_SL g714 ( 
.A1(n_631),
.A2(n_382),
.B1(n_370),
.B2(n_313),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_638),
.B(n_493),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_614),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_571),
.B(n_442),
.Y(n_717)
);

AOI22x1_ASAP7_75t_L g718 ( 
.A1(n_632),
.A2(n_486),
.B1(n_481),
.B2(n_502),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_640),
.B(n_445),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_640),
.B(n_520),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_517),
.A2(n_452),
.B1(n_436),
.B2(n_502),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_601),
.B(n_488),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_533),
.B(n_488),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_605),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_511),
.B(n_488),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_560),
.B(n_487),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_625),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_535),
.B(n_488),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_611),
.Y(n_729)
);

AOI22x1_ASAP7_75t_L g730 ( 
.A1(n_644),
.A2(n_486),
.B1(n_481),
.B2(n_502),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_535),
.B(n_437),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_614),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_611),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_621),
.Y(n_734)
);

O2A1O1Ixp5_ASAP7_75t_L g735 ( 
.A1(n_564),
.A2(n_489),
.B(n_487),
.C(n_490),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_524),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_585),
.B(n_487),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_600),
.A2(n_618),
.B1(n_641),
.B2(n_518),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_621),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_636),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_645),
.B(n_453),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_626),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_535),
.B(n_517),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_524),
.A2(n_480),
.B1(n_500),
.B2(n_499),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_535),
.B(n_453),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_656),
.B(n_453),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_562),
.B(n_480),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_535),
.B(n_480),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_516),
.B(n_452),
.C(n_481),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_591),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_570),
.B(n_482),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_535),
.B(n_482),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_516),
.B(n_505),
.Y(n_753)
);

INVxp33_ASAP7_75t_L g754 ( 
.A(n_567),
.Y(n_754)
);

BUFx6f_ASAP7_75t_SL g755 ( 
.A(n_517),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_539),
.B(n_487),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_626),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_539),
.B(n_489),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_630),
.A2(n_482),
.B(n_500),
.C(n_499),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_579),
.B(n_505),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_630),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_584),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_568),
.B(n_509),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_539),
.B(n_489),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_535),
.B(n_483),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_539),
.B(n_489),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_524),
.A2(n_500),
.B1(n_499),
.B2(n_497),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_SL g768 ( 
.A(n_592),
.B(n_483),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_517),
.A2(n_497),
.B1(n_491),
.B2(n_486),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_584),
.B(n_483),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_635),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_513),
.B(n_497),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_593),
.B(n_491),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_539),
.B(n_490),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_547),
.B(n_491),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_637),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_550),
.B(n_490),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_636),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_546),
.B(n_227),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_624),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_589),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_589),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_595),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_546),
.B(n_555),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_562),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_624),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_546),
.B(n_240),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_546),
.B(n_240),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_610),
.A2(n_272),
.B1(n_265),
.B2(n_261),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_595),
.Y(n_791)
);

INVx8_ASAP7_75t_L g792 ( 
.A(n_610),
.Y(n_792)
);

NOR2x1p5_ASAP7_75t_L g793 ( 
.A(n_592),
.B(n_231),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_530),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_612),
.B(n_235),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_534),
.B(n_238),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_554),
.A2(n_307),
.B(n_247),
.C(n_250),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_616),
.B(n_634),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_616),
.B(n_245),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_580),
.B(n_254),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_586),
.A2(n_304),
.B(n_272),
.C(n_307),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_513),
.B(n_434),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_581),
.B(n_255),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_R g804 ( 
.A(n_540),
.B(n_175),
.Y(n_804)
);

AND2x2_ASAP7_75t_SL g805 ( 
.A(n_521),
.B(n_243),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_596),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_569),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_561),
.B(n_267),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_590),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_629),
.A2(n_250),
.B1(n_317),
.B2(n_265),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_613),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_591),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_546),
.B(n_243),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_726),
.A2(n_590),
.B(n_575),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_696),
.B(n_561),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_662),
.Y(n_818)
);

BUFx4f_ASAP7_75t_L g819 ( 
.A(n_660),
.Y(n_819)
);

NAND2x1p5_ASAP7_75t_L g820 ( 
.A(n_658),
.B(n_591),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_658),
.B(n_570),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_676),
.A2(n_652),
.B(n_651),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_762),
.B(n_600),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_726),
.A2(n_737),
.B(n_785),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_717),
.B(n_561),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_803),
.A2(n_652),
.B(n_655),
.C(n_651),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_707),
.A2(n_653),
.B(n_655),
.C(n_512),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_735),
.A2(n_653),
.B(n_525),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_737),
.A2(n_575),
.B(n_569),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_685),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_710),
.B(n_650),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_720),
.A2(n_583),
.B(n_512),
.C(n_558),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_793),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_683),
.A2(n_583),
.B(n_558),
.C(n_551),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_785),
.A2(n_575),
.B(n_569),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_684),
.A2(n_608),
.B(n_576),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_781),
.B(n_561),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_689),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_684),
.A2(n_608),
.B(n_576),
.Y(n_839)
);

BUFx4f_ASAP7_75t_L g840 ( 
.A(n_746),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_689),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_805),
.B(n_594),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_799),
.A2(n_649),
.B(n_532),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_759),
.A2(n_525),
.B(n_519),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_670),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_787),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_794),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_725),
.A2(n_657),
.B(n_615),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_682),
.B(n_586),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_727),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_769),
.A2(n_570),
.B1(n_586),
.B2(n_617),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_723),
.A2(n_657),
.B(n_615),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_713),
.A2(n_657),
.B(n_615),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_782),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_671),
.Y(n_855)
);

AOI21xp33_ASAP7_75t_L g856 ( 
.A1(n_661),
.A2(n_647),
.B(n_570),
.Y(n_856)
);

OAI21xp33_ASAP7_75t_L g857 ( 
.A1(n_753),
.A2(n_594),
.B(n_586),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_686),
.A2(n_566),
.B(n_549),
.C(n_522),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_727),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_786),
.B(n_620),
.Y(n_860)
);

CKINVDCx10_ASAP7_75t_R g861 ( 
.A(n_804),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_786),
.B(n_570),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_658),
.B(n_603),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_661),
.A2(n_603),
.B(n_604),
.C(n_617),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_759),
.A2(n_527),
.B(n_526),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_721),
.A2(n_541),
.B(n_527),
.Y(n_866)
);

AOI21x1_ASAP7_75t_L g867 ( 
.A1(n_756),
.A2(n_643),
.B(n_639),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_719),
.B(n_603),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_663),
.B(n_603),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_665),
.B(n_604),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_768),
.A2(n_642),
.B1(n_610),
.B2(n_604),
.Y(n_871)
);

OAI21xp33_ASAP7_75t_L g872 ( 
.A1(n_796),
.A2(n_617),
.B(n_289),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_792),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_770),
.B(n_573),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_773),
.B(n_639),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_747),
.B(n_722),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_659),
.A2(n_668),
.B(n_687),
.C(n_704),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_758),
.A2(n_548),
.B(n_545),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_747),
.B(n_610),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_663),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_758),
.A2(n_553),
.B(n_548),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_808),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_764),
.A2(n_774),
.B(n_766),
.Y(n_883)
);

AND2x2_ASAP7_75t_SL g884 ( 
.A(n_805),
.B(n_247),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_767),
.A2(n_679),
.B(n_749),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_673),
.B(n_610),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_673),
.B(n_610),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_664),
.A2(n_563),
.B(n_557),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_666),
.B(n_741),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_741),
.B(n_610),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_775),
.B(n_642),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_659),
.B(n_523),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_692),
.A2(n_643),
.B1(n_578),
.B2(n_551),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_663),
.B(n_642),
.Y(n_894)
);

CKINVDCx10_ASAP7_75t_R g895 ( 
.A(n_754),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_731),
.A2(n_563),
.B(n_549),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_745),
.A2(n_552),
.B(n_531),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_668),
.B(n_531),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_677),
.B(n_751),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_695),
.A2(n_566),
.B(n_552),
.C(n_578),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_677),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_782),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_791),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_690),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_677),
.B(n_642),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_751),
.B(n_642),
.Y(n_906)
);

AO21x1_ASAP7_75t_L g907 ( 
.A1(n_744),
.A2(n_768),
.B(n_743),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_778),
.B(n_642),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_810),
.A2(n_536),
.B(n_528),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_760),
.B(n_642),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_751),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_691),
.A2(n_559),
.B(n_572),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_791),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_680),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_709),
.B(n_572),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_800),
.A2(n_654),
.B1(n_256),
.B2(n_260),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_714),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_748),
.A2(n_559),
.B(n_654),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_701),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_715),
.B(n_559),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_697),
.A2(n_556),
.B(n_555),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_697),
.A2(n_556),
.B(n_555),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_675),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_705),
.A2(n_443),
.B(n_439),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_798),
.B(n_555),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_675),
.B(n_555),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_763),
.B(n_556),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_706),
.B(n_708),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_699),
.B(n_556),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_697),
.A2(n_609),
.B(n_582),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_SL g931 ( 
.A(n_712),
.B(n_268),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_700),
.A2(n_609),
.B(n_582),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_700),
.A2(n_609),
.B(n_582),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_724),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_712),
.B(n_582),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_L g936 ( 
.A1(n_809),
.A2(n_292),
.B(n_290),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_755),
.A2(n_323),
.B1(n_293),
.B2(n_298),
.Y(n_937)
);

O2A1O1Ixp5_ASAP7_75t_L g938 ( 
.A1(n_674),
.A2(n_256),
.B(n_317),
.C(n_304),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_752),
.A2(n_765),
.B(n_733),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_674),
.B(n_750),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_813),
.B(n_299),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_700),
.A2(n_609),
.B(n_582),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_702),
.A2(n_609),
.B(n_627),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_L g944 ( 
.A(n_795),
.B(n_448),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_750),
.B(n_300),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_728),
.Y(n_946)
);

CKINVDCx10_ASAP7_75t_R g947 ( 
.A(n_755),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_814),
.B(n_310),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_755),
.A2(n_336),
.B1(n_318),
.B2(n_319),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_736),
.B(n_321),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_792),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_811),
.B(n_325),
.Y(n_952)
);

BUFx6f_ASAP7_75t_SL g953 ( 
.A(n_736),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_808),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_792),
.A2(n_337),
.B1(n_332),
.B2(n_343),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_729),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_792),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_734),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_739),
.A2(n_339),
.B(n_341),
.C(n_342),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_808),
.B(n_814),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_702),
.A2(n_627),
.B(n_577),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_742),
.B(n_757),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_761),
.A2(n_443),
.B(n_439),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_806),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_698),
.B(n_448),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_771),
.B(n_448),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_790),
.B(n_186),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_776),
.A2(n_627),
.B(n_577),
.Y(n_968)
);

AOI21xp33_ASAP7_75t_L g969 ( 
.A1(n_797),
.A2(n_195),
.B(n_188),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_806),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_777),
.A2(n_627),
.B(n_577),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_SL g972 ( 
.A1(n_801),
.A2(n_447),
.B(n_443),
.C(n_455),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_702),
.A2(n_711),
.B(n_772),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_711),
.A2(n_627),
.B(n_577),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_681),
.B(n_577),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_783),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_667),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_801),
.A2(n_439),
.B(n_443),
.C(n_446),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_784),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_807),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_711),
.A2(n_716),
.B(n_693),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_807),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_812),
.A2(n_627),
.B(n_577),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_738),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_667),
.A2(n_703),
.B(n_693),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_817),
.A2(n_718),
.B1(n_730),
.B2(n_812),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_864),
.A2(n_694),
.B(n_703),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_847),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_876),
.A2(n_694),
.B(n_716),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_SL g990 ( 
.A(n_825),
.B(n_780),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_818),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_819),
.B(n_780),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_819),
.B(n_840),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_868),
.A2(n_740),
.B(n_672),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_977),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_840),
.B(n_738),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_846),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_849),
.A2(n_738),
.B1(n_669),
.B2(n_732),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_957),
.B(n_669),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_845),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_874),
.B(n_672),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_855),
.Y(n_1002)
);

O2A1O1Ixp5_ASAP7_75t_L g1003 ( 
.A1(n_907),
.A2(n_815),
.B(n_788),
.C(n_789),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_904),
.B(n_678),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_821),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_884),
.A2(n_681),
.B1(n_779),
.B2(n_740),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_869),
.B(n_681),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_842),
.A2(n_681),
.B1(n_779),
.B2(n_732),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_928),
.A2(n_688),
.B1(n_678),
.B2(n_802),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_917),
.B(n_688),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_823),
.B(n_681),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_848),
.A2(n_681),
.B(n_455),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_838),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_924),
.A2(n_963),
.B(n_824),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_968),
.A2(n_681),
.B(n_455),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_875),
.B(n_16),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_861),
.B(n_197),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_R g1018 ( 
.A(n_833),
.B(n_198),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_860),
.B(n_17),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_873),
.B(n_212),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_957),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_889),
.B(n_18),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_899),
.B(n_214),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_873),
.B(n_220),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_869),
.B(n_221),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_838),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_837),
.B(n_225),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_838),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_821),
.B(n_253),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_968),
.A2(n_455),
.B(n_449),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_901),
.B(n_20),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_880),
.B(n_23),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_911),
.B(n_23),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_936),
.A2(n_449),
.B(n_447),
.C(n_446),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_SL g1035 ( 
.A1(n_826),
.A2(n_449),
.B(n_447),
.C(n_446),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_854),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_914),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_SL g1038 ( 
.A1(n_941),
.A2(n_449),
.B(n_447),
.C(n_446),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_906),
.B(n_234),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_867),
.A2(n_439),
.B(n_440),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_906),
.B(n_236),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_929),
.B(n_27),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_872),
.A2(n_27),
.B(n_29),
.C(n_34),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_931),
.B(n_241),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_831),
.B(n_34),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_871),
.B(n_251),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_902),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_946),
.B(n_37),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_850),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_863),
.B(n_326),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_919),
.B(n_38),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_952),
.B(n_39),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_934),
.B(n_40),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_956),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_928),
.A2(n_312),
.B1(n_259),
.B2(n_263),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_937),
.B(n_315),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_850),
.Y(n_1057)
);

O2A1O1Ixp5_ASAP7_75t_L g1058 ( 
.A1(n_975),
.A2(n_46),
.B(n_48),
.C(n_50),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_862),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_971),
.A2(n_302),
.B(n_264),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_959),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_971),
.A2(n_305),
.B(n_269),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_903),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_913),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_850),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_937),
.B(n_309),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_857),
.A2(n_301),
.B(n_277),
.C(n_271),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_938),
.A2(n_54),
.B(n_58),
.C(n_61),
.Y(n_1068)
);

NAND2x1p5_ASAP7_75t_L g1069 ( 
.A(n_957),
.B(n_335),
.Y(n_1069)
);

CKINVDCx11_ASAP7_75t_R g1070 ( 
.A(n_895),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_822),
.A2(n_61),
.B(n_334),
.C(n_331),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_820),
.B(n_324),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_923),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_852),
.A2(n_296),
.B(n_273),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_950),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_958),
.B(n_327),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_949),
.A2(n_183),
.B(n_329),
.C(n_286),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_947),
.B(n_285),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_821),
.B(n_335),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_820),
.B(n_441),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_964),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_851),
.A2(n_183),
.B1(n_335),
.B2(n_253),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_962),
.B(n_916),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_885),
.A2(n_335),
.B(n_253),
.C(n_433),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_885),
.A2(n_335),
.B1(n_440),
.B2(n_433),
.C(n_441),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_SL g1086 ( 
.A1(n_830),
.A2(n_441),
.B1(n_440),
.B2(n_433),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_923),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_851),
.A2(n_183),
.B1(n_440),
.B2(n_433),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_SL g1089 ( 
.A1(n_891),
.A2(n_183),
.B(n_67),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_822),
.A2(n_440),
.B(n_433),
.C(n_441),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_L g1091 ( 
.A(n_841),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_976),
.Y(n_1092)
);

INVx4_ASAP7_75t_SL g1093 ( 
.A(n_953),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_973),
.A2(n_441),
.B(n_440),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_979),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_870),
.B(n_183),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_930),
.A2(n_441),
.B(n_440),
.Y(n_1097)
);

AO32x1_ASAP7_75t_L g1098 ( 
.A1(n_893),
.A2(n_183),
.A3(n_441),
.B1(n_80),
.B2(n_86),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_894),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_932),
.A2(n_62),
.B(n_78),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_951),
.B(n_90),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_841),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_890),
.A2(n_183),
.B1(n_96),
.B2(n_97),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_980),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_966),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_856),
.A2(n_183),
.B(n_106),
.C(n_110),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_953),
.Y(n_1107)
);

INVx8_ASAP7_75t_L g1108 ( 
.A(n_859),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_949),
.A2(n_183),
.B(n_115),
.C(n_120),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_945),
.A2(n_92),
.B(n_121),
.C(n_127),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_879),
.B(n_145),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_951),
.B(n_146),
.Y(n_1112)
);

AOI22x1_ASAP7_75t_L g1113 ( 
.A1(n_836),
.A2(n_148),
.B1(n_153),
.B2(n_156),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_910),
.A2(n_157),
.B1(n_165),
.B2(n_905),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_955),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_933),
.A2(n_942),
.B(n_920),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_886),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_964),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_887),
.B(n_944),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_859),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_915),
.A2(n_981),
.B(n_922),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_925),
.B(n_892),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_898),
.B(n_877),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_882),
.B(n_954),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_SL g1125 ( 
.A1(n_969),
.A2(n_935),
.B(n_984),
.C(n_926),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_921),
.A2(n_983),
.B(n_883),
.Y(n_1126)
);

CKINVDCx6p67_ASAP7_75t_R g1127 ( 
.A(n_948),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_983),
.A2(n_943),
.B(n_927),
.Y(n_1128)
);

NAND2x1_ASAP7_75t_SL g1129 ( 
.A(n_967),
.B(n_882),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_829),
.A2(n_835),
.B(n_974),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_939),
.B(n_982),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1011),
.A2(n_856),
.B(n_908),
.C(n_939),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1010),
.B(n_982),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1052),
.A2(n_982),
.B1(n_970),
.B2(n_896),
.Y(n_1134)
);

AO32x2_ASAP7_75t_L g1135 ( 
.A1(n_998),
.A2(n_893),
.A3(n_972),
.B1(n_865),
.B2(n_844),
.Y(n_1135)
);

NOR2x1_ASAP7_75t_R g1136 ( 
.A(n_1070),
.B(n_1107),
.Y(n_1136)
);

CKINVDCx11_ASAP7_75t_R g1137 ( 
.A(n_1093),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1014),
.A2(n_985),
.B(n_828),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_993),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1115),
.A2(n_940),
.B1(n_896),
.B2(n_888),
.Y(n_1140)
);

CKINVDCx6p67_ASAP7_75t_R g1141 ( 
.A(n_1057),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1059),
.B(n_970),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_988),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1105),
.B(n_970),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1056),
.A2(n_827),
.B(n_888),
.C(n_834),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_995),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1036),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1130),
.A2(n_881),
.B(n_878),
.Y(n_1148)
);

AND2x2_ASAP7_75t_SL g1149 ( 
.A(n_996),
.B(n_965),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1047),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_SL g1151 ( 
.A(n_1073),
.B(n_954),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1116),
.A2(n_866),
.B(n_844),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1031),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1032),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1066),
.B(n_960),
.Y(n_1155)
);

AOI31xp67_ASAP7_75t_L g1156 ( 
.A1(n_1008),
.A2(n_978),
.A3(n_866),
.B(n_865),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1128),
.A2(n_918),
.B(n_912),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_992),
.B(n_897),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_991),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1027),
.B(n_897),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_L g1161 ( 
.A(n_1021),
.B(n_853),
.Y(n_1161)
);

NOR4xp25_ASAP7_75t_L g1162 ( 
.A(n_1043),
.B(n_832),
.C(n_858),
.D(n_900),
.Y(n_1162)
);

CKINVDCx11_ASAP7_75t_R g1163 ( 
.A(n_1093),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1000),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1121),
.A2(n_918),
.B(n_816),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1002),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1019),
.A2(n_839),
.B(n_909),
.C(n_961),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1015),
.A2(n_1123),
.B(n_986),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1117),
.B(n_1122),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1073),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1009),
.A2(n_1084),
.A3(n_986),
.B(n_1131),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1101),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1082),
.A2(n_1016),
.B1(n_1022),
.B2(n_1083),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1042),
.A2(n_1094),
.B(n_1012),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1073),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1037),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1067),
.A2(n_989),
.A3(n_994),
.B(n_1106),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1063),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1088),
.A2(n_1044),
.B1(n_1048),
.B2(n_1020),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1064),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1114),
.A2(n_987),
.A3(n_1096),
.B(n_1111),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1013),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_990),
.A2(n_1090),
.B(n_1035),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1005),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1054),
.B(n_1023),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1085),
.A2(n_1003),
.B(n_1030),
.Y(n_1186)
);

AOI31xp67_ASAP7_75t_L g1187 ( 
.A1(n_1103),
.A2(n_1006),
.A3(n_1046),
.B(n_1080),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1092),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1097),
.A2(n_1125),
.B(n_1100),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1095),
.B(n_1050),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1113),
.A2(n_1069),
.B(n_1034),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1074),
.A2(n_1068),
.B(n_1058),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1051),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1061),
.A2(n_1071),
.B(n_1055),
.C(n_1045),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1069),
.A2(n_999),
.B(n_1112),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1078),
.B(n_1075),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1118),
.A2(n_1001),
.A3(n_1053),
.B(n_1055),
.Y(n_1197)
);

AO21x1_ASAP7_75t_L g1198 ( 
.A1(n_1074),
.A2(n_1109),
.B(n_1077),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1013),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1033),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1129),
.A2(n_1089),
.B(n_1119),
.C(n_1060),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1062),
.A2(n_1110),
.B(n_1038),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1087),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1017),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1093),
.B(n_1087),
.Y(n_1205)
);

INVx3_ASAP7_75t_SL g1206 ( 
.A(n_1127),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1101),
.A2(n_1029),
.B1(n_1079),
.B2(n_1091),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1098),
.A2(n_1007),
.B(n_1091),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1102),
.Y(n_1209)
);

NOR3xp33_ASAP7_75t_L g1210 ( 
.A(n_1025),
.B(n_1039),
.C(n_1041),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1098),
.A2(n_1124),
.B(n_1024),
.Y(n_1211)
);

OA22x2_ASAP7_75t_L g1212 ( 
.A1(n_1117),
.A2(n_1029),
.B1(n_1079),
.B2(n_1099),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1112),
.A2(n_1076),
.B(n_1124),
.Y(n_1213)
);

AO21x2_ASAP7_75t_L g1214 ( 
.A1(n_1072),
.A2(n_1098),
.B(n_1086),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1020),
.A2(n_1024),
.B(n_1120),
.C(n_1004),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_999),
.A2(n_1079),
.A3(n_1029),
.B(n_1101),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1120),
.B(n_1108),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1087),
.B(n_1049),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1108),
.B(n_1026),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1081),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1021),
.A2(n_1108),
.B(n_1026),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1028),
.B(n_1049),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1065),
.A2(n_696),
.B(n_676),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1018),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1011),
.A2(n_696),
.B1(n_884),
.B2(n_843),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1107),
.Y(n_1226)
);

NAND3x1_ASAP7_75t_L g1227 ( 
.A(n_1052),
.B(n_823),
.C(n_622),
.Y(n_1227)
);

INVx3_ASAP7_75t_SL g1228 ( 
.A(n_1107),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1014),
.A2(n_1126),
.B(n_1130),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1073),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1073),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_991),
.Y(n_1232)
);

AO32x2_ASAP7_75t_L g1233 ( 
.A1(n_998),
.A2(n_1086),
.A3(n_1009),
.B1(n_986),
.B2(n_1114),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1011),
.A2(n_696),
.B(n_843),
.C(n_565),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1070),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_988),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_998),
.A2(n_1009),
.A3(n_1084),
.B(n_907),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_998),
.A2(n_1009),
.A3(n_1084),
.B(n_907),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1014),
.A2(n_1126),
.B(n_1130),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1014),
.A2(n_1126),
.B(n_1130),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1011),
.A2(n_696),
.B(n_843),
.C(n_565),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1011),
.B(n_1105),
.Y(n_1244)
);

NAND2x1_ASAP7_75t_L g1245 ( 
.A(n_1124),
.B(n_1120),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1011),
.A2(n_696),
.B1(n_884),
.B2(n_817),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1011),
.A2(n_696),
.B(n_843),
.C(n_565),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1011),
.B(n_1105),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1056),
.B(n_571),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1250)
);

AOI221x1_ASAP7_75t_L g1251 ( 
.A1(n_998),
.A2(n_696),
.B1(n_738),
.B2(n_843),
.C(n_857),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1010),
.B(n_717),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1011),
.A2(n_696),
.B(n_843),
.C(n_565),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1014),
.A2(n_1126),
.B(n_1130),
.Y(n_1255)
);

NAND3x1_ASAP7_75t_L g1256 ( 
.A(n_1052),
.B(n_823),
.C(n_622),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1021),
.B(n_1120),
.Y(n_1257)
);

AOI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1040),
.A2(n_1116),
.B(n_1130),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_991),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1011),
.B(n_819),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1011),
.A2(n_696),
.B1(n_884),
.B2(n_817),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1011),
.A2(n_696),
.B(n_843),
.C(n_565),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_988),
.B(n_997),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1011),
.A2(n_755),
.B(n_864),
.Y(n_1264)
);

AND2x2_ASAP7_75t_SL g1265 ( 
.A(n_1011),
.B(n_884),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1070),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1010),
.B(n_717),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_988),
.B(n_997),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1011),
.A2(n_696),
.B1(n_884),
.B2(n_817),
.Y(n_1271)
);

OAI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1056),
.A2(n_631),
.B1(n_567),
.B2(n_823),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1011),
.A2(n_884),
.B1(n_714),
.B2(n_823),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_991),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1073),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1104),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1073),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_991),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1128),
.A2(n_661),
.B(n_696),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1249),
.A2(n_1265),
.B1(n_1271),
.B2(n_1261),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1272),
.A2(n_1273),
.B1(n_1149),
.B2(n_1246),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1159),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1137),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1225),
.A2(n_1256),
.B1(n_1227),
.B2(n_1260),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_1204),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1225),
.A2(n_1268),
.B1(n_1252),
.B2(n_1160),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1164),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1155),
.A2(n_1242),
.B1(n_1234),
.B2(n_1253),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1247),
.A2(n_1262),
.B1(n_1140),
.B2(n_1145),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1143),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_SL g1291 ( 
.A(n_1235),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1153),
.B(n_1154),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1166),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1173),
.A2(n_1179),
.B1(n_1193),
.B2(n_1153),
.Y(n_1294)
);

INVx4_ASAP7_75t_SL g1295 ( 
.A(n_1216),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1173),
.A2(n_1172),
.B1(n_1244),
.B2(n_1248),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1196),
.A2(n_1140),
.B1(n_1207),
.B2(n_1210),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1263),
.Y(n_1298)
);

BUFx8_ASAP7_75t_SL g1299 ( 
.A(n_1266),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1172),
.A2(n_1248),
.B1(n_1244),
.B2(n_1185),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1220),
.Y(n_1301)
);

INVx4_ASAP7_75t_L g1302 ( 
.A(n_1220),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1239),
.A2(n_1279),
.B(n_1269),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1169),
.B(n_1190),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1270),
.A2(n_1207),
.B1(n_1264),
.B2(n_1243),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1176),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1188),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1232),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1259),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1200),
.A2(n_1251),
.B1(n_1169),
.B2(n_1278),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1212),
.A2(n_1133),
.B1(n_1178),
.B2(n_1147),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1146),
.A2(n_1150),
.B1(n_1180),
.B2(n_1276),
.Y(n_1312)
);

CKINVDCx6p67_ASAP7_75t_R g1313 ( 
.A(n_1206),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1218),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1205),
.A2(n_1224),
.B1(n_1226),
.B2(n_1209),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1228),
.A2(n_1136),
.B1(n_1213),
.B2(n_1274),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1198),
.A2(n_1184),
.B1(n_1158),
.B2(n_1142),
.Y(n_1317)
);

CKINVDCx6p67_ASAP7_75t_R g1318 ( 
.A(n_1163),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1144),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1214),
.A2(n_1192),
.B1(n_1213),
.B2(n_1233),
.Y(n_1320)
);

BUFx4f_ASAP7_75t_SL g1321 ( 
.A(n_1139),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1141),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1144),
.A2(n_1152),
.B1(n_1223),
.B2(n_1245),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1182),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1134),
.A2(n_1151),
.B1(n_1214),
.B2(n_1215),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1192),
.A2(n_1233),
.B1(n_1152),
.B2(n_1186),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1250),
.A2(n_1267),
.B1(n_1254),
.B2(n_1132),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1139),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1194),
.A2(n_1168),
.B1(n_1223),
.B2(n_1211),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1217),
.A2(n_1208),
.B1(n_1201),
.B2(n_1257),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1170),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1186),
.A2(n_1175),
.B1(n_1275),
.B2(n_1170),
.Y(n_1332)
);

INVx4_ASAP7_75t_SL g1333 ( 
.A(n_1216),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1175),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_SL g1335 ( 
.A(n_1175),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1203),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1203),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1203),
.A2(n_1275),
.B1(n_1277),
.B2(n_1231),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1275),
.A2(n_1230),
.B1(n_1231),
.B2(n_1233),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1230),
.A2(n_1257),
.B1(n_1221),
.B2(n_1202),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1217),
.A2(n_1219),
.B1(n_1161),
.B2(n_1183),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1136),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1199),
.B(n_1222),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1135),
.A2(n_1202),
.B1(n_1238),
.B2(n_1237),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1216),
.Y(n_1345)
);

INVx8_ASAP7_75t_L g1346 ( 
.A(n_1195),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1187),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1197),
.Y(n_1348)
);

INVx6_ASAP7_75t_L g1349 ( 
.A(n_1162),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1135),
.A2(n_1157),
.B1(n_1165),
.B2(n_1238),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1135),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1162),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1237),
.A2(n_1238),
.B1(n_1189),
.B2(n_1191),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1237),
.A2(n_1138),
.B1(n_1156),
.B2(n_1171),
.Y(n_1354)
);

CKINVDCx11_ASAP7_75t_R g1355 ( 
.A(n_1167),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1148),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1181),
.A2(n_1177),
.B1(n_1240),
.B2(n_1229),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1174),
.Y(n_1358)
);

INVx4_ASAP7_75t_L g1359 ( 
.A(n_1241),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1255),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1181),
.A2(n_884),
.B1(n_1265),
.B2(n_1273),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1258),
.A2(n_1243),
.B(n_1239),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1159),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1159),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1159),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1159),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1197),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1139),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1249),
.A2(n_696),
.B1(n_1265),
.B2(n_1261),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1159),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1220),
.Y(n_1376)
);

BUFx8_ASAP7_75t_L g1377 ( 
.A(n_1235),
.Y(n_1377)
);

BUFx12f_ASAP7_75t_L g1378 ( 
.A(n_1137),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1225),
.A2(n_1246),
.B1(n_1271),
.B2(n_1261),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1252),
.B(n_1268),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1137),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1249),
.A2(n_696),
.B(n_1273),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1153),
.B(n_1154),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1235),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1143),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1235),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1153),
.B(n_1154),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1265),
.A2(n_884),
.B1(n_1273),
.B2(n_1272),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1249),
.A2(n_696),
.B1(n_1265),
.B2(n_1261),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1236),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1362),
.A2(n_1329),
.B(n_1358),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1346),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1295),
.B(n_1333),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1362),
.A2(n_1303),
.B(n_1327),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1355),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1295),
.B(n_1333),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1303),
.A2(n_1356),
.B(n_1353),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1394),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1304),
.B(n_1298),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1394),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1351),
.B(n_1344),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1324),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1344),
.B(n_1282),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1385),
.A2(n_1372),
.B1(n_1393),
.B2(n_1280),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1369),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1369),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1306),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1307),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_SL g1414 ( 
.A1(n_1289),
.A2(n_1288),
.B(n_1361),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1346),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1308),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1309),
.B(n_1363),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1364),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1375),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1319),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1383),
.B(n_1286),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1292),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1348),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1386),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1330),
.A2(n_1341),
.A3(n_1305),
.B(n_1359),
.Y(n_1426)
);

INVx4_ASAP7_75t_SL g1427 ( 
.A(n_1345),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1349),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1349),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1346),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1342),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1325),
.B(n_1360),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1320),
.B(n_1350),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1323),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1323),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1334),
.B(n_1317),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1345),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1350),
.B(n_1391),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1352),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1326),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1326),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1370),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1290),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1353),
.A2(n_1332),
.B(n_1354),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1310),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1389),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1354),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1314),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1339),
.B(n_1286),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1339),
.B(n_1296),
.Y(n_1450)
);

AO21x1_ASAP7_75t_L g1451 ( 
.A1(n_1380),
.A2(n_1284),
.B(n_1297),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1347),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1296),
.B(n_1294),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1357),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1357),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1299),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1332),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1294),
.B(n_1300),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1300),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1312),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1370),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1340),
.Y(n_1462)
);

AO21x1_ASAP7_75t_SL g1463 ( 
.A1(n_1340),
.A2(n_1281),
.B(n_1365),
.Y(n_1463)
);

CKINVDCx6p67_ASAP7_75t_R g1464 ( 
.A(n_1322),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1338),
.A2(n_1343),
.B(n_1311),
.Y(n_1465)
);

CKINVDCx11_ASAP7_75t_R g1466 ( 
.A(n_1387),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1365),
.A2(n_1367),
.B1(n_1371),
.B2(n_1392),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1315),
.B(n_1367),
.Y(n_1468)
);

BUFx8_ASAP7_75t_SL g1469 ( 
.A(n_1283),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1371),
.A2(n_1381),
.B1(n_1392),
.B2(n_1388),
.C(n_1382),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1370),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1321),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1402),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1423),
.B(n_1328),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1448),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1470),
.A2(n_1374),
.B1(n_1373),
.B2(n_1379),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1408),
.A2(n_1388),
.B1(n_1382),
.B2(n_1381),
.C(n_1379),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1425),
.B(n_1316),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1469),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1448),
.Y(n_1480)
);

AND2x4_ASAP7_75t_SL g1481 ( 
.A(n_1399),
.B(n_1318),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1466),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1451),
.A2(n_1384),
.B1(n_1378),
.B2(n_1313),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1464),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1464),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1421),
.B(n_1336),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1467),
.A2(n_1301),
.B1(n_1302),
.B2(n_1376),
.C(n_1337),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1409),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1453),
.A2(n_1321),
.B1(n_1335),
.B2(n_1291),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1438),
.B(n_1336),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1438),
.B(n_1337),
.Y(n_1493)
);

OR2x2_ASAP7_75t_SL g1494 ( 
.A(n_1399),
.B(n_1390),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1409),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1414),
.A2(n_1291),
.B(n_1377),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1406),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1451),
.A2(n_1331),
.B1(n_1335),
.B2(n_1377),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1427),
.B(n_1285),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1442),
.Y(n_1500)
);

AO32x2_ASAP7_75t_L g1501 ( 
.A1(n_1396),
.A2(n_1285),
.A3(n_1430),
.B1(n_1471),
.B2(n_1442),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1439),
.B(n_1422),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1462),
.A2(n_1453),
.B(n_1398),
.Y(n_1503)
);

CKINVDCx6p67_ASAP7_75t_R g1504 ( 
.A(n_1472),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_SL g1505 ( 
.A1(n_1461),
.A2(n_1471),
.B(n_1443),
.C(n_1446),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1424),
.B(n_1396),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1462),
.A2(n_1398),
.B(n_1458),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_L g1508 ( 
.A(n_1399),
.B(n_1431),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1458),
.A2(n_1433),
.B(n_1452),
.C(n_1450),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1468),
.A2(n_1399),
.B1(n_1449),
.B2(n_1450),
.Y(n_1510)
);

NOR2x1_ASAP7_75t_SL g1511 ( 
.A(n_1399),
.B(n_1463),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1411),
.B(n_1417),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1445),
.A2(n_1435),
.B(n_1434),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1419),
.B(n_1407),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1428),
.B(n_1429),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1419),
.B(n_1407),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1405),
.B(n_1429),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1452),
.A2(n_1449),
.B(n_1441),
.C(n_1440),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1405),
.B(n_1452),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1452),
.B(n_1432),
.Y(n_1520)
);

BUFx8_ASAP7_75t_SL g1521 ( 
.A(n_1456),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1397),
.B(n_1400),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1401),
.A2(n_1444),
.B(n_1435),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1414),
.A2(n_1441),
.B1(n_1440),
.B2(n_1459),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1412),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1459),
.A2(n_1454),
.B1(n_1455),
.B2(n_1463),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1397),
.B(n_1400),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1412),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1421),
.B(n_1413),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1473),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1490),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1473),
.B(n_1434),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1490),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1495),
.B(n_1413),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1477),
.A2(n_1432),
.B(n_1436),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1497),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1512),
.B(n_1514),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1495),
.B(n_1416),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1516),
.B(n_1455),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1502),
.B(n_1503),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1502),
.B(n_1416),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1523),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1503),
.B(n_1447),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1522),
.B(n_1527),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1501),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1526),
.A2(n_1460),
.B1(n_1457),
.B2(n_1465),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1519),
.B(n_1447),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1507),
.B(n_1520),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1475),
.B(n_1410),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1526),
.A2(n_1460),
.B1(n_1457),
.B2(n_1465),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1529),
.B(n_1418),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1529),
.B(n_1418),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1517),
.B(n_1395),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1488),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1525),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1491),
.B(n_1415),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1395),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1482),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1486),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1480),
.B(n_1426),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1477),
.A2(n_1432),
.B1(n_1420),
.B2(n_1403),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1487),
.B(n_1426),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1487),
.B(n_1426),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1492),
.B(n_1426),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1513),
.B(n_1426),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1549),
.B(n_1513),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1567),
.A2(n_1509),
.B(n_1505),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1530),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1531),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1560),
.B(n_1484),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1527),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1500),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1549),
.B(n_1509),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1563),
.A2(n_1476),
.B1(n_1524),
.B2(n_1536),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1531),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1545),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1532),
.B(n_1541),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1545),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1545),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1548),
.A2(n_1524),
.B1(n_1510),
.B2(n_1493),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1561),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1550),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1474),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1567),
.A2(n_1518),
.B1(n_1483),
.B2(n_1478),
.C(n_1489),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1532),
.B(n_1542),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1561),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1518),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1563),
.B(n_1498),
.C(n_1491),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1534),
.Y(n_1593)
);

INVx5_ASAP7_75t_SL g1594 ( 
.A(n_1545),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1560),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1534),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1560),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1543),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1537),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1547),
.B(n_1559),
.C(n_1565),
.D(n_1564),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1555),
.B(n_1426),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1546),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1506),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1555),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1552),
.A2(n_1515),
.B1(n_1489),
.B2(n_1437),
.Y(n_1605)
);

NAND3xp33_ASAP7_75t_L g1606 ( 
.A(n_1536),
.B(n_1505),
.C(n_1508),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1586),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1571),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1588),
.B(n_1539),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1555),
.Y(n_1612)
);

NOR2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1606),
.B(n_1479),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1578),
.Y(n_1614)
);

NAND2xp33_ASAP7_75t_R g1615 ( 
.A(n_1572),
.B(n_1485),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1562),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1571),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1604),
.B(n_1562),
.Y(n_1618)
);

NAND2xp67_ASAP7_75t_L g1619 ( 
.A(n_1586),
.B(n_1481),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1578),
.B(n_1564),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1539),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1586),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1578),
.B(n_1564),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1577),
.Y(n_1624)
);

AND2x4_ASAP7_75t_SL g1625 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1578),
.B(n_1565),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1601),
.B(n_1553),
.Y(n_1628)
);

NOR4xp25_ASAP7_75t_SL g1629 ( 
.A(n_1587),
.B(n_1558),
.C(n_1494),
.D(n_1484),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1580),
.B(n_1565),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1553),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1600),
.B(n_1554),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1577),
.B(n_1557),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1590),
.B(n_1551),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1592),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1593),
.B(n_1557),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1580),
.B(n_1566),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1590),
.B(n_1551),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1580),
.B(n_1566),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1600),
.B(n_1554),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1580),
.B(n_1603),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1598),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1598),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1613),
.A2(n_1576),
.B1(n_1591),
.B2(n_1605),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1634),
.B(n_1568),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1632),
.A2(n_1576),
.B1(n_1544),
.B2(n_1569),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1608),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1607),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1607),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1622),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1634),
.B(n_1568),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1638),
.B(n_1583),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1608),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1638),
.B(n_1589),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1617),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1594),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1622),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1624),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1614),
.B(n_1606),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1627),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1627),
.Y(n_1669)
);

NOR2xp67_ASAP7_75t_L g1670 ( 
.A(n_1614),
.B(n_1581),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1635),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1624),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1609),
.B(n_1570),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_L g1674 ( 
.A1(n_1632),
.A2(n_1641),
.B(n_1591),
.Y(n_1674)
);

NOR5xp2_ASAP7_75t_L g1675 ( 
.A(n_1629),
.B(n_1599),
.C(n_1556),
.D(n_1596),
.E(n_1593),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1625),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1633),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1625),
.B(n_1594),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1633),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1636),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1637),
.B(n_1573),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1610),
.B(n_1585),
.Y(n_1684)
);

AO21x1_ASAP7_75t_SL g1685 ( 
.A1(n_1632),
.A2(n_1574),
.B(n_1596),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1611),
.B(n_1575),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1635),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1611),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1674),
.B(n_1647),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_L g1690 ( 
.A(n_1674),
.B(n_1621),
.C(n_1597),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1685),
.B(n_1616),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1647),
.A2(n_1629),
.B1(n_1641),
.B2(n_1575),
.Y(n_1692)
);

INVxp67_ASAP7_75t_SL g1693 ( 
.A(n_1675),
.Y(n_1693)
);

XOR2xp5_ASAP7_75t_L g1694 ( 
.A(n_1646),
.B(n_1595),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1655),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.B(n_1621),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1651),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1685),
.B(n_1616),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1667),
.A2(n_1544),
.B1(n_1582),
.B2(n_1644),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1649),
.B(n_1628),
.Y(n_1701)
);

OR2x6_ASAP7_75t_L g1702 ( 
.A(n_1646),
.B(n_1595),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1656),
.B(n_1628),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1686),
.B(n_1612),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1651),
.Y(n_1705)
);

NAND4xp75_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1670),
.C(n_1683),
.D(n_1662),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1655),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1686),
.B(n_1595),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1597),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1616),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1612),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1658),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1658),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1676),
.B(n_1595),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1656),
.B(n_1628),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1655),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1660),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1676),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1660),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1688),
.B(n_1612),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1662),
.B(n_1637),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1678),
.B(n_1637),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1678),
.B(n_1640),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1661),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1706),
.B(n_1595),
.Y(n_1725)
);

OAI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1700),
.A2(n_1631),
.B1(n_1673),
.B2(n_1664),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1717),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1717),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1689),
.A2(n_1544),
.B1(n_1688),
.B2(n_1687),
.Y(n_1729)
);

OAI321xp33_ASAP7_75t_L g1730 ( 
.A1(n_1692),
.A2(n_1664),
.A3(n_1659),
.B1(n_1657),
.B2(n_1677),
.C(n_1681),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1699),
.B(n_1677),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1724),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1710),
.B(n_1682),
.Y(n_1733)
);

NOR2x1p5_ASAP7_75t_L g1734 ( 
.A(n_1706),
.B(n_1595),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1724),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_1521),
.Y(n_1736)
);

NAND2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1709),
.B(n_1670),
.Y(n_1737)
);

O2A1O1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1693),
.A2(n_1673),
.B(n_1672),
.C(n_1666),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1714),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1708),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1690),
.A2(n_1682),
.B(n_1618),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1694),
.A2(n_1644),
.B(n_1661),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1718),
.Y(n_1743)
);

AOI322xp5_ASAP7_75t_L g1744 ( 
.A1(n_1691),
.A2(n_1640),
.A3(n_1684),
.B1(n_1618),
.B2(n_1540),
.C1(n_1668),
.C2(n_1687),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1710),
.B(n_1682),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1696),
.B(n_1521),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1702),
.Y(n_1747)
);

OAI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1720),
.A2(n_1680),
.B(n_1679),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1697),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1682),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1727),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1731),
.B(n_1696),
.Y(n_1752)
);

OAI322xp33_ASAP7_75t_L g1753 ( 
.A1(n_1726),
.A2(n_1703),
.A3(n_1715),
.B1(n_1701),
.B2(n_1704),
.C1(n_1694),
.C2(n_1712),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1746),
.B(n_1702),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1731),
.B(n_1701),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1733),
.B(n_1691),
.Y(n_1756)
);

AOI32xp33_ASAP7_75t_L g1757 ( 
.A1(n_1730),
.A2(n_1698),
.A3(n_1711),
.B1(n_1703),
.B2(n_1715),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1728),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1732),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1740),
.B(n_1705),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1743),
.B(n_1713),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1735),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1749),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1750),
.Y(n_1765)
);

OAI221xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1738),
.A2(n_1744),
.B1(n_1741),
.B2(n_1748),
.C(n_1729),
.Y(n_1766)
);

AOI321xp33_ASAP7_75t_L g1767 ( 
.A1(n_1750),
.A2(n_1698),
.A3(n_1716),
.B1(n_1707),
.B2(n_1695),
.C(n_1719),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1739),
.B(n_1631),
.Y(n_1768)
);

OAI211xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1742),
.A2(n_1736),
.B(n_1734),
.C(n_1737),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1745),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1742),
.B1(n_1747),
.B2(n_1695),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1759),
.A2(n_1737),
.B1(n_1702),
.B2(n_1707),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1755),
.B(n_1721),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1761),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1754),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1766),
.A2(n_1716),
.B1(n_1687),
.B2(n_1668),
.C(n_1665),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1754),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1766),
.A2(n_1672),
.B(n_1666),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1753),
.A2(n_1679),
.B(n_1681),
.C(n_1680),
.Y(n_1779)
);

AO22x1_ASAP7_75t_L g1780 ( 
.A1(n_1765),
.A2(n_1723),
.B1(n_1722),
.B2(n_1721),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1768),
.Y(n_1781)
);

INVxp67_ASAP7_75t_SL g1782 ( 
.A(n_1759),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1778),
.B(n_1757),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1775),
.B(n_1752),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1782),
.B(n_1781),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1773),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1774),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1780),
.Y(n_1788)
);

NOR3xp33_ASAP7_75t_SL g1789 ( 
.A(n_1772),
.B(n_1769),
.C(n_1764),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1777),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_L g1791 ( 
.A(n_1771),
.B(n_1770),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1776),
.B(n_1756),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1791),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1783),
.A2(n_1668),
.B1(n_1665),
.B2(n_1758),
.Y(n_1794)
);

NAND4xp75_ASAP7_75t_L g1795 ( 
.A(n_1789),
.B(n_1760),
.C(n_1763),
.D(n_1751),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1783),
.A2(n_1767),
.B(n_1779),
.C(n_1762),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_SL g1797 ( 
.A1(n_1784),
.A2(n_1723),
.B(n_1722),
.C(n_1665),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1785),
.A2(n_1792),
.B(n_1787),
.C(n_1790),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1796),
.A2(n_1788),
.B1(n_1786),
.B2(n_1648),
.C(n_1671),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1793),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1798),
.A2(n_1671),
.B(n_1669),
.C(n_1663),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1794),
.A2(n_1669),
.B1(n_1663),
.B2(n_1654),
.C(n_1653),
.Y(n_1802)
);

AOI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1797),
.A2(n_1652),
.B(n_1648),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1795),
.A2(n_1654),
.B1(n_1653),
.B2(n_1652),
.C(n_1602),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1800),
.Y(n_1805)
);

OAI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1799),
.A2(n_1614),
.B(n_1618),
.C(n_1642),
.Y(n_1806)
);

NAND4xp75_ASAP7_75t_L g1807 ( 
.A(n_1803),
.B(n_1640),
.C(n_1642),
.D(n_1623),
.Y(n_1807)
);

XNOR2xp5_ASAP7_75t_L g1808 ( 
.A(n_1804),
.B(n_1619),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1801),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1802),
.B(n_1496),
.C(n_1631),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1805),
.B(n_1642),
.Y(n_1811)
);

NOR3xp33_ASAP7_75t_L g1812 ( 
.A(n_1807),
.B(n_1645),
.C(n_1643),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1811),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1806),
.B1(n_1808),
.B2(n_1810),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1814),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1814),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1816),
.A2(n_1812),
.B1(n_1615),
.B2(n_1504),
.Y(n_1817)
);

XOR2x2_ASAP7_75t_L g1818 ( 
.A(n_1815),
.B(n_1511),
.Y(n_1818)
);

OAI22x1_ASAP7_75t_L g1819 ( 
.A1(n_1818),
.A2(n_1630),
.B1(n_1643),
.B2(n_1639),
.Y(n_1819)
);

XNOR2xp5_ASAP7_75t_L g1820 ( 
.A(n_1819),
.B(n_1817),
.Y(n_1820)
);

OAI21x1_ASAP7_75t_L g1821 ( 
.A1(n_1820),
.A2(n_1585),
.B(n_1620),
.Y(n_1821)
);

AOI21xp33_ASAP7_75t_L g1822 ( 
.A1(n_1821),
.A2(n_1645),
.B(n_1643),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1645),
.B1(n_1635),
.B2(n_1639),
.C(n_1602),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1639),
.B(n_1623),
.C(n_1626),
.Y(n_1824)
);


endmodule