module fake_jpeg_8017_n_32 (n_3, n_2, n_1, n_0, n_4, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_15),
.C(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_15),
.B1(n_13),
.B2(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_17),
.B(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_7),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_24),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.A3(n_25),
.B1(n_21),
.B2(n_9),
.C1(n_8),
.C2(n_10),
.Y(n_29)
);

AOI21x1_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_19),
.B(n_12),
.Y(n_28)
);

AOI322xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_0),
.A3(n_1),
.B1(n_26),
.B2(n_28),
.C1(n_22),
.C2(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_31),
.Y(n_32)
);


endmodule