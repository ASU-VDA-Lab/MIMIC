module fake_jpeg_5301_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

AND2x6_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_25),
.B1(n_20),
.B2(n_26),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_59),
.B1(n_19),
.B2(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_15),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_22),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_21),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_40),
.B1(n_34),
.B2(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_56),
.B1(n_46),
.B2(n_52),
.Y(n_99)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_74),
.B1(n_76),
.B2(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_81),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_48),
.B1(n_29),
.B2(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_61),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_21),
.B(n_17),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_92),
.B1(n_99),
.B2(n_66),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_45),
.B1(n_44),
.B2(n_51),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_58),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_71),
.C(n_30),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_64),
.B1(n_69),
.B2(n_68),
.Y(n_107)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_21),
.Y(n_117)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_87),
.B1(n_90),
.B2(n_94),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_72),
.A3(n_31),
.B1(n_33),
.B2(n_55),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_120),
.B(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_23),
.C(n_30),
.Y(n_141)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_64),
.B1(n_17),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_115),
.B1(n_86),
.B2(n_85),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_84),
.B(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_118),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_41),
.B1(n_55),
.B2(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_40),
.B1(n_34),
.B2(n_57),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_99),
.B1(n_97),
.B2(n_40),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_31),
.B(n_33),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_38),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_93),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_137),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_131),
.B1(n_134),
.B2(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_125),
.B1(n_118),
.B2(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_93),
.B1(n_29),
.B2(n_33),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_136),
.B(n_24),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_111),
.B(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_102),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_116),
.C(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_0),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_12),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_112),
.A2(n_29),
.B1(n_34),
.B2(n_63),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_125),
.C(n_109),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_1),
.B(n_2),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_161),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_134),
.B1(n_131),
.B2(n_148),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_124),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_116),
.B1(n_25),
.B2(n_63),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_170),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_25),
.B(n_0),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_127),
.B(n_24),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.C(n_138),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_135),
.C(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_91),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_146),
.B(n_136),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_180),
.B(n_157),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_185),
.B1(n_152),
.B2(n_149),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_179),
.C(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_182),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_142),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_132),
.B1(n_91),
.B2(n_78),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_91),
.C(n_63),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_188),
.C(n_3),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_25),
.B1(n_78),
.B2(n_42),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_42),
.C(n_78),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_194),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_156),
.Y(n_194)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_205),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_167),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_176),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_177),
.C(n_183),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_210),
.C(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_177),
.C(n_187),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_171),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_196),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_150),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_191),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_154),
.C(n_162),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_162),
.C(n_185),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_194),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_230),
.B(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_224),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_175),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_3),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_42),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_233),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_4),
.B(n_5),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_216),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_4),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_243),
.B(n_244),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_6),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_14),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_237),
.A3(n_239),
.B1(n_242),
.B2(n_235),
.C1(n_12),
.C2(n_6),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_14),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_7),
.B(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_7),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_251),
.C(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_250),
.C(n_10),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_10),
.Y(n_254)
);


endmodule