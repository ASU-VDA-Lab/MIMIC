module fake_jpeg_13526_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_0),
.Y(n_6)
);

BUFx12_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_SL g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_17),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_5),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_13),
.A2(n_5),
.B1(n_0),
.B2(n_4),
.Y(n_19)
);

AOI22x1_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_10),
.B1(n_12),
.B2(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_10),
.B1(n_12),
.B2(n_7),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_24),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_23),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_7),
.A3(n_22),
.B1(n_9),
.B2(n_20),
.C1(n_17),
.C2(n_15),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_34),
.B(n_28),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_28),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_29),
.C(n_30),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

BUFx24_ASAP7_75t_SL g41 ( 
.A(n_35),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_42),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B(n_22),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_25),
.B(n_4),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_7),
.C(n_9),
.Y(n_47)
);


endmodule