module fake_jpeg_9944_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_0),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_11),
.B1(n_16),
.B2(n_13),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_10),
.B1(n_21),
.B2(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.C(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_39),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_30),
.B1(n_28),
.B2(n_20),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_39),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_28),
.B1(n_34),
.B2(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_44),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

AO221x1_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_43),
.B2(n_46),
.C(n_25),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI321xp33_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_42),
.A3(n_45),
.B1(n_15),
.B2(n_17),
.C(n_18),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_15),
.Y(n_56)
);

AOI31xp67_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_15),
.A3(n_6),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_18),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_58),
.C(n_6),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_7),
.B(n_3),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_4),
.Y(n_61)
);


endmodule