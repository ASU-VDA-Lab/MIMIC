module fake_aes_1833_n_1210 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1210);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1210;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_659;
wire n_432;
wire n_386;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_724;
wire n_599;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1125;
wire n_773;
wire n_847;
wire n_1097;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1094;
wire n_1169;
wire n_652;
wire n_968;
wire n_975;
wire n_303;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_1188;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_1155;
wire n_1101;
wire n_1159;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1160;
wire n_1184;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_703;
wire n_482;
wire n_415;
wire n_394;
wire n_478;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1186;
wire n_864;
wire n_1167;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_1157;
wire n_876;
wire n_986;
wire n_886;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_1206;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_1178;
wire n_1209;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_621;
wire n_666;
wire n_423;
wire n_420;
wire n_342;
wire n_799;
wire n_880;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_937;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_881;
wire n_716;
wire n_899;
wire n_806;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_1199;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_597;
wire n_349;
wire n_723;
wire n_972;
wire n_1069;
wire n_1021;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_1208;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_875;
wire n_924;
wire n_841;
wire n_947;
wire n_1043;
wire n_582;
wire n_378;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_335;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_994;
wire n_930;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_991;
wire n_515;
wire n_670;
wire n_843;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_1204;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_153), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_120), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_4), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_40), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_191), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_164), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_132), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_231), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_157), .Y(n_297) );
INVxp33_ASAP7_75t_SL g298 ( .A(n_126), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_25), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_128), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_208), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_136), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_233), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_46), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_180), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_88), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_36), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_185), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_193), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_37), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_56), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_163), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_41), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_113), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_144), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_14), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_275), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_211), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_244), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_34), .Y(n_322) );
INVxp33_ASAP7_75t_SL g323 ( .A(n_67), .Y(n_323) );
INVxp33_ASAP7_75t_L g324 ( .A(n_222), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_7), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_154), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_133), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_206), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_260), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_215), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_121), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_149), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_19), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_148), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_212), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_177), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_16), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_69), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_86), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_169), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_270), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_188), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_109), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_55), .Y(n_344) );
INVxp33_ASAP7_75t_SL g345 ( .A(n_262), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_226), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_176), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_283), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_129), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_115), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_237), .B(n_79), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_216), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_278), .Y(n_353) );
INVxp33_ASAP7_75t_L g354 ( .A(n_285), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_256), .Y(n_355) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_236), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_277), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_282), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_97), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_229), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_242), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_196), .Y(n_362) );
INVxp33_ASAP7_75t_L g363 ( .A(n_186), .Y(n_363) );
CKINVDCx14_ASAP7_75t_R g364 ( .A(n_89), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_166), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_247), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_89), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_170), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_82), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_264), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_168), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_281), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_209), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_130), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_65), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_241), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_173), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_158), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_28), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_142), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_156), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_41), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_45), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_261), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_183), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_147), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_114), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_204), .Y(n_388) );
INVxp33_ASAP7_75t_SL g389 ( .A(n_55), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_171), .Y(n_390) );
CKINVDCx14_ASAP7_75t_R g391 ( .A(n_42), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_268), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_252), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_98), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_56), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_235), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_238), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_182), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_250), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_263), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_179), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_72), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_239), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_21), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_219), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_61), .Y(n_406) );
INVxp33_ASAP7_75t_L g407 ( .A(n_66), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_155), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_11), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_214), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_100), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_65), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_20), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_131), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_101), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_112), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_162), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_174), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_27), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_284), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_85), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_11), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_2), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_232), .Y(n_424) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_234), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_127), .Y(n_426) );
CKINVDCx14_ASAP7_75t_R g427 ( .A(n_12), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_210), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_224), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_33), .Y(n_430) );
CKINVDCx14_ASAP7_75t_R g431 ( .A(n_1), .Y(n_431) );
INVxp33_ASAP7_75t_SL g432 ( .A(n_43), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_377), .B(n_0), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_315), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_315), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_300), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_350), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_300), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_305), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_364), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_299), .B(n_0), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_391), .Y(n_443) );
INVx4_ASAP7_75t_L g444 ( .A(n_359), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_305), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_308), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_407), .B(n_1), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_292), .B(n_2), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_308), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_316), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_316), .A2(n_3), .B(n_5), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_319), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_319), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_292), .B(n_5), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_315), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_320), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_315), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_320), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_369), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_321), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_321), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_326), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_315), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_290), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_299), .B(n_6), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_374), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_290), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_294), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_374), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_459), .B(n_294), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_441), .B(n_369), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_464), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_466), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_437), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_464), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_464), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_464), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_467), .Y(n_480) );
INVx4_ASAP7_75t_SL g481 ( .A(n_466), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_467), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_467), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_441), .B(n_306), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_459), .B(n_301), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g488 ( .A(n_451), .B(n_326), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_443), .B(n_324), .Y(n_489) );
AND2x6_ASAP7_75t_L g490 ( .A(n_442), .B(n_327), .Y(n_490) );
AND2x6_ASAP7_75t_L g491 ( .A(n_442), .B(n_327), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_427), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_467), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_442), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_441), .B(n_423), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
NAND3x1_ASAP7_75t_L g498 ( .A(n_433), .B(n_335), .C(n_334), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_431), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_443), .B(n_440), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_468), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_440), .B(n_354), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_442), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_468), .Y(n_505) );
NAND2xp33_ASAP7_75t_SL g506 ( .A(n_447), .B(n_329), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_437), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_436), .B(n_414), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
AND2x6_ASAP7_75t_L g510 ( .A(n_465), .B(n_334), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_468), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g512 ( .A1(n_433), .A2(n_291), .B1(n_375), .B2(n_411), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_466), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_465), .B(n_423), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_468), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_474), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_474), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_489), .B(n_447), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_473), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_490), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_474), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_494), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_475), .Y(n_523) );
INVx4_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_512), .B(n_448), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_485), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_494), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_502), .B(n_436), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_492), .B(n_438), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_503), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_507), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_499), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_485), .B(n_465), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_492), .B(n_465), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_503), .Y(n_536) );
NAND3xp33_ASAP7_75t_SL g537 ( .A(n_506), .B(n_368), .C(n_361), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_485), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_473), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_472), .B(n_438), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_485), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_496), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_496), .B(n_289), .Y(n_543) );
BUFx3_ASAP7_75t_L g544 ( .A(n_490), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_490), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_496), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_500), .B(n_439), .Y(n_547) );
AND2x6_ASAP7_75t_SL g548 ( .A(n_512), .B(n_448), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_503), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_494), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_508), .A2(n_454), .B(n_446), .C(n_449), .Y(n_552) );
AO22x1_ASAP7_75t_L g553 ( .A1(n_490), .A2(n_345), .B1(n_298), .B2(n_323), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_514), .Y(n_556) );
OR2x2_ASAP7_75t_SL g557 ( .A(n_470), .B(n_451), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_476), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_509), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_470), .B(n_445), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_509), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_509), .Y(n_562) );
OR2x6_ASAP7_75t_L g563 ( .A(n_498), .B(n_454), .Y(n_563) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_494), .B(n_451), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_490), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_491), .B(n_446), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_513), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_491), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_491), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_476), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_491), .Y(n_571) );
BUFx3_ASAP7_75t_L g572 ( .A(n_491), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_477), .Y(n_573) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_513), .Y(n_574) );
AOI21x1_ASAP7_75t_L g575 ( .A1(n_477), .A2(n_450), .B(n_449), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_513), .Y(n_576) );
OAI22xp5_ASAP7_75t_SL g577 ( .A1(n_488), .A2(n_389), .B1(n_432), .B2(n_323), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_479), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_497), .A2(n_450), .B(n_453), .C(n_452), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_479), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_480), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_491), .Y(n_582) );
AND2x6_ASAP7_75t_SL g583 ( .A(n_487), .B(n_306), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_491), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_497), .Y(n_585) );
BUFx4f_ASAP7_75t_L g586 ( .A(n_491), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_480), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_482), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_482), .Y(n_589) );
INVx4_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_510), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_510), .B(n_452), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_484), .Y(n_593) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_510), .Y(n_594) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_594), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_535), .A2(n_504), .B(n_497), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_534), .A2(n_510), .B1(n_504), .B2(n_497), .Y(n_597) );
BUFx3_ASAP7_75t_L g598 ( .A(n_594), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_594), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_584), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_584), .Y(n_601) );
OR2x6_ASAP7_75t_L g602 ( .A(n_524), .B(n_504), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_594), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_525), .B(n_504), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_560), .B(n_510), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
BUFx2_ASAP7_75t_L g608 ( .A(n_534), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_560), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_538), .A2(n_432), .B1(n_510), .B2(n_307), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_524), .B(n_484), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_590), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_532), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_563), .A2(n_510), .B1(n_453), .B2(n_458), .Y(n_614) );
BUFx6f_ASAP7_75t_SL g615 ( .A(n_524), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_594), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_520), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_528), .B(n_487), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_592), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_580), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_580), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_556), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_531), .Y(n_625) );
BUFx3_ASAP7_75t_L g626 ( .A(n_520), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_538), .A2(n_311), .B1(n_337), .B2(n_312), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_523), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_518), .B(n_498), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_525), .B(n_498), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_581), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_587), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_592), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_544), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_577), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_533), .Y(n_636) );
AND2x2_ASAP7_75t_SL g637 ( .A(n_555), .B(n_451), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_529), .A2(n_488), .B(n_493), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_572), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_546), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_547), .B(n_456), .Y(n_641) );
BUFx12f_ASAP7_75t_L g642 ( .A(n_523), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_587), .B(n_311), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_526), .B(n_488), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_590), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_588), .Y(n_646) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_526), .A2(n_363), .B(n_345), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_583), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_563), .A2(n_458), .B1(n_460), .B2(n_456), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_579), .A2(n_552), .B(n_539), .C(n_519), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_519), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_541), .B(n_460), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_537), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_553), .B(n_461), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
OR2x6_ASAP7_75t_L g656 ( .A(n_541), .B(n_488), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_539), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_SL g658 ( .A1(n_522), .A2(n_351), .B(n_462), .C(n_461), .Y(n_658) );
BUFx2_ASAP7_75t_L g659 ( .A(n_553), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_563), .A2(n_312), .B1(n_338), .B2(n_337), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_558), .A2(n_493), .B(n_505), .C(n_501), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_543), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_590), .B(n_501), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_563), .B(n_338), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_540), .B(n_462), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_558), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_570), .B(n_505), .Y(n_667) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_572), .Y(n_668) );
OR2x6_ASAP7_75t_L g669 ( .A(n_545), .B(n_314), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_570), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_555), .A2(n_451), .B1(n_515), .B2(n_511), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_516), .A2(n_515), .B(n_511), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_573), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_542), .B(n_419), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_555), .B(n_298), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_522), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_593), .B(n_419), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_522), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_527), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_578), .B(n_451), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_586), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_586), .Y(n_682) );
NAND2xp33_ASAP7_75t_L g683 ( .A(n_582), .B(n_295), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_527), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_589), .B(n_382), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_586), .Y(n_686) );
INVx8_ASAP7_75t_L g687 ( .A(n_582), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_565), .Y(n_688) );
CKINVDCx6p67_ASAP7_75t_R g689 ( .A(n_565), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_516), .A2(n_483), .B(n_471), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_568), .Y(n_691) );
INVx5_ASAP7_75t_L g692 ( .A(n_568), .Y(n_692) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_571), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_548), .B(n_383), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_571), .Y(n_695) );
OR2x6_ASAP7_75t_L g696 ( .A(n_569), .B(n_314), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_569), .B(n_322), .Y(n_697) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_566), .B(n_367), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_550), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_530), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_SL g701 ( .A1(n_517), .A2(n_340), .B(n_341), .C(n_335), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_550), .B(n_322), .Y(n_702) );
BUFx12f_ASAP7_75t_L g703 ( .A(n_591), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g704 ( .A(n_591), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_585), .A2(n_444), .B1(n_333), .B2(n_339), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_609), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_628), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_635), .B(n_585), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_604), .A2(n_564), .B1(n_359), .B2(n_379), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_630), .A2(n_564), .B1(n_359), .B2(n_409), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_595), .Y(n_712) );
NOR2x1_ASAP7_75t_SL g713 ( .A(n_669), .B(n_575), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_649), .A2(n_557), .B1(n_575), .B2(n_328), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_702), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_608), .B(n_521), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_613), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_702), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_702), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_648), .A2(n_333), .B1(n_339), .B2(n_325), .Y(n_720) );
CKINVDCx6p67_ASAP7_75t_R g721 ( .A(n_642), .Y(n_721) );
INVx3_ASAP7_75t_L g722 ( .A(n_611), .Y(n_722) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_694), .A2(n_395), .B1(n_415), .B2(n_413), .C(n_412), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_619), .B(n_421), .Y(n_724) );
CKINVDCx6p67_ASAP7_75t_R g725 ( .A(n_642), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_643), .Y(n_726) );
OAI21x1_ASAP7_75t_L g727 ( .A1(n_638), .A2(n_536), .B(n_521), .Y(n_727) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_595), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g729 ( .A(n_692), .B(n_530), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_664), .B(n_422), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_629), .A2(n_549), .B(n_536), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_627), .B(n_557), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_659), .A2(n_549), .B1(n_576), .B2(n_562), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_660), .B(n_325), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_649), .A2(n_336), .B1(n_370), .B2(n_332), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_685), .B(n_344), .Y(n_736) );
INVx2_ASAP7_75t_SL g737 ( .A(n_628), .Y(n_737) );
OR2x6_ASAP7_75t_L g738 ( .A(n_687), .B(n_304), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_621), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_622), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_611), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_651), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_657), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_610), .A2(n_336), .B1(n_370), .B2(n_332), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_602), .B(n_530), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_673), .B(n_344), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_666), .A2(n_404), .B1(n_406), .B2(n_402), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_SL g748 ( .A1(n_658), .A2(n_296), .B(n_297), .C(n_293), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_614), .A2(n_420), .B1(n_424), .B2(n_417), .Y(n_749) );
BUFx2_ASAP7_75t_SL g750 ( .A(n_615), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_670), .Y(n_751) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_696), .A2(n_430), .B1(n_317), .B2(n_394), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_674), .B(n_304), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_666), .A2(n_394), .B1(n_444), .B2(n_340), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_606), .A2(n_444), .B1(n_341), .B2(n_343), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_602), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_636), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_614), .A2(n_386), .B1(n_372), .B2(n_302), .Y(n_758) );
BUFx3_ASAP7_75t_L g759 ( .A(n_625), .Y(n_759) );
OR2x6_ASAP7_75t_L g760 ( .A(n_687), .B(n_342), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_640), .Y(n_761) );
NOR2x1_ASAP7_75t_SL g762 ( .A(n_602), .B(n_530), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_653), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_677), .B(n_6), .Y(n_764) );
OAI21xp5_ASAP7_75t_L g765 ( .A1(n_661), .A2(n_401), .B(n_399), .Y(n_765) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_623), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_607), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_616), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_652), .B(n_530), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_647), .A2(n_426), .B1(n_428), .B2(n_416), .C(n_403), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_624), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_654), .A2(n_387), .B1(n_396), .B2(n_384), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_697), .A2(n_444), .B1(n_416), .B2(n_426), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_652), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_623), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_597), .A2(n_331), .B1(n_352), .B2(n_330), .Y(n_776) );
AOI222xp33_ASAP7_75t_L g777 ( .A1(n_641), .A2(n_428), .B1(n_403), .B2(n_429), .C1(n_425), .C2(n_365), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_697), .A2(n_632), .B1(n_646), .B2(n_631), .Y(n_778) );
INVx3_ASAP7_75t_L g779 ( .A(n_693), .Y(n_779) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_595), .Y(n_780) );
OR2x6_ASAP7_75t_L g781 ( .A(n_687), .B(n_429), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_697), .Y(n_782) );
AO31x2_ASAP7_75t_L g783 ( .A1(n_661), .A2(n_463), .A3(n_455), .B(n_457), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_631), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_650), .A2(n_346), .B(n_347), .C(n_310), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_637), .A2(n_387), .B1(n_396), .B2(n_384), .Y(n_786) );
INVx4_ASAP7_75t_L g787 ( .A(n_689), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_597), .A2(n_358), .B1(n_366), .B2(n_356), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_691), .A2(n_574), .B1(n_561), .B2(n_567), .Y(n_789) );
INVx6_ASAP7_75t_L g790 ( .A(n_703), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_696), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_632), .A2(n_444), .B1(n_469), .B2(n_466), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_646), .Y(n_793) );
INVx1_ASAP7_75t_SL g794 ( .A(n_655), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_655), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_689), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_696), .A2(n_400), .B1(n_349), .B2(n_353), .Y(n_797) );
OAI22xp33_ASAP7_75t_L g798 ( .A1(n_656), .A2(n_400), .B1(n_355), .B2(n_362), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_637), .A2(n_371), .B1(n_373), .B2(n_348), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_662), .B(n_559), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_667), .A2(n_561), .B1(n_567), .B2(n_559), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_680), .A2(n_561), .B(n_559), .Y(n_802) );
AOI221x1_ASAP7_75t_L g803 ( .A1(n_650), .A2(n_469), .B1(n_466), .B2(n_378), .C(n_380), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g804 ( .A1(n_658), .A2(n_561), .B(n_559), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_665), .B(n_559), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_671), .A2(n_381), .B(n_376), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_676), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_705), .A2(n_469), .B1(n_466), .B2(n_388), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_L g809 ( .A1(n_596), .A2(n_390), .B(n_392), .C(n_385), .Y(n_809) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_705), .A2(n_410), .B1(n_393), .B2(n_397), .C(n_398), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_633), .A2(n_561), .B1(n_574), .B2(n_567), .Y(n_811) );
INVx5_ASAP7_75t_L g812 ( .A(n_595), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_679), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_656), .A2(n_574), .B1(n_567), .B2(n_303), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_678), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_620), .B(n_7), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_656), .A2(n_567), .B1(n_574), .B2(n_360), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_678), .Y(n_818) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_701), .A2(n_418), .B1(n_469), .B2(n_313), .C(n_318), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_688), .A2(n_574), .B1(n_309), .B2(n_313), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_698), .A2(n_469), .B1(n_309), .B2(n_318), .Y(n_821) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_723), .A2(n_701), .B1(n_675), .B2(n_671), .C(n_672), .Y(n_822) );
BUFx2_ASAP7_75t_L g823 ( .A(n_707), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_732), .A2(n_675), .B1(n_703), .B2(n_699), .Y(n_824) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_712), .Y(n_825) );
BUFx4f_ASAP7_75t_SL g826 ( .A(n_721), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_799), .A2(n_684), .B1(n_699), .B2(n_704), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_799), .A2(n_684), .B1(n_699), .B2(n_704), .Y(n_828) );
BUFx2_ASAP7_75t_L g829 ( .A(n_796), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_757), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_761), .Y(n_831) );
AND2x4_ASAP7_75t_L g832 ( .A(n_722), .B(n_692), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_752), .A2(n_644), .B1(n_692), .B2(n_693), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_760), .A2(n_693), .B1(n_695), .B2(n_663), .Y(n_834) );
OAI33xp33_ASAP7_75t_L g835 ( .A1(n_752), .A2(n_301), .A3(n_357), .B1(n_405), .B2(n_408), .B3(n_455), .Y(n_835) );
OR2x6_ASAP7_75t_L g836 ( .A(n_760), .B(n_695), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g837 ( .A1(n_720), .A2(n_683), .B1(n_600), .B2(n_645), .C(n_601), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_726), .B(n_695), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_767), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_717), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_760), .A2(n_601), .B1(n_605), .B2(n_600), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_766), .A2(n_690), .B(n_603), .Y(n_842) );
BUFx3_ASAP7_75t_L g843 ( .A(n_725), .Y(n_843) );
AO21x1_ASAP7_75t_L g844 ( .A1(n_798), .A2(n_463), .B(n_455), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_722), .Y(n_845) );
OR2x6_ASAP7_75t_L g846 ( .A(n_781), .B(n_618), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_742), .B(n_612), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_708), .Y(n_848) );
AO31x2_ASAP7_75t_L g849 ( .A1(n_803), .A2(n_463), .A3(n_455), .B(n_457), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_730), .A2(n_469), .B1(n_626), .B2(n_618), .C(n_634), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_736), .A2(n_469), .B1(n_639), .B2(n_634), .C(n_618), .Y(n_851) );
OAI211xp5_ASAP7_75t_L g852 ( .A1(n_720), .A2(n_463), .B(n_457), .C(n_435), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_753), .A2(n_668), .B1(n_634), .B2(n_639), .C(n_700), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_739), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_768), .Y(n_855) );
AO21x2_ASAP7_75t_L g856 ( .A1(n_806), .A2(n_483), .B(n_471), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_774), .A2(n_617), .B1(n_598), .B2(n_603), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_787), .A2(n_682), .B1(n_686), .B2(n_681), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_774), .A2(n_617), .B1(n_598), .B2(n_603), .Y(n_859) );
OAI211xp5_ASAP7_75t_L g860 ( .A1(n_777), .A2(n_435), .B(n_434), .C(n_700), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g861 ( .A1(n_770), .A2(n_435), .B(n_434), .C(n_668), .Y(n_861) );
NAND3xp33_ASAP7_75t_SL g862 ( .A(n_763), .B(n_483), .C(n_471), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_724), .A2(n_668), .B1(n_603), .B2(n_599), .C(n_434), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_734), .A2(n_599), .B1(n_435), .B2(n_495), .C(n_478), .Y(n_864) );
OR2x6_ASAP7_75t_L g865 ( .A(n_738), .B(n_8), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_738), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_866) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_709), .A2(n_435), .B1(n_495), .B2(n_478), .C(n_486), .Y(n_867) );
INVx3_ASAP7_75t_L g868 ( .A(n_741), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g869 ( .A1(n_706), .A2(n_435), .B1(n_495), .B2(n_478), .C(n_486), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_759), .B(n_9), .Y(n_870) );
AOI21xp5_ASAP7_75t_SL g871 ( .A1(n_766), .A2(n_435), .B(n_107), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_737), .A2(n_481), .B1(n_486), .B2(n_478), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g873 ( .A1(n_791), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_764), .A2(n_481), .B1(n_486), .B2(n_478), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_798), .A2(n_481), .B1(n_486), .B2(n_16), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_771), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_740), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_778), .A2(n_18), .B1(n_15), .B2(n_17), .Y(n_878) );
INVx3_ASAP7_75t_L g879 ( .A(n_741), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_784), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_750), .A2(n_18), .B1(n_15), .B2(n_17), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_802), .A2(n_481), .B(n_108), .Y(n_882) );
INVx3_ASAP7_75t_L g883 ( .A(n_745), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_778), .A2(n_22), .B1(n_19), .B2(n_21), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_804), .A2(n_110), .B(n_106), .Y(n_885) );
OA21x2_ASAP7_75t_L g886 ( .A1(n_727), .A2(n_116), .B(n_111), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_715), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_746), .B(n_26), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_718), .A2(n_26), .B1(n_27), .B2(n_29), .Y(n_889) );
AOI221xp5_ASAP7_75t_SL g890 ( .A1(n_785), .A2(n_29), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_719), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_747), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_797), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_743), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_756), .A2(n_38), .B1(n_40), .B2(n_42), .Y(n_895) );
BUFx6f_ASAP7_75t_L g896 ( .A(n_712), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_810), .A2(n_44), .B1(n_47), .B2(n_48), .C(n_49), .Y(n_897) );
AOI21xp33_ASAP7_75t_L g898 ( .A1(n_714), .A2(n_50), .B(n_51), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_710), .A2(n_50), .B(n_52), .Y(n_899) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_786), .A2(n_53), .B1(n_54), .B2(n_57), .C(n_58), .Y(n_900) );
INVx6_ASAP7_75t_L g901 ( .A(n_790), .Y(n_901) );
BUFx6f_ASAP7_75t_L g902 ( .A(n_712), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_795), .Y(n_903) );
AOI21x1_ASAP7_75t_L g904 ( .A1(n_814), .A2(n_118), .B(n_117), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_751), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_765), .A2(n_58), .B1(n_59), .B2(n_60), .C(n_61), .Y(n_906) );
NOR2x1_ASAP7_75t_SL g907 ( .A(n_812), .B(n_60), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_790), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g909 ( .A1(n_744), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_797), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_910) );
INVx3_ASAP7_75t_L g911 ( .A(n_745), .Y(n_911) );
AO31x2_ASAP7_75t_L g912 ( .A1(n_801), .A2(n_70), .A3(n_71), .B(n_72), .Y(n_912) );
AO31x2_ASAP7_75t_L g913 ( .A1(n_713), .A2(n_809), .A3(n_817), .B(n_820), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_816), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_762), .A2(n_70), .B1(n_71), .B2(n_73), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_776), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g917 ( .A1(n_735), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_775), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_813), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_794), .A2(n_77), .B1(n_80), .B2(n_81), .Y(n_920) );
NAND2xp33_ASAP7_75t_L g921 ( .A(n_812), .B(n_80), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_782), .B(n_81), .Y(n_922) );
BUFx4f_ASAP7_75t_SL g923 ( .A(n_793), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_788), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_924) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_748), .A2(n_84), .B1(n_85), .B2(n_86), .C(n_87), .Y(n_925) );
INVx8_ASAP7_75t_L g926 ( .A(n_865), .Y(n_926) );
NAND5xp2_ASAP7_75t_L g927 ( .A(n_827), .B(n_772), .C(n_819), .D(n_773), .E(n_710), .Y(n_927) );
BUFx3_ASAP7_75t_L g928 ( .A(n_826), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g929 ( .A1(n_881), .A2(n_754), .B(n_749), .C(n_821), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_880), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_830), .Y(n_931) );
AOI21xp33_ASAP7_75t_SL g932 ( .A1(n_865), .A2(n_758), .B(n_87), .Y(n_932) );
AND2x4_ASAP7_75t_L g933 ( .A(n_836), .B(n_779), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_831), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_839), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_855), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_876), .Y(n_937) );
INVx5_ASAP7_75t_L g938 ( .A(n_836), .Y(n_938) );
INVxp67_ASAP7_75t_L g939 ( .A(n_840), .Y(n_939) );
BUFx8_ASAP7_75t_L g940 ( .A(n_843), .Y(n_940) );
BUFx2_ASAP7_75t_L g941 ( .A(n_923), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_894), .B(n_711), .Y(n_942) );
NAND3xp33_ASAP7_75t_L g943 ( .A(n_890), .B(n_821), .C(n_754), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_903), .Y(n_944) );
AO21x2_ASAP7_75t_L g945 ( .A1(n_898), .A2(n_731), .B(n_769), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_848), .Y(n_946) );
OA21x2_ASAP7_75t_L g947 ( .A1(n_890), .A2(n_711), .B(n_792), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_836), .A2(n_755), .B1(n_805), .B2(n_733), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_832), .B(n_812), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g950 ( .A1(n_846), .A2(n_800), .B1(n_716), .B2(n_808), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_905), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_846), .A2(n_818), .B1(n_815), .B2(n_807), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_866), .A2(n_792), .B1(n_811), .B2(n_789), .C(n_729), .Y(n_953) );
OAI222xp33_ASAP7_75t_L g954 ( .A1(n_846), .A2(n_812), .B1(n_91), .B2(n_92), .C1(n_93), .C2(n_94), .Y(n_954) );
AOI222xp33_ASAP7_75t_L g955 ( .A1(n_878), .A2(n_90), .B1(n_92), .B2(n_93), .C1(n_94), .C2(n_95), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_854), .Y(n_956) );
AOI222xp33_ASAP7_75t_L g957 ( .A1(n_878), .A2(n_90), .B1(n_96), .B2(n_97), .C1(n_98), .C2(n_99), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_919), .Y(n_958) );
OAI21xp5_ASAP7_75t_L g959 ( .A1(n_898), .A2(n_783), .B(n_780), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_922), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_870), .B(n_99), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_829), .B(n_783), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_888), .B(n_783), .Y(n_963) );
NAND3xp33_ASAP7_75t_L g964 ( .A(n_925), .B(n_780), .C(n_728), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_847), .B(n_783), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_877), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_842), .A2(n_780), .B(n_728), .Y(n_967) );
OR2x6_ASAP7_75t_L g968 ( .A(n_833), .B(n_712), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_914), .B(n_100), .Y(n_969) );
OAI21xp33_ASAP7_75t_SL g970 ( .A1(n_899), .A2(n_780), .B(n_728), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_900), .A2(n_728), .B1(n_102), .B2(n_103), .Y(n_971) );
OAI21xp5_ASAP7_75t_L g972 ( .A1(n_822), .A2(n_101), .B(n_102), .Y(n_972) );
INVxp67_ASAP7_75t_L g973 ( .A(n_823), .Y(n_973) );
OA21x2_ASAP7_75t_L g974 ( .A1(n_885), .A2(n_202), .B(n_287), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_922), .Y(n_975) );
INVxp67_ASAP7_75t_SL g976 ( .A(n_921), .Y(n_976) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_884), .A2(n_103), .B1(n_104), .B2(n_105), .C(n_119), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_884), .Y(n_978) );
OAI221xp5_ASAP7_75t_L g979 ( .A1(n_893), .A2(n_122), .B1(n_123), .B2(n_124), .C(n_125), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_838), .B(n_288), .Y(n_980) );
OR2x2_ASAP7_75t_L g981 ( .A(n_845), .B(n_286), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_828), .A2(n_134), .B1(n_135), .B2(n_137), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_845), .B(n_138), .Y(n_983) );
OAI21xp5_ASAP7_75t_L g984 ( .A1(n_899), .A2(n_139), .B(n_140), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_868), .B(n_141), .Y(n_985) );
INVx4_ASAP7_75t_L g986 ( .A(n_908), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_912), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_879), .B(n_143), .Y(n_988) );
AOI222xp33_ASAP7_75t_L g989 ( .A1(n_906), .A2(n_145), .B1(n_146), .B2(n_150), .C1(n_151), .C2(n_152), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g990 ( .A1(n_917), .A2(n_159), .B1(n_160), .B2(n_161), .C(n_165), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_912), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_909), .A2(n_167), .B1(n_172), .B2(n_175), .C(n_178), .Y(n_992) );
OAI211xp5_ASAP7_75t_L g993 ( .A1(n_910), .A2(n_181), .B(n_184), .C(n_187), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_912), .Y(n_994) );
NAND3xp33_ASAP7_75t_L g995 ( .A(n_892), .B(n_189), .C(n_190), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_833), .A2(n_192), .B1(n_194), .B2(n_195), .Y(n_996) );
AOI33xp33_ASAP7_75t_L g997 ( .A1(n_895), .A2(n_197), .A3(n_198), .B1(n_199), .B2(n_200), .B3(n_201), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_875), .A2(n_203), .B1(n_205), .B2(n_207), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_883), .B(n_280), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_918), .A2(n_213), .B1(n_217), .B2(n_218), .C(n_220), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1001 ( .A1(n_837), .A2(n_221), .B1(n_223), .B2(n_225), .Y(n_1001) );
NAND4xp25_ASAP7_75t_SL g1002 ( .A(n_873), .B(n_227), .C(n_228), .D(n_230), .Y(n_1002) );
INVx2_ASAP7_75t_L g1003 ( .A(n_911), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_911), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_832), .B(n_918), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_907), .Y(n_1006) );
OR2x2_ASAP7_75t_SL g1007 ( .A(n_901), .B(n_240), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_849), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_920), .A2(n_243), .B1(n_245), .B2(n_246), .C(n_248), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_860), .A2(n_249), .B1(n_251), .B2(n_253), .C(n_254), .Y(n_1010) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_968), .Y(n_1011) );
NOR3xp33_ASAP7_75t_SL g1012 ( .A(n_954), .B(n_920), .C(n_852), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_931), .B(n_897), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_934), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_987), .B(n_913), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_935), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1008), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_991), .B(n_994), .Y(n_1018) );
NAND4xp25_ASAP7_75t_L g1019 ( .A(n_955), .B(n_924), .C(n_916), .D(n_891), .Y(n_1019) );
NAND2xp5_ASAP7_75t_SL g1020 ( .A(n_976), .B(n_834), .Y(n_1020) );
NAND2x1p5_ASAP7_75t_L g1021 ( .A(n_938), .B(n_825), .Y(n_1021) );
AOI221xp5_ASAP7_75t_L g1022 ( .A1(n_932), .A2(n_889), .B1(n_887), .B2(n_835), .C(n_915), .Y(n_1022) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_939), .A2(n_824), .B1(n_844), .B2(n_862), .C(n_841), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_930), .B(n_913), .Y(n_1024) );
OAI33xp33_ASAP7_75t_L g1025 ( .A1(n_962), .A2(n_859), .A3(n_857), .B1(n_913), .B2(n_849), .B3(n_861), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_936), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_937), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_951), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_967), .Y(n_1029) );
OAI31xp33_ASAP7_75t_L g1030 ( .A1(n_927), .A2(n_859), .A3(n_857), .B(n_882), .Y(n_1030) );
OAI321xp33_ASAP7_75t_L g1031 ( .A1(n_972), .A2(n_904), .A3(n_853), .B1(n_850), .B2(n_874), .C(n_851), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_965), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_944), .B(n_849), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_958), .B(n_856), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_965), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_967), .Y(n_1036) );
INVxp67_ASAP7_75t_L g1037 ( .A(n_941), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_960), .B(n_856), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_946), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_926), .A2(n_863), .B1(n_858), .B2(n_864), .Y(n_1040) );
A2O1A1Ixp33_ASAP7_75t_L g1041 ( .A1(n_977), .A2(n_867), .B(n_869), .C(n_872), .Y(n_1041) );
INVx1_ASAP7_75t_SL g1042 ( .A(n_986), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_956), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1044 ( .A1(n_973), .A2(n_871), .B1(n_886), .B2(n_896), .C(n_902), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_963), .B(n_902), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_966), .Y(n_1046) );
NOR3xp33_ASAP7_75t_L g1047 ( .A(n_927), .B(n_886), .C(n_255), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_969), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_968), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_959), .B(n_902), .Y(n_1050) );
NOR3xp33_ASAP7_75t_L g1051 ( .A(n_961), .B(n_257), .C(n_258), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_968), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_977), .A2(n_896), .B1(n_825), .B2(n_265), .C(n_266), .Y(n_1053) );
NAND3xp33_ASAP7_75t_L g1054 ( .A(n_957), .B(n_267), .C(n_269), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_959), .B(n_271), .Y(n_1055) );
INVx3_ASAP7_75t_L g1056 ( .A(n_938), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_940), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_975), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_926), .A2(n_273), .B1(n_274), .B2(n_276), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1003), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_978), .Y(n_1061) );
OAI33xp33_ASAP7_75t_L g1062 ( .A1(n_971), .A2(n_279), .A3(n_996), .B1(n_942), .B2(n_948), .B3(n_998), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1005), .B(n_1004), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_942), .Y(n_1064) );
OAI31xp33_ASAP7_75t_L g1065 ( .A1(n_929), .A2(n_1002), .A3(n_996), .B(n_1010), .Y(n_1065) );
OAI33xp33_ASAP7_75t_L g1066 ( .A1(n_948), .A2(n_998), .A3(n_1001), .B1(n_1006), .B2(n_943), .B3(n_999), .Y(n_1066) );
NOR2x1_ASAP7_75t_SL g1067 ( .A(n_938), .B(n_981), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_945), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_945), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_949), .B(n_933), .Y(n_1070) );
AOI31xp67_ASAP7_75t_L g1071 ( .A1(n_1010), .A2(n_979), .A3(n_982), .B(n_952), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_933), .B(n_938), .Y(n_1072) );
OR2x6_ASAP7_75t_L g1073 ( .A(n_984), .B(n_964), .Y(n_1073) );
NAND4xp25_ASAP7_75t_L g1074 ( .A(n_989), .B(n_1009), .C(n_1000), .D(n_992), .Y(n_1074) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_1007), .B(n_980), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_947), .B(n_970), .Y(n_1076) );
AO21x2_ASAP7_75t_L g1077 ( .A1(n_984), .A2(n_993), .B(n_950), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_988), .Y(n_1078) );
INVx3_ASAP7_75t_L g1079 ( .A(n_1029), .Y(n_1079) );
NAND2xp5_ASAP7_75t_SL g1080 ( .A(n_1065), .B(n_997), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1018), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1061), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1024), .B(n_947), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_1042), .B(n_928), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1061), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1024), .B(n_1032), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_1032), .B(n_983), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1035), .B(n_985), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g1089 ( .A(n_1037), .B(n_995), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1058), .B(n_953), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1035), .B(n_974), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1014), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1016), .B(n_990), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_1050), .B(n_1049), .Y(n_1094) );
NOR2x1_ASAP7_75t_L g1095 ( .A(n_1075), .B(n_974), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_1064), .B(n_1063), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1064), .B(n_1063), .Y(n_1097) );
NOR2xp33_ASAP7_75t_L g1098 ( .A(n_1057), .B(n_1048), .Y(n_1098) );
INVxp67_ASAP7_75t_L g1099 ( .A(n_1026), .Y(n_1099) );
INVx3_ASAP7_75t_SL g1100 ( .A(n_1056), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1015), .B(n_1018), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1034), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1027), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1028), .B(n_1043), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1015), .B(n_1050), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1033), .B(n_1076), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1033), .B(n_1076), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1039), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1045), .B(n_1038), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1017), .B(n_1052), .Y(n_1110) );
INVx1_ASAP7_75t_SL g1111 ( .A(n_1070), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_1049), .B(n_1052), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1045), .B(n_1011), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1011), .B(n_1046), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1029), .Y(n_1115) );
NOR2xp33_ASAP7_75t_L g1116 ( .A(n_1072), .B(n_1013), .Y(n_1116) );
NOR2x1_ASAP7_75t_L g1117 ( .A(n_1056), .B(n_1054), .Y(n_1117) );
NOR2x1_ASAP7_75t_L g1118 ( .A(n_1056), .B(n_1074), .Y(n_1118) );
OAI21xp5_ASAP7_75t_L g1119 ( .A1(n_1047), .A2(n_1012), .B(n_1040), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1060), .B(n_1078), .Y(n_1120) );
OAI211xp5_ASAP7_75t_L g1121 ( .A1(n_1019), .A2(n_1030), .B(n_1023), .C(n_1022), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1068), .B(n_1069), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1036), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_1055), .B(n_1036), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1068), .B(n_1077), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1126 ( .A(n_1021), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1021), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1067), .Y(n_1128) );
NOR2xp33_ASAP7_75t_L g1129 ( .A(n_1084), .B(n_1062), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1081), .B(n_1077), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1081), .B(n_1077), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1106), .B(n_1073), .Y(n_1132) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1115), .Y(n_1133) );
OAI311xp33_ASAP7_75t_L g1134 ( .A1(n_1119), .A2(n_1053), .A3(n_1059), .B1(n_1044), .C1(n_1041), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1108), .Y(n_1135) );
AND2x2_ASAP7_75t_SL g1136 ( .A(n_1124), .B(n_1051), .Y(n_1136) );
NOR2x1_ASAP7_75t_L g1137 ( .A(n_1118), .B(n_1073), .Y(n_1137) );
INVxp67_ASAP7_75t_L g1138 ( .A(n_1098), .Y(n_1138) );
INVx1_ASAP7_75t_SL g1139 ( .A(n_1100), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1106), .B(n_1073), .Y(n_1140) );
NOR4xp25_ASAP7_75t_L g1141 ( .A(n_1121), .B(n_1020), .C(n_1031), .D(n_1041), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1096), .B(n_1025), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1108), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1107), .B(n_1101), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1107), .B(n_1066), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1082), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1109), .B(n_1071), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1101), .B(n_1071), .Y(n_1148) );
OA21x2_ASAP7_75t_L g1149 ( .A1(n_1125), .A2(n_1090), .B(n_1123), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1097), .B(n_1099), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1082), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1105), .B(n_1086), .Y(n_1152) );
OAI21xp33_ASAP7_75t_L g1153 ( .A1(n_1080), .A2(n_1095), .B(n_1116), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1085), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1105), .B(n_1083), .Y(n_1155) );
HB1xp67_ASAP7_75t_L g1156 ( .A(n_1114), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1092), .Y(n_1157) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1113), .B(n_1102), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1123), .Y(n_1159) );
CKINVDCx14_ASAP7_75t_R g1160 ( .A(n_1126), .Y(n_1160) );
NOR2xp67_ASAP7_75t_L g1161 ( .A(n_1128), .B(n_1125), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1155), .B(n_1094), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1157), .Y(n_1163) );
INVx1_ASAP7_75t_SL g1164 ( .A(n_1139), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1142), .Y(n_1165) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1160), .B(n_1120), .Y(n_1166) );
INVx1_ASAP7_75t_SL g1167 ( .A(n_1150), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1158), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1144), .B(n_1124), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1145), .B(n_1148), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1171 ( .A(n_1138), .B(n_1111), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1172 ( .A(n_1156), .Y(n_1172) );
OAI32xp33_ASAP7_75t_L g1173 ( .A1(n_1147), .A2(n_1127), .A3(n_1087), .B1(n_1093), .B2(n_1104), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1142), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1145), .B(n_1102), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1158), .Y(n_1176) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1129), .B(n_1103), .Y(n_1177) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1133), .Y(n_1178) );
OAI321xp33_ASAP7_75t_L g1179 ( .A1(n_1153), .A2(n_1089), .A3(n_1110), .B1(n_1088), .B2(n_1122), .C(n_1091), .Y(n_1179) );
INVx1_ASAP7_75t_SL g1180 ( .A(n_1152), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_1141), .A2(n_1117), .B1(n_1088), .B2(n_1112), .Y(n_1181) );
O2A1O1Ixp33_ASAP7_75t_L g1182 ( .A1(n_1141), .A2(n_1079), .B(n_1112), .C(n_1134), .Y(n_1182) );
O2A1O1Ixp33_ASAP7_75t_L g1183 ( .A1(n_1134), .A2(n_1137), .B(n_1131), .C(n_1130), .Y(n_1183) );
INVx1_ASAP7_75t_SL g1184 ( .A(n_1152), .Y(n_1184) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_1136), .A2(n_1137), .B1(n_1140), .B2(n_1132), .Y(n_1185) );
XNOR2xp5_ASAP7_75t_L g1186 ( .A(n_1136), .B(n_1132), .Y(n_1186) );
NAND2xp5_ASAP7_75t_SL g1187 ( .A(n_1161), .B(n_1140), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1135), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1149), .B(n_1143), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_1177), .A2(n_1183), .B1(n_1173), .B2(n_1182), .C(n_1174), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1189), .Y(n_1191) );
NAND2xp33_ASAP7_75t_SL g1192 ( .A(n_1186), .B(n_1187), .Y(n_1192) );
NOR2x1p5_ASAP7_75t_L g1193 ( .A(n_1170), .B(n_1174), .Y(n_1193) );
NOR3xp33_ASAP7_75t_L g1194 ( .A(n_1179), .B(n_1173), .C(n_1165), .Y(n_1194) );
OAI211xp5_ASAP7_75t_L g1195 ( .A1(n_1185), .A2(n_1181), .B(n_1164), .C(n_1165), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1163), .Y(n_1196) );
XNOR2xp5_ASAP7_75t_L g1197 ( .A(n_1186), .B(n_1167), .Y(n_1197) );
AOI322xp5_ASAP7_75t_L g1198 ( .A1(n_1166), .A2(n_1180), .A3(n_1184), .B1(n_1171), .B2(n_1175), .C1(n_1176), .C2(n_1168), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1172), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1196), .Y(n_1200) );
INVxp67_ASAP7_75t_L g1201 ( .A(n_1199), .Y(n_1201) );
AOI222xp33_ASAP7_75t_L g1202 ( .A1(n_1192), .A2(n_1190), .B1(n_1195), .B2(n_1197), .C1(n_1191), .C2(n_1193), .Y(n_1202) );
OAI211xp5_ASAP7_75t_L g1203 ( .A1(n_1202), .A2(n_1198), .B(n_1194), .C(n_1191), .Y(n_1203) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1201), .B(n_1169), .Y(n_1204) );
AOI211x1_ASAP7_75t_L g1205 ( .A1(n_1203), .A2(n_1162), .B(n_1188), .C(n_1200), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1205), .B(n_1204), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_1206), .A2(n_1178), .B1(n_1146), .B2(n_1151), .Y(n_1207) );
BUFx2_ASAP7_75t_SL g1208 ( .A(n_1207), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1208), .Y(n_1209) );
AOI21xp5_ASAP7_75t_L g1210 ( .A1(n_1209), .A2(n_1154), .B(n_1159), .Y(n_1210) );
endmodule