module fake_jpeg_31981_n_383 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_383);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_383;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_49),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_23),
.B(n_9),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_50),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_58),
.B(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_71),
.Y(n_80)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_76),
.Y(n_115)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_0),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_92),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_34),
.B1(n_22),
.B2(n_37),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_108),
.B1(n_29),
.B2(n_36),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_30),
.B1(n_24),
.B2(n_40),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_87),
.A2(n_100),
.B1(n_43),
.B2(n_72),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_30),
.B1(n_40),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_30),
.B1(n_40),
.B2(n_32),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_32),
.B1(n_35),
.B2(n_21),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_0),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_35),
.B1(n_21),
.B2(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_28),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_35),
.B1(n_42),
.B2(n_38),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

CKINVDCx6p67_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_42),
.B1(n_38),
.B2(n_33),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_122),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_154),
.Y(n_163)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_50),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_128),
.Y(n_162)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_29),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_36),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_80),
.B(n_16),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_36),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_144),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_78),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_64),
.B1(n_52),
.B2(n_53),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_151),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_67),
.B1(n_77),
.B2(n_70),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_145),
.B1(n_120),
.B2(n_119),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_43),
.B1(n_54),
.B2(n_57),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_92),
.B(n_65),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_92),
.A2(n_43),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_19),
.C(n_8),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_153),
.Y(n_173)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_8),
.B1(n_18),
.B2(n_17),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_7),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_104),
.A2(n_99),
.B1(n_98),
.B2(n_109),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_82),
.A2(n_7),
.B(n_17),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_6),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_104),
.B1(n_109),
.B2(n_103),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_170),
.B(n_133),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_87),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_191),
.C(n_135),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_105),
.B(n_102),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_121),
.B1(n_125),
.B2(n_144),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_185),
.B1(n_187),
.B2(n_81),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_128),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_83),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_189),
.B1(n_154),
.B2(n_152),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_85),
.B1(n_86),
.B2(n_113),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_106),
.B1(n_86),
.B2(n_112),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_113),
.B1(n_83),
.B2(n_118),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_103),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_81),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_133),
.B(n_126),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_196),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_129),
.B1(n_127),
.B2(n_153),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_200),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_191),
.B1(n_182),
.B2(n_172),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_138),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_204),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_133),
.B1(n_81),
.B2(n_150),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_206),
.B1(n_160),
.B2(n_189),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_130),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_205),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_165),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_211),
.B(n_216),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_132),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_133),
.B(n_112),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_155),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_215),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_179),
.C(n_169),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_170),
.B(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_101),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_163),
.A2(n_123),
.B(n_101),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_171),
.B(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_124),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_233),
.B(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_163),
.B1(n_192),
.B2(n_167),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_235),
.B1(n_199),
.B2(n_198),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_243),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_181),
.B(n_173),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_234),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_164),
.B1(n_173),
.B2(n_169),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_181),
.B1(n_174),
.B2(n_185),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_197),
.B(n_209),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_242),
.A2(n_195),
.B1(n_206),
.B2(n_219),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_196),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_184),
.B(n_177),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_239),
.B(n_229),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_161),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_203),
.B(n_240),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_265),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_200),
.C(n_216),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_256),
.C(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_242),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_213),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_235),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_205),
.C(n_207),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_257),
.B(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_217),
.C(n_211),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_261),
.B(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_208),
.B(n_218),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_215),
.C(n_220),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_274),
.C(n_225),
.Y(n_288)
);

BUFx4f_ASAP7_75t_SL g263 ( 
.A(n_239),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_231),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_172),
.C(n_161),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_232),
.B(n_244),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_221),
.A2(n_197),
.B(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_271),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_204),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_183),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_182),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_262),
.C(n_258),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_288),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_230),
.B1(n_240),
.B2(n_237),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_279),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_271),
.B(n_255),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_237),
.B1(n_242),
.B2(n_238),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_248),
.A2(n_238),
.B1(n_232),
.B2(n_230),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_294),
.Y(n_299)
);

XOR2x2_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_226),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_264),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_244),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_251),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_224),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_224),
.B(n_234),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_234),
.B(n_267),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_253),
.A2(n_234),
.B1(n_222),
.B2(n_246),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_234),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_263),
.A3(n_264),
.B1(n_256),
.B2(n_257),
.C1(n_234),
.C2(n_261),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_302),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_255),
.B(n_259),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_308),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_310),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_285),
.A2(n_268),
.B(n_269),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_312),
.A2(n_296),
.B1(n_290),
.B2(n_284),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_227),
.C(n_252),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_317),
.C(n_293),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_270),
.B1(n_246),
.B2(n_227),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_287),
.B1(n_297),
.B2(n_286),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_183),
.C(n_178),
.Y(n_317)
);

BUFx12_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_330),
.C(n_307),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_325),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_306),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_323),
.A2(n_327),
.B1(n_329),
.B2(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_299),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_292),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_304),
.A2(n_280),
.B1(n_283),
.B2(n_281),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_304),
.A2(n_280),
.B1(n_283),
.B2(n_288),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_275),
.C(n_276),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_312),
.A2(n_282),
.B1(n_277),
.B2(n_178),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_282),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_301),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_320),
.A2(n_302),
.B(n_308),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_340),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_344),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_299),
.B(n_313),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_332),
.A2(n_313),
.B(n_305),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_341),
.A2(n_342),
.B(n_350),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_335),
.A2(n_317),
.B(n_314),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_346),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_326),
.B(n_309),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_326),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_310),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_349),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_316),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_330),
.B(n_303),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_327),
.B(n_311),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_323),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_354),
.B(n_357),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_346),
.B(n_329),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_356),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_338),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_318),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_361),
.A2(n_324),
.B(n_165),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_360),
.C(n_359),
.Y(n_362)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_362),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_353),
.A2(n_331),
.B1(n_322),
.B2(n_277),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_367),
.Y(n_374)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_334),
.C(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_366),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_334),
.C(n_345),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_165),
.B(n_156),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_9),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_96),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_371),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_375),
.C(n_14),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_13),
.Y(n_375)
);

OAI322xp33_ASAP7_75t_L g376 ( 
.A1(n_372),
.A2(n_5),
.A3(n_19),
.B1(n_16),
.B2(n_15),
.C1(n_14),
.C2(n_136),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

AOI21x1_ASAP7_75t_L g381 ( 
.A1(n_378),
.A2(n_379),
.B(n_374),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_335),
.C2(n_305),
.Y(n_379)
);

NOR3xp33_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_374),
.C(n_377),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_380),
.Y(n_383)
);


endmodule