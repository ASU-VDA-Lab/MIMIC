module fake_jpeg_20195_n_105 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_22),
.B1(n_14),
.B2(n_15),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx2_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_20),
.B1(n_17),
.B2(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_7),
.C(n_10),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_26),
.Y(n_49)
);

A2O1A1O1Ixp25_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_29),
.B(n_27),
.C(n_13),
.D(n_17),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_46),
.C(n_40),
.Y(n_51)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_63),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_43),
.B1(n_39),
.B2(n_44),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_16),
.B(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_1),
.B(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_11),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_11),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_60),
.B1(n_35),
.B2(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_51),
.B1(n_55),
.B2(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_53),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_52),
.C(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_50),
.B1(n_57),
.B2(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_61),
.B1(n_54),
.B2(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_70),
.B(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_85),
.B1(n_83),
.B2(n_87),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_80),
.C(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_100)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_85),
.A3(n_86),
.B1(n_76),
.B2(n_77),
.C(n_71),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_99),
.B(n_75),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_75),
.B(n_67),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_77),
.B(n_67),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_35),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);


endmodule