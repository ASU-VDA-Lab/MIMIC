module real_jpeg_25994_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_40),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_1),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_40),
.B1(n_68),
.B2(n_69),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_3),
.A2(n_10),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_3),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_3),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_3),
.A2(n_25),
.B1(n_68),
.B2(n_69),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_6),
.B(n_29),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_63),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_69),
.C(n_83),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_53),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_6),
.A2(n_107),
.B1(n_216),
.B2(n_222),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_7),
.A2(n_68),
.B1(n_69),
.B2(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_90),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_9),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_122)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_11),
.A2(n_47),
.B1(n_97),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_11),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_11),
.A2(n_47),
.B1(n_68),
.B2(n_69),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_12),
.A2(n_68),
.B1(n_69),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_76),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_68),
.B1(n_69),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_14),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_74),
.Y(n_103)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_15),
.Y(n_121)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_145),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_143),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_19),
.B(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_77),
.C(n_101),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_20),
.B(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_44),
.B2(n_45),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_23),
.B(n_44),
.C(n_60),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_24),
.Y(n_100)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_27),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_27),
.A2(n_29),
.B1(n_39),
.B2(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_36),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_28),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_94)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_34),
.B(n_62),
.C(n_64),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_30),
.B(n_63),
.CON(n_171),
.SN(n_171)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_33),
.C(n_43),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_31),
.A2(n_52),
.A3(n_55),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_57),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_48),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_48),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_48),
.A2(n_92),
.B1(n_93),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_49),
.A2(n_53),
.B1(n_161),
.B2(n_171),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_51),
.B(n_54),
.Y(n_172)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_53),
.B(n_139),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_55),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_55),
.B(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_63),
.B(n_86),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_63),
.B(n_121),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_67),
.B(n_110),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_67),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_69),
.B1(n_83),
.B2(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_68),
.B(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_73),
.A2(n_121),
.B(n_123),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_77),
.A2(n_78),
.B1(n_101),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.C(n_94),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_79),
.A2(n_80),
.B1(n_91),
.B2(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_88),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_81),
.A2(n_126),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_81),
.A2(n_178),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_81),
.A2(n_126),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_81),
.A2(n_126),
.B1(n_177),
.B2(n_198),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_94),
.B(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_101),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_106),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_107),
.A2(n_109),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_107),
.A2(n_119),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_107),
.A2(n_213),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_141),
.B2(n_142),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_129),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_124),
.B2(n_128),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_140),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_242),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_165),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_162),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_149),
.B(n_162),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_150),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_153),
.B(n_155),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_183),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_237),
.B(n_241),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_192),
.B(n_236),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_179),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_168),
.B(n_179),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.C(n_176),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_173),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_175),
.B(n_176),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_187),
.C(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_231),
.B(n_235),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_209),
.B(n_230),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_199),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_218),
.B(n_229),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_217),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_228),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_239),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);


endmodule