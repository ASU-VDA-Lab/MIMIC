module fake_jpeg_16913_n_217 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NAND2x1_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_53),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_24),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_1),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_1),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_3),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_3),
.C(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_5),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_30),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_4),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_37),
.B1(n_21),
.B2(n_20),
.Y(n_85)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_67),
.B1(n_84),
.B2(n_90),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_34),
.B(n_23),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_93),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_37),
.B1(n_21),
.B2(n_18),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_97),
.B1(n_83),
.B2(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_20),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_100),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_8),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_58),
.B1(n_41),
.B2(n_23),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_102),
.A2(n_111),
.B1(n_105),
.B2(n_119),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_103),
.B(n_73),
.Y(n_147)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_116),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_10),
.B1(n_66),
.B2(n_64),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_65),
.B(n_79),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_129),
.A3(n_68),
.B1(n_67),
.B2(n_84),
.Y(n_133)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_65),
.B(n_86),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_130),
.B(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_70),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_96),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_76),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_68),
.B(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_145),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_96),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_102),
.B1(n_127),
.B2(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_77),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_94),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_141),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_149),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_73),
.B(n_77),
.Y(n_148)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_115),
.B1(n_113),
.B2(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_155),
.B1(n_156),
.B2(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_112),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_104),
.B1(n_114),
.B2(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_117),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_102),
.A2(n_120),
.B1(n_130),
.B2(n_125),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_173),
.B(n_154),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_139),
.C(n_148),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_177),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_145),
.B(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_134),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_172),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_159),
.B1(n_135),
.B2(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_181),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_178),
.A2(n_140),
.B1(n_135),
.B2(n_141),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_173),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_178),
.A2(n_135),
.B1(n_155),
.B2(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_147),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_190),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_132),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_195),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_144),
.B(n_152),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_196),
.B(n_162),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_132),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_199),
.B(n_196),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_167),
.C(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_176),
.B1(n_182),
.B2(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_193),
.B1(n_160),
.B2(n_194),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_195),
.C(n_163),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_205),
.A2(n_199),
.B(n_204),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_168),
.B(n_165),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_209),
.A2(n_206),
.B(n_200),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_210),
.A2(n_207),
.B(n_179),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_208),
.B(n_201),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_216),
.Y(n_217)
);


endmodule