module fake_ibex_873_n_18 (n_4, n_2, n_5, n_0, n_3, n_1, n_18);

input n_4;
input n_2;
input n_5;
input n_0;
input n_3;
input n_1;

output n_18;

wire n_13;
wire n_7;
wire n_11;
wire n_17;
wire n_6;
wire n_8;
wire n_15;
wire n_14;
wire n_10;
wire n_9;
wire n_16;
wire n_12;

INVx2_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_6),
.B(n_10),
.Y(n_14)
);

OAI211xp5_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_11),
.B(n_8),
.C(n_2),
.Y(n_15)
);

AND2x4_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

AO221x2_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_15),
.Y(n_18)
);


endmodule