module fake_jpeg_21919_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_12),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_24),
.B1(n_30),
.B2(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_44),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_28),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_49),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_51),
.Y(n_52)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_12),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_23),
.C(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_54),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_42),
.B1(n_36),
.B2(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_23),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_59),
.C(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_29),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_69),
.B(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_73),
.B1(n_61),
.B2(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_79),
.B1(n_73),
.B2(n_54),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_62),
.C(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_81),
.C(n_64),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_42),
.B1(n_59),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_68),
.B1(n_32),
.B2(n_31),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_63),
.A3(n_17),
.B1(n_10),
.B2(n_8),
.C1(n_5),
.C2(n_6),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_8),
.C(n_2),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_27),
.B(n_25),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_47),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_83),
.B(n_87),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_27),
.C(n_25),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_66),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_76),
.C(n_80),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_67),
.B1(n_51),
.B2(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_67),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_92),
.C(n_25),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_80),
.B(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_84),
.B(n_85),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_16),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_96),
.B(n_22),
.C(n_21),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_22),
.C(n_21),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_98),
.B(n_19),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_0),
.B(n_2),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_19),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_3),
.Y(n_100)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.A3(n_3),
.B1(n_4),
.B2(n_7),
.C(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_4),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_18),
.Y(n_104)
);


endmodule