module real_aes_7022_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g483 ( .A1(n_0), .A2(n_147), .B(n_484), .C(n_487), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_1), .B(n_479), .Y(n_488) );
INVx1_ASAP7_75t_L g436 ( .A(n_2), .Y(n_436) );
INVx1_ASAP7_75t_L g145 ( .A(n_3), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_4), .B(n_148), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_5), .A2(n_447), .B(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_6), .A2(n_732), .B1(n_735), .B2(n_736), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_6), .Y(n_736) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_7), .A2(n_155), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_8), .A2(n_37), .B1(n_135), .B2(n_183), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_9), .B(n_155), .Y(n_163) );
AND2x6_ASAP7_75t_L g150 ( .A(n_10), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_11), .A2(n_150), .B(n_452), .C(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_12), .A2(n_41), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_12), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_13), .B(n_38), .Y(n_437) );
INVx1_ASAP7_75t_L g126 ( .A(n_14), .Y(n_126) );
INVx1_ASAP7_75t_L g129 ( .A(n_15), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_16), .B(n_131), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_17), .B(n_148), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_18), .B(n_122), .Y(n_229) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_19), .A2(n_121), .A3(n_155), .B1(n_174), .B2(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_20), .B(n_135), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_21), .B(n_122), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_22), .A2(n_57), .B1(n_135), .B2(n_183), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g185 ( .A1(n_23), .A2(n_84), .B1(n_131), .B2(n_135), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_24), .B(n_135), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_25), .A2(n_174), .B(n_452), .C(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_26), .A2(n_174), .B(n_452), .C(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_28), .B(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_29), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_29), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_30), .A2(n_447), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_31), .B(n_176), .Y(n_217) );
INVx2_ASAP7_75t_L g133 ( .A(n_32), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_33), .A2(n_450), .B(n_454), .C(n_460), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_34), .B(n_135), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_35), .B(n_176), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_36), .B(n_194), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_39), .B(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_40), .Y(n_500) );
INVx1_ASAP7_75t_L g734 ( .A(n_41), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_42), .B(n_148), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g762 ( .A1(n_43), .A2(n_763), .B1(n_765), .B2(n_766), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_43), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_44), .B(n_447), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_45), .A2(n_109), .B1(n_110), .B2(n_431), .Y(n_108) );
INVx1_ASAP7_75t_L g431 ( .A(n_45), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_45), .A2(n_47), .B1(n_431), .B2(n_764), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_46), .A2(n_450), .B(n_460), .C(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_47), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_48), .B(n_135), .Y(n_158) );
INVx1_ASAP7_75t_L g485 ( .A(n_49), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_50), .A2(n_92), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g516 ( .A(n_51), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_52), .B(n_135), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_53), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_54), .B(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_55), .B(n_447), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_56), .B(n_143), .Y(n_162) );
AOI22xp33_ASAP7_75t_SL g227 ( .A1(n_58), .A2(n_62), .B1(n_131), .B2(n_135), .Y(n_227) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_59), .A2(n_105), .B1(n_745), .B2(n_755), .C1(n_772), .C2(n_778), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_59), .Y(n_475) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_59), .A2(n_69), .B1(n_475), .B2(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_60), .B(n_135), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_61), .B(n_135), .Y(n_191) );
INVx1_ASAP7_75t_L g151 ( .A(n_63), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_64), .B(n_447), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_65), .B(n_479), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_66), .A2(n_137), .B(n_143), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_67), .B(n_135), .Y(n_146) );
INVx1_ASAP7_75t_L g125 ( .A(n_68), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_69), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_70), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_71), .B(n_148), .Y(n_458) );
AO32x2_ASAP7_75t_L g180 ( .A1(n_72), .A2(n_155), .A3(n_174), .B1(n_181), .B2(n_186), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_73), .B(n_149), .Y(n_497) );
INVx1_ASAP7_75t_L g170 ( .A(n_74), .Y(n_170) );
INVx1_ASAP7_75t_L g212 ( .A(n_75), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_76), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_77), .B(n_457), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_78), .A2(n_452), .B(n_460), .C(n_550), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g106 ( .A1(n_79), .A2(n_107), .B1(n_727), .B2(n_728), .C1(n_737), .C2(n_741), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_80), .B(n_131), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_81), .Y(n_524) );
INVx1_ASAP7_75t_L g750 ( .A(n_82), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_83), .B(n_456), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_85), .B(n_183), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_86), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_87), .B(n_131), .Y(n_216) );
INVx2_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_89), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_90), .B(n_173), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_91), .B(n_131), .Y(n_159) );
OR2x2_ASAP7_75t_L g434 ( .A(n_93), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g726 ( .A(n_93), .Y(n_726) );
OR2x2_ASAP7_75t_L g754 ( .A(n_93), .B(n_744), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_94), .A2(n_103), .B1(n_131), .B2(n_132), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_95), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g455 ( .A(n_96), .Y(n_455) );
INVxp67_ASAP7_75t_L g527 ( .A(n_97), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_98), .B(n_131), .Y(n_168) );
INVx1_ASAP7_75t_L g493 ( .A(n_99), .Y(n_493) );
INVx1_ASAP7_75t_L g551 ( .A(n_100), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_101), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g518 ( .A(n_102), .B(n_176), .Y(n_518) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_432), .B1(n_438), .B2(n_725), .Y(n_107) );
INVx1_ASAP7_75t_L g738 ( .A(n_108), .Y(n_738) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_109), .A2(n_110), .B1(n_761), .B2(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_SL g110 ( .A(n_111), .B(n_397), .Y(n_110) );
NOR3xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_301), .C(n_385), .Y(n_111) );
NAND4xp25_ASAP7_75t_L g112 ( .A(n_113), .B(n_244), .C(n_266), .D(n_282), .Y(n_112) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_177), .B1(n_203), .B2(n_222), .C(n_230), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_153), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_116), .B(n_222), .Y(n_256) );
NAND4xp25_ASAP7_75t_L g296 ( .A(n_116), .B(n_284), .C(n_297), .D(n_299), .Y(n_296) );
INVxp67_ASAP7_75t_L g413 ( .A(n_116), .Y(n_413) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g295 ( .A(n_117), .B(n_233), .Y(n_295) );
AND2x2_ASAP7_75t_L g319 ( .A(n_117), .B(n_153), .Y(n_319) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g286 ( .A(n_118), .B(n_221), .Y(n_286) );
AND2x2_ASAP7_75t_L g326 ( .A(n_118), .B(n_307), .Y(n_326) );
AND2x2_ASAP7_75t_L g343 ( .A(n_118), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_118), .B(n_154), .Y(n_367) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g220 ( .A(n_119), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g238 ( .A(n_119), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g250 ( .A(n_119), .B(n_154), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_119), .B(n_164), .Y(n_272) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_127), .B(n_152), .Y(n_119) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_120), .A2(n_165), .B(n_175), .Y(n_164) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_121), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_123), .B(n_124), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_141), .B(n_150), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_134), .C(n_137), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_130), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_130), .A2(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g136 ( .A(n_133), .Y(n_136) );
INVx1_ASAP7_75t_L g144 ( .A(n_133), .Y(n_144) );
INVx3_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_135), .Y(n_553) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g183 ( .A(n_136), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
AND2x6_ASAP7_75t_L g452 ( .A(n_136), .B(n_453), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_137), .A2(n_551), .B(n_552), .C(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_138), .A2(n_215), .B(n_216), .Y(n_214) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g457 ( .A(n_139), .Y(n_457) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g149 ( .A(n_140), .Y(n_149) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx1_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
AND2x2_ASAP7_75t_L g448 ( .A(n_140), .B(n_144), .Y(n_448) );
INVx1_ASAP7_75t_L g453 ( .A(n_140), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_146), .C(n_147), .Y(n_141) );
O2A1O1Ixp5_ASAP7_75t_L g169 ( .A1(n_142), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_142), .A2(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_147), .A2(n_161), .B(n_162), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_147), .A2(n_173), .B1(n_201), .B2(n_202), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_147), .A2(n_173), .B1(n_226), .B2(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_148), .A2(n_158), .B(n_159), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_148), .A2(n_167), .B(n_168), .Y(n_166) );
O2A1O1Ixp5_ASAP7_75t_SL g210 ( .A1(n_148), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_148), .B(n_527), .Y(n_526) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_149), .A2(n_173), .B1(n_182), .B2(n_185), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_150), .A2(n_157), .B(n_160), .Y(n_156) );
BUFx3_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_150), .A2(n_190), .B(n_195), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_150), .A2(n_210), .B(n_214), .Y(n_209) );
AND2x4_ASAP7_75t_L g447 ( .A(n_150), .B(n_448), .Y(n_447) );
INVx4_ASAP7_75t_SL g461 ( .A(n_150), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_150), .B(n_448), .Y(n_494) );
AND2x2_ASAP7_75t_L g253 ( .A(n_153), .B(n_254), .Y(n_253) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_153), .A2(n_303), .B1(n_306), .B2(n_308), .C(n_312), .Y(n_302) );
AND2x2_ASAP7_75t_L g361 ( .A(n_153), .B(n_326), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_153), .B(n_343), .Y(n_395) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_164), .Y(n_153) );
INVx3_ASAP7_75t_L g221 ( .A(n_154), .Y(n_221) );
AND2x2_ASAP7_75t_L g270 ( .A(n_154), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g324 ( .A(n_154), .B(n_239), .Y(n_324) );
AND2x2_ASAP7_75t_L g382 ( .A(n_154), .B(n_383), .Y(n_382) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_163), .Y(n_154) );
INVx4_ASAP7_75t_L g224 ( .A(n_155), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_155), .A2(n_503), .B(n_504), .Y(n_502) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_155), .Y(n_521) );
AND2x2_ASAP7_75t_L g222 ( .A(n_164), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g239 ( .A(n_164), .Y(n_239) );
INVx1_ASAP7_75t_L g294 ( .A(n_164), .Y(n_294) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_164), .Y(n_300) );
AND2x2_ASAP7_75t_L g345 ( .A(n_164), .B(n_221), .Y(n_345) );
OR2x2_ASAP7_75t_L g384 ( .A(n_164), .B(n_223), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_174), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_172), .A2(n_196), .B(n_197), .Y(n_195) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g486 ( .A(n_173), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_174), .B(n_224), .C(n_225), .Y(n_243) );
INVx2_ASAP7_75t_L g186 ( .A(n_176), .Y(n_186) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_176), .A2(n_189), .B(n_198), .Y(n_188) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_176), .A2(n_209), .B(n_217), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_176), .A2(n_446), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g476 ( .A(n_176), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_176), .A2(n_513), .B(n_514), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_177), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_187), .Y(n_177) );
AND2x2_ASAP7_75t_L g380 ( .A(n_178), .B(n_377), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_178), .B(n_362), .Y(n_412) );
BUFx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g311 ( .A(n_179), .B(n_235), .Y(n_311) );
AND2x2_ASAP7_75t_L g360 ( .A(n_179), .B(n_206), .Y(n_360) );
INVx1_ASAP7_75t_L g406 ( .A(n_179), .Y(n_406) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
AND2x2_ASAP7_75t_L g261 ( .A(n_180), .B(n_235), .Y(n_261) );
INVx1_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
AND2x2_ASAP7_75t_L g284 ( .A(n_180), .B(n_199), .Y(n_284) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_184), .Y(n_459) );
INVx2_ASAP7_75t_L g487 ( .A(n_184), .Y(n_487) );
INVx1_ASAP7_75t_L g473 ( .A(n_186), .Y(n_473) );
AND2x2_ASAP7_75t_L g352 ( .A(n_187), .B(n_260), .Y(n_352) );
INVx2_ASAP7_75t_L g417 ( .A(n_187), .Y(n_417) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
AND2x2_ASAP7_75t_L g234 ( .A(n_188), .B(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g247 ( .A(n_188), .B(n_207), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_188), .B(n_206), .Y(n_275) );
INVx1_ASAP7_75t_L g281 ( .A(n_188), .Y(n_281) );
INVx1_ASAP7_75t_L g298 ( .A(n_188), .Y(n_298) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_188), .Y(n_310) );
INVx2_ASAP7_75t_L g378 ( .A(n_188), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g235 ( .A(n_199), .Y(n_235) );
BUFx2_ASAP7_75t_L g332 ( .A(n_199), .Y(n_332) );
AND2x2_ASAP7_75t_L g377 ( .A(n_199), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_218), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_205), .B(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_205), .A2(n_376), .B(n_390), .Y(n_400) );
AND2x2_ASAP7_75t_L g425 ( .A(n_205), .B(n_311), .Y(n_425) );
BUFx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g347 ( .A(n_207), .Y(n_347) );
AND2x2_ASAP7_75t_L g376 ( .A(n_207), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_208), .Y(n_260) );
INVx2_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_208), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g233 ( .A(n_219), .Y(n_233) );
OR2x2_ASAP7_75t_L g246 ( .A(n_219), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g314 ( .A(n_219), .B(n_310), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_219), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g415 ( .A(n_219), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_219), .B(n_352), .Y(n_427) );
AND2x2_ASAP7_75t_L g306 ( .A(n_220), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g329 ( .A(n_220), .B(n_222), .Y(n_329) );
INVx2_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
AND2x2_ASAP7_75t_L g269 ( .A(n_221), .B(n_242), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_221), .B(n_294), .Y(n_350) );
AND2x2_ASAP7_75t_L g264 ( .A(n_222), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g411 ( .A(n_222), .Y(n_411) );
AND2x2_ASAP7_75t_L g423 ( .A(n_222), .B(n_286), .Y(n_423) );
AND2x2_ASAP7_75t_L g249 ( .A(n_223), .B(n_239), .Y(n_249) );
INVx1_ASAP7_75t_L g344 ( .A(n_223), .Y(n_344) );
AO21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_228), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_224), .B(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g479 ( .A(n_224), .Y(n_479) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_224), .A2(n_492), .B(n_499), .Y(n_491) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_224), .A2(n_548), .B(n_555), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_224), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g242 ( .A(n_229), .B(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_236), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_233), .B(n_280), .Y(n_289) );
OR2x2_ASAP7_75t_L g421 ( .A(n_233), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g338 ( .A(n_234), .B(n_279), .Y(n_338) );
AND2x2_ASAP7_75t_L g346 ( .A(n_234), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g405 ( .A(n_234), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g429 ( .A(n_234), .B(n_276), .Y(n_429) );
NOR2xp67_ASAP7_75t_L g387 ( .A(n_235), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g416 ( .A(n_235), .B(n_279), .Y(n_416) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
AND2x2_ASAP7_75t_L g268 ( .A(n_238), .B(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g430 ( .A(n_238), .Y(n_430) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g265 ( .A(n_241), .Y(n_265) );
AND2x2_ASAP7_75t_L g316 ( .A(n_241), .B(n_249), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_241), .B(n_384), .Y(n_410) );
INVx2_ASAP7_75t_L g255 ( .A(n_242), .Y(n_255) );
INVx3_ASAP7_75t_L g307 ( .A(n_242), .Y(n_307) );
OR2x2_ASAP7_75t_L g335 ( .A(n_242), .B(n_336), .Y(n_335) );
AOI311xp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_248), .A3(n_250), .B(n_251), .C(n_262), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_245), .A2(n_283), .B(n_285), .C(n_287), .Y(n_282) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_SL g267 ( .A(n_247), .Y(n_267) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g285 ( .A(n_249), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_249), .B(n_265), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_249), .B(n_250), .Y(n_418) );
AND2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_254), .Y(n_340) );
AOI21xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_256), .B(n_257), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g398 ( .A(n_254), .B(n_286), .Y(n_398) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_255), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g292 ( .A(n_255), .Y(n_292) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g283 ( .A(n_259), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
AND2x4_ASAP7_75t_L g390 ( .A(n_261), .B(n_359), .Y(n_390) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_264), .A2(n_330), .B1(n_342), .B2(n_346), .C1(n_348), .C2(n_352), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_270), .C(n_273), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_267), .B(n_311), .Y(n_334) );
INVx1_ASAP7_75t_L g356 ( .A(n_269), .Y(n_356) );
INVx1_ASAP7_75t_L g290 ( .A(n_271), .Y(n_290) );
OR2x2_ASAP7_75t_L g355 ( .A(n_272), .B(n_356), .Y(n_355) );
OAI21xp33_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_276), .B(n_280), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g291 ( .A(n_274), .B(n_292), .C(n_293), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_274), .A2(n_311), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_278), .Y(n_331) );
AND2x2_ASAP7_75t_SL g297 ( .A(n_279), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g388 ( .A(n_279), .Y(n_388) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_279), .Y(n_404) );
INVx2_ASAP7_75t_L g362 ( .A(n_280), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_284), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g336 ( .A(n_286), .Y(n_336) );
OAI221xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B1(n_291), .B2(n_295), .C(n_296), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_290), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g424 ( .A(n_290), .Y(n_424) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g305 ( .A(n_297), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_297), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g363 ( .A(n_297), .B(n_311), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_297), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g396 ( .A(n_297), .B(n_331), .Y(n_396) );
BUFx3_ASAP7_75t_L g359 ( .A(n_298), .Y(n_359) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND5xp2_ASAP7_75t_L g301 ( .A(n_302), .B(n_320), .C(n_341), .D(n_353), .E(n_368), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI32xp33_ASAP7_75t_L g393 ( .A1(n_305), .A2(n_332), .A3(n_348), .B1(n_394), .B2(n_396), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_307), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g317 ( .A(n_311), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B1(n_317), .B2(n_318), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_327), .B1(n_329), .B2(n_330), .C(n_333), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g392 ( .A(n_324), .B(n_343), .Y(n_392) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_329), .A2(n_390), .B1(n_408), .B2(n_413), .C(n_414), .Y(n_407) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx2_ASAP7_75t_L g373 ( .A(n_332), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_337), .B2(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g351 ( .A(n_343), .Y(n_351) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B1(n_361), .B2(n_362), .C1(n_363), .C2(n_364), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_362), .A2(n_409), .B1(n_411), .B2(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_379), .B(n_381), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B(n_391), .C(n_393), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_401), .C(n_426), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_398), .Y(n_402) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_407), .C(n_419), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B(n_418), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22x1_ASAP7_75t_SL g737 ( .A1(n_432), .A2(n_439), .B1(n_738), .B2(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g725 ( .A(n_435), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g744 ( .A(n_435), .Y(n_744) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR3x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_639), .C(n_682), .Y(n_439) );
NAND5xp2_ASAP7_75t_L g440 ( .A(n_441), .B(n_566), .C(n_596), .D(n_613), .E(n_628), .Y(n_440) );
AOI221xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_489), .B1(n_529), .B2(n_535), .C(n_539), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_464), .Y(n_442) );
OR2x2_ASAP7_75t_L g544 ( .A(n_443), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g583 ( .A(n_443), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g601 ( .A(n_443), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_443), .B(n_537), .Y(n_618) );
OR2x2_ASAP7_75t_L g630 ( .A(n_443), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_443), .B(n_589), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_443), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_443), .B(n_567), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_443), .B(n_575), .Y(n_681) );
AND2x2_ASAP7_75t_L g713 ( .A(n_443), .B(n_477), .Y(n_713) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_443), .Y(n_721) );
INVx5_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_444), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g541 ( .A(n_444), .B(n_519), .Y(n_541) );
BUFx2_ASAP7_75t_L g563 ( .A(n_444), .Y(n_563) );
AND2x2_ASAP7_75t_L g592 ( .A(n_444), .B(n_465), .Y(n_592) );
AND2x2_ASAP7_75t_L g647 ( .A(n_444), .B(n_545), .Y(n_647) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_462), .Y(n_444) );
BUFx2_ASAP7_75t_L g468 ( .A(n_447), .Y(n_468) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_451), .A2(n_461), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_451), .A2(n_461), .B(n_524), .C(n_525), .Y(n_523) );
INVx5_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_458), .C(n_459), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_456), .A2(n_459), .B(n_516), .C(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_464), .B(n_601), .Y(n_610) );
OAI32xp33_ASAP7_75t_L g624 ( .A1(n_464), .A2(n_560), .A3(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_464), .B(n_626), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_464), .B(n_544), .Y(n_667) );
INVx1_ASAP7_75t_SL g696 ( .A(n_464), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_464), .B(n_491), .C(n_647), .D(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_477), .Y(n_464) );
INVx5_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
AND2x2_ASAP7_75t_L g567 ( .A(n_465), .B(n_478), .Y(n_567) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_465), .Y(n_646) );
AND2x2_ASAP7_75t_L g716 ( .A(n_465), .B(n_663), .Y(n_716) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_474), .Y(n_465) );
AOI21xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_469), .B(n_473), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x4_ASAP7_75t_L g589 ( .A(n_477), .B(n_538), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_477), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g623 ( .A(n_477), .B(n_545), .Y(n_623) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g537 ( .A(n_478), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g575 ( .A(n_478), .B(n_547), .Y(n_575) );
AND2x2_ASAP7_75t_L g584 ( .A(n_478), .B(n_546), .Y(n_584) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_488), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g652 ( .A1(n_489), .A2(n_653), .B1(n_655), .B2(n_657), .C1(n_660), .C2(n_661), .Y(n_652) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_508), .Y(n_489) );
AND2x2_ASAP7_75t_L g585 ( .A(n_490), .B(n_586), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_490), .B(n_563), .C(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
INVx5_ASAP7_75t_SL g534 ( .A(n_491), .Y(n_534) );
OAI322xp33_ASAP7_75t_L g539 ( .A1(n_491), .A2(n_540), .A3(n_542), .B1(n_543), .B2(n_557), .C1(n_560), .C2(n_562), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_491), .B(n_532), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_491), .B(n_520), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_495), .Y(n_492) );
INVx2_ASAP7_75t_L g532 ( .A(n_501), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_501), .B(n_510), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_508), .B(n_570), .Y(n_625) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g604 ( .A(n_509), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
OR2x2_ASAP7_75t_L g533 ( .A(n_510), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_510), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g572 ( .A(n_510), .B(n_520), .Y(n_572) );
AND2x2_ASAP7_75t_L g595 ( .A(n_510), .B(n_532), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_510), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_510), .B(n_570), .Y(n_611) );
AND2x2_ASAP7_75t_L g619 ( .A(n_510), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_510), .B(n_579), .Y(n_669) );
INVx5_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g559 ( .A(n_511), .B(n_534), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_511), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g586 ( .A(n_511), .B(n_520), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_511), .B(n_633), .Y(n_674) );
OR2x2_ASAP7_75t_L g690 ( .A(n_511), .B(n_634), .Y(n_690) );
AND2x2_ASAP7_75t_SL g697 ( .A(n_511), .B(n_651), .Y(n_697) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_511), .Y(n_704) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
AND2x2_ASAP7_75t_L g558 ( .A(n_519), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g608 ( .A(n_519), .B(n_532), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_519), .B(n_534), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_519), .B(n_570), .Y(n_692) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_520), .B(n_534), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_520), .B(n_532), .Y(n_580) );
OR2x2_ASAP7_75t_L g634 ( .A(n_520), .B(n_532), .Y(n_634) );
AND2x2_ASAP7_75t_L g651 ( .A(n_520), .B(n_531), .Y(n_651) );
INVxp67_ASAP7_75t_L g673 ( .A(n_520), .Y(n_673) );
AND2x2_ASAP7_75t_L g700 ( .A(n_520), .B(n_570), .Y(n_700) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_520), .Y(n_707) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_528), .Y(n_520) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_531), .B(n_581), .Y(n_654) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g570 ( .A(n_532), .B(n_534), .Y(n_570) );
OR2x2_ASAP7_75t_L g637 ( .A(n_532), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g581 ( .A(n_533), .Y(n_581) );
OR2x2_ASAP7_75t_L g642 ( .A(n_533), .B(n_634), .Y(n_642) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g542 ( .A(n_537), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_537), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g543 ( .A(n_538), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_538), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_538), .B(n_545), .Y(n_577) );
INVx2_ASAP7_75t_L g622 ( .A(n_538), .Y(n_622) );
AND2x2_ASAP7_75t_L g635 ( .A(n_538), .B(n_575), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_538), .B(n_584), .Y(n_660) );
INVx1_ASAP7_75t_L g612 ( .A(n_543), .Y(n_612) );
INVx2_ASAP7_75t_SL g599 ( .A(n_544), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_545), .Y(n_602) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_546), .Y(n_565) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g663 ( .A(n_547), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g632 ( .A(n_559), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_559), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_559), .A2(n_641), .B1(n_643), .B2(n_648), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_559), .B(n_651), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_560), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g594 ( .A(n_561), .Y(n_594) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OR2x2_ASAP7_75t_L g576 ( .A(n_563), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_563), .B(n_567), .Y(n_627) );
AND2x2_ASAP7_75t_L g650 ( .A(n_563), .B(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B(n_573), .C(n_587), .Y(n_566) );
INVx1_ASAP7_75t_L g590 ( .A(n_567), .Y(n_590) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_567), .A2(n_699), .B1(n_701), .B2(n_702), .C(n_705), .Y(n_698) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g717 ( .A(n_570), .Y(n_717) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g666 ( .A(n_572), .B(n_605), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_578), .C(n_582), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OAI32xp33_ASAP7_75t_L g691 ( .A1(n_580), .A2(n_581), .A3(n_644), .B1(n_681), .B2(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
AND2x2_ASAP7_75t_L g723 ( .A(n_583), .B(n_622), .Y(n_723) );
AND2x2_ASAP7_75t_L g670 ( .A(n_584), .B(n_622), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_584), .B(n_592), .Y(n_688) );
AOI31xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_590), .A3(n_591), .B(n_593), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_589), .B(n_601), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_589), .B(n_599), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_589), .A2(n_619), .B1(n_709), .B2(n_712), .C(n_714), .Y(n_708) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g614 ( .A(n_594), .B(n_615), .Y(n_614) );
AOI222xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_603), .B1(n_606), .B2(n_609), .C1(n_611), .C2(n_612), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g679 ( .A(n_598), .Y(n_679) );
INVx1_ASAP7_75t_L g701 ( .A(n_601), .Y(n_701) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_604), .A2(n_715), .B1(n_717), .B2(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g620 ( .A(n_605), .Y(n_620) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B1(n_619), .B2(n_621), .C(n_624), .Y(n_613) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g658 ( .A(n_616), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g710 ( .A(n_616), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g685 ( .A(n_621), .Y(n_685) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g649 ( .A(n_622), .Y(n_649) );
INVx1_ASAP7_75t_L g631 ( .A(n_623), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_626), .B(n_713), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_632), .B1(n_635), .B2(n_636), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g722 ( .A(n_635), .Y(n_722) );
INVxp33_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_637), .B(n_681), .Y(n_680) );
OAI32xp33_ASAP7_75t_L g671 ( .A1(n_638), .A2(n_672), .A3(n_673), .B1(n_674), .B2(n_675), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_652), .C(n_664), .D(n_676), .Y(n_639) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
NAND2xp33_ASAP7_75t_SL g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_647), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
CKINVDCx16_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_661), .A2(n_677), .B1(n_694), .B2(n_697), .C(n_698), .Y(n_693) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g712 ( .A(n_663), .B(n_713), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B1(n_668), .B2(n_670), .C(n_671), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_673), .B(n_704), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g682 ( .A(n_683), .B(n_693), .C(n_708), .D(n_719), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B(n_689), .C(n_691), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g724 ( .A(n_711), .Y(n_724) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_724), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g740 ( .A(n_725), .Y(n_740) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_726), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
CKINVDCx14_ASAP7_75t_R g735 ( .A(n_732), .Y(n_735) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
NOR2xp33_ASAP7_75t_SL g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_SL g777 ( .A(n_749), .Y(n_777) );
INVx1_ASAP7_75t_L g776 ( .A(n_751), .Y(n_776) );
OA21x2_ASAP7_75t_L g779 ( .A1(n_751), .A2(n_777), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g768 ( .A(n_752), .Y(n_768) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_754), .Y(n_771) );
BUFx2_ASAP7_75t_L g780 ( .A(n_754), .Y(n_780) );
OAI21xp5_ASAP7_75t_SL g755 ( .A1(n_756), .A2(n_768), .B(n_769), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B1(n_760), .B2(n_767), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_757), .Y(n_767) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_763), .Y(n_766) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
CKINVDCx6p67_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
endmodule