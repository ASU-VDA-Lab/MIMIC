module real_jpeg_1843_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_64),
.B1(n_67),
.B2(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_1),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_81),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_29),
.B1(n_64),
.B2(n_67),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_64),
.B1(n_67),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_5),
.B(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_48),
.C(n_50),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_47),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_64),
.C(n_66),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_5),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_5),
.B(n_84),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_118),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_64),
.B1(n_67),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_12),
.A2(n_58),
.B1(n_64),
.B2(n_67),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_55),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_14),
.A2(n_55),
.B1(n_64),
.B2(n_67),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_122),
.B1(n_201),
.B2(n_202),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_20),
.B(n_97),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_88),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_21),
.B(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_72),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_44),
.C(n_59),
.Y(n_119)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_38),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_32),
.A3(n_34),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_30),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_32),
.B1(n_48),
.B2(n_52),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_31),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_31),
.B(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_38),
.A2(n_113),
.B(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_59),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_57),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_45),
.A2(n_103),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_91),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_50),
.B1(n_65),
.B2(n_66),
.Y(n_70)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_50),
.B(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_56),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_68),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_61),
.A2(n_69),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_68),
.B(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_63),
.A2(n_130),
.B1(n_157),
.B2(n_165),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_64),
.B(n_171),
.Y(n_170)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_129),
.B(n_131),
.Y(n_128)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_118),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_88),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_82),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_82),
.A2(n_83),
.B1(n_149),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_83),
.A2(n_96),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_140),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_86),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_84),
.A2(n_139),
.B(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_95),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_109),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_143),
.B(n_200),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_141),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_141),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_133),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_133),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_195),
.B(n_199),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_185),
.B(n_194),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_167),
.B(n_184),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_160),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_152),
.B1(n_158),
.B2(n_159),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_155),
.C(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_178),
.B(n_183),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_173),
.B(n_177),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_176),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_187),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_198),
.Y(n_199)
);


endmodule