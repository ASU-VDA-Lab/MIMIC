module fake_netlist_5_381_n_169 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_169);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_169;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_154;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_64;
wire n_102;
wire n_106;
wire n_77;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_115;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_97;
wire n_63;
wire n_141;
wire n_166;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_8),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_0),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_3),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_4),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_7),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_7),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_37),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_53),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_52),
.B(n_47),
.C(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_74),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_51),
.A3(n_49),
.B1(n_9),
.B2(n_19),
.C(n_17),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_13),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_27),
.B(n_24),
.C(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_65),
.B(n_67),
.C(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_73),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_68),
.B(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_56),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_56),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

OAI21x1_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_60),
.B(n_66),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_56),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_87),
.B(n_80),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_89),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_72),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_75),
.C(n_78),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_103),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_99),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_77),
.B(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_95),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_112),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2xp67_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_108),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_63),
.C(n_70),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_95),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_108),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_128),
.C(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_126),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_84),
.C(n_55),
.Y(n_139)
);

AND5x1_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_63),
.C(n_97),
.D(n_108),
.E(n_122),
.Y(n_140)
);

NOR3x1_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_125),
.C(n_136),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_122),
.B(n_108),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_132),
.Y(n_143)
);

AND5x1_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_63),
.C(n_105),
.D(n_61),
.E(n_94),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_105),
.B1(n_61),
.B2(n_91),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_105),
.Y(n_155)
);

OA211x2_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_105),
.B(n_101),
.C(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

AND3x4_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_101),
.C(n_150),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_151),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_101),
.Y(n_160)
);

OAI22x1_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_88),
.B1(n_104),
.B2(n_71),
.Y(n_161)
);

NAND5xp2_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_71),
.C(n_82),
.D(n_104),
.E(n_96),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_104),
.B(n_71),
.C(n_82),
.Y(n_163)
);

NOR4xp25_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_159),
.C(n_158),
.D(n_155),
.Y(n_164)
);

AO21x2_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_159),
.B(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_160),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_156),
.B(n_82),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_161),
.B(n_162),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_R g169 ( 
.A1(n_168),
.A2(n_166),
.B1(n_167),
.B2(n_71),
.C(n_82),
.Y(n_169)
);


endmodule