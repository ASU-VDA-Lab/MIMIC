module fake_netlist_5_2182_n_1679 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1679);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1679;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_30),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_50),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_93),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_58),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_25),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_18),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_52),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_108),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_62),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_81),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_61),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_126),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_49),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_32),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_36),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_26),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_51),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_71),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_77),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_29),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_55),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_125),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_29),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_78),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_2),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_53),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_9),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_60),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_149),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_57),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_19),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_25),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_48),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_44),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_107),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_72),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_35),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_23),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_152),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_21),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_101),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_34),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_114),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_113),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_0),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_36),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_6),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_86),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_98),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_146),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_134),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_35),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_132),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_97),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_155),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_127),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_37),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_23),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_119),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_142),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_64),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_73),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_3),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_0),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_49),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_79),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_43),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_143),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_43),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_137),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_68),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_59),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_21),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_96),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_88),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_80),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_24),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_157),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_95),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_42),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_70),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_115),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_37),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_54),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_45),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_32),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_91),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_16),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_39),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_52),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_85),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_47),
.Y(n_305)
);

BUFx2_ASAP7_75t_SL g306 ( 
.A(n_27),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_41),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_33),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_129),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_154),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_65),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_24),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_4),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_22),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_236),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_221),
.B(n_206),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_236),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_192),
.B(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_182),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_199),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_202),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_208),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_200),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_187),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_173),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_210),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_212),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_213),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_187),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_187),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_217),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_187),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_313),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_218),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_223),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_228),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_178),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_195),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_191),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_229),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_290),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_232),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_191),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_238),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_227),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_227),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_231),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_241),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_242),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_247),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_248),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_250),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_255),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_195),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_231),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_235),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_235),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_159),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_256),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_239),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_192),
.B(n_1),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_163),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_239),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_165),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_168),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_180),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_258),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_263),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_198),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_261),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_197),
.B(n_5),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_201),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_262),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_270),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_271),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_220),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_222),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_224),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_275),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_237),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_327),
.B(n_282),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_325),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_328),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_329),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_333),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_345),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_158),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_315),
.A2(n_243),
.B(n_233),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_337),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_378),
.B(n_263),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_349),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_315),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_316),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_351),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_320),
.B(n_158),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_353),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_317),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_317),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_321),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_350),
.B(n_162),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_357),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_322),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_364),
.B(n_197),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_322),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_334),
.B(n_162),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_324),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_324),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_326),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_323),
.B(n_301),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_361),
.Y(n_437)
);

CKINVDCx6p67_ASAP7_75t_R g438 ( 
.A(n_340),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_326),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_362),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_363),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_377),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_348),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_375),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_383),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_348),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_335),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_342),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_343),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_381),
.A2(n_354),
.B(n_352),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_390),
.B(n_205),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_433),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_371),
.B1(n_174),
.B2(n_268),
.Y(n_466)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_390),
.B(n_436),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_433),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_404),
.A2(n_174),
.B1(n_303),
.B2(n_299),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_404),
.A2(n_312),
.B1(n_245),
.B2(n_259),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_406),
.Y(n_476)
);

NOR2x1p5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_160),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_392),
.B(n_422),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_404),
.A2(n_278),
.B1(n_308),
.B2(n_307),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_433),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_442),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_423),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_429),
.B(n_205),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_404),
.A2(n_305),
.B1(n_291),
.B2(n_276),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_418),
.B(n_359),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_401),
.A2(n_369),
.B1(n_384),
.B2(n_360),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_429),
.A2(n_267),
.B(n_352),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

INVx4_ASAP7_75t_SL g496 ( 
.A(n_431),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_429),
.B(n_358),
.Y(n_497)
);

BUFx8_ASAP7_75t_SL g498 ( 
.A(n_393),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_418),
.B(n_385),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_412),
.A2(n_193),
.B1(n_190),
.B2(n_185),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_425),
.B(n_401),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_402),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_425),
.B(n_346),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_347),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_432),
.B(n_205),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

INVxp33_ASAP7_75t_SL g510 ( 
.A(n_456),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_394),
.B(n_205),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_435),
.B(n_379),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_404),
.A2(n_306),
.B1(n_387),
.B2(n_386),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_442),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_402),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_382),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_444),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_445),
.B(n_388),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_439),
.B(n_205),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_395),
.B(n_164),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_439),
.B(n_167),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_172),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_397),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_448),
.B(n_382),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_438),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_417),
.A2(n_280),
.B1(n_294),
.B2(n_302),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_397),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_396),
.B(n_166),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

INVx4_ASAP7_75t_SL g533 ( 
.A(n_391),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_445),
.A2(n_160),
.B1(n_161),
.B2(n_302),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_447),
.A2(n_196),
.B1(n_274),
.B2(n_284),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_460),
.B(n_414),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_398),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_460),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_400),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_460),
.B(n_181),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_430),
.B(n_386),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_447),
.A2(n_387),
.B1(n_388),
.B2(n_257),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_428),
.B(n_203),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_413),
.B(n_354),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_416),
.B(n_166),
.Y(n_547)
);

AND2x6_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_204),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_420),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_391),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_399),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_427),
.B(n_219),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_437),
.B(n_169),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_430),
.B(n_355),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_450),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_399),
.B(n_403),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_403),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_450),
.A2(n_277),
.B1(n_226),
.B2(n_230),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_452),
.B(n_244),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_452),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_455),
.B(n_249),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

AND2x6_ASAP7_75t_L g565 ( 
.A(n_455),
.B(n_264),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_441),
.Y(n_566)
);

AND2x2_ASAP7_75t_SL g567 ( 
.A(n_458),
.B(n_269),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_405),
.B(n_273),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_446),
.B(n_279),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_451),
.A2(n_252),
.B1(n_314),
.B2(n_194),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_459),
.B(n_355),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_458),
.B(n_283),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_459),
.B(n_287),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_407),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_407),
.B(n_293),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_408),
.B(n_311),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_449),
.B(n_163),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_408),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_449),
.B(n_163),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_409),
.B(n_356),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_449),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_409),
.B(n_356),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_453),
.A2(n_373),
.B1(n_370),
.B2(n_367),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_410),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_410),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_411),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_411),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_419),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_419),
.B(n_169),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_453),
.B(n_365),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_453),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_457),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_390),
.B(n_170),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_392),
.B(n_170),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_421),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_429),
.B(n_365),
.Y(n_599)
);

INVx4_ASAP7_75t_SL g600 ( 
.A(n_433),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_436),
.A2(n_373),
.B1(n_370),
.B2(n_367),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_392),
.B(n_171),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_392),
.B(n_171),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_429),
.B(n_366),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_429),
.B(n_366),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_470),
.A2(n_254),
.B(n_266),
.C(n_304),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_543),
.B(n_161),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_480),
.B(n_176),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_470),
.A2(n_596),
.B1(n_491),
.B2(n_499),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_596),
.B(n_240),
.C(n_207),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_605),
.B(n_163),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_176),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_501),
.B(n_177),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_536),
.A2(n_310),
.B(n_309),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_584),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_501),
.B(n_605),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_564),
.B(n_177),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_539),
.B(n_163),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_498),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_491),
.B(n_183),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_537),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_520),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_605),
.B(n_183),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_499),
.B(n_184),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_560),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_605),
.B(n_184),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_554),
.B(n_175),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_539),
.B(n_163),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_605),
.B(n_506),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_599),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_520),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_597),
.B(n_185),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_513),
.B(n_163),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_502),
.B(n_175),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_497),
.B(n_546),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_520),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_561),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_513),
.A2(n_310),
.B1(n_309),
.B2(n_304),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_474),
.A2(n_300),
.B1(n_190),
.B2(n_296),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_193),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_602),
.B(n_272),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_523),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_603),
.B(n_272),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_463),
.B(n_478),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_518),
.Y(n_651)
);

BUFx8_ASAP7_75t_L g652 ( 
.A(n_540),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_466),
.B(n_253),
.C(n_209),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_509),
.B(n_63),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_474),
.A2(n_300),
.B1(n_281),
.B2(n_296),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_466),
.B(n_251),
.C(n_211),
.Y(n_656)
);

NAND2x1_ASAP7_75t_L g657 ( 
.A(n_582),
.B(n_66),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_462),
.A2(n_292),
.B1(n_289),
.B2(n_281),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_547),
.B(n_285),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_479),
.B(n_285),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_547),
.B(n_286),
.Y(n_661)
);

AND2x4_ASAP7_75t_SL g662 ( 
.A(n_594),
.B(n_263),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_483),
.B(n_286),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_523),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_485),
.B(n_289),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_SL g666 ( 
.A1(n_567),
.A2(n_297),
.B1(n_295),
.B2(n_186),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_467),
.B(n_214),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_559),
.B(n_163),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_467),
.B(n_527),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_604),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_553),
.B(n_292),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_486),
.B(n_234),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_488),
.B(n_246),
.Y(n_673)
);

OAI22x1_ASAP7_75t_L g674 ( 
.A1(n_515),
.A2(n_297),
.B1(n_295),
.B2(n_288),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_564),
.B(n_83),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_525),
.B(n_216),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_489),
.B(n_225),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_493),
.B(n_215),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_541),
.B(n_260),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_527),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_507),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_553),
.B(n_265),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_495),
.B(n_288),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_559),
.B(n_284),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_509),
.B(n_576),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_576),
.B(n_274),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_604),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_580),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_505),
.B(n_189),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_569),
.B(n_549),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_598),
.B(n_189),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_587),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_530),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_582),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_566),
.B(n_122),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_572),
.B(n_188),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_469),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_522),
.B(n_188),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_583),
.B(n_186),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_SL g700 ( 
.A(n_566),
.B(n_179),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_469),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_481),
.B(n_179),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_586),
.B(n_156),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_586),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_472),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_508),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_522),
.B(n_552),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_588),
.B(n_150),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_5),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_462),
.B(n_148),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_476),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_481),
.B(n_490),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_490),
.B(n_144),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_593),
.B(n_139),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_473),
.B(n_138),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_593),
.B(n_133),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_550),
.B(n_121),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_476),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_500),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_571),
.B(n_7),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_557),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_473),
.B(n_103),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_550),
.B(n_100),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_484),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_558),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_504),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_568),
.B(n_92),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_550),
.B(n_89),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_550),
.B(n_87),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_558),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_582),
.Y(n_733)
);

INVx8_ASAP7_75t_L g734 ( 
.A(n_574),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_487),
.A2(n_84),
.B1(n_76),
.B2(n_75),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_589),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_492),
.B(n_12),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_503),
.B(n_67),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_526),
.B(n_13),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_487),
.B(n_53),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_556),
.B(n_48),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_494),
.B(n_14),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_567),
.B(n_16),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_571),
.B(n_17),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_559),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_568),
.B(n_22),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_594),
.B(n_26),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_512),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_511),
.B(n_28),
.Y(n_750)
);

BUFx8_ASAP7_75t_L g751 ( 
.A(n_510),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_582),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_511),
.B(n_31),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_496),
.B(n_33),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_713),
.A2(n_468),
.B(n_465),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_609),
.A2(n_516),
.B(n_544),
.C(n_601),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_620),
.A2(n_538),
.B(n_532),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_SL g758 ( 
.A(n_751),
.B(n_528),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_634),
.A2(n_508),
.B1(n_569),
.B2(n_528),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_620),
.A2(n_542),
.B(n_475),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_SL g761 ( 
.A1(n_715),
.A2(n_581),
.B(n_579),
.C(n_534),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_749),
.B(n_516),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_749),
.A2(n_569),
.B1(n_591),
.B2(n_574),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_710),
.A2(n_544),
.B(n_601),
.C(n_524),
.Y(n_764)
);

O2A1O1Ixp5_ASAP7_75t_SL g765 ( 
.A1(n_743),
.A2(n_575),
.B(n_579),
.C(n_581),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_614),
.B(n_475),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_614),
.B(n_482),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_681),
.B(n_482),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_633),
.A2(n_545),
.B(n_521),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_618),
.A2(n_464),
.B(n_461),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_708),
.A2(n_574),
.B1(n_577),
.B2(n_570),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_633),
.A2(n_471),
.B(n_521),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_614),
.A2(n_595),
.B(n_471),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_681),
.B(n_563),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_614),
.A2(n_595),
.B(n_517),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_640),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_680),
.B(n_531),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_669),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_621),
.A2(n_595),
.B(n_517),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_625),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_708),
.A2(n_628),
.B1(n_623),
.B2(n_707),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_621),
.A2(n_595),
.B(n_514),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_623),
.A2(n_628),
.B1(n_685),
.B2(n_680),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_637),
.B(n_565),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_635),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_710),
.A2(n_575),
.B(n_578),
.C(n_585),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_637),
.B(n_565),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_676),
.A2(n_582),
.B(n_563),
.Y(n_788)
);

NAND2x1_ASAP7_75t_L g789 ( 
.A(n_752),
.B(n_559),
.Y(n_789)
);

NOR2x1_ASAP7_75t_R g790 ( 
.A(n_622),
.B(n_477),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_635),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_667),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_676),
.A2(n_565),
.B(n_563),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_722),
.A2(n_585),
.B(n_534),
.C(n_529),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_743),
.A2(n_535),
.B(n_529),
.C(n_563),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_721),
.B(n_38),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_646),
.B(n_649),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_646),
.B(n_565),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_685),
.A2(n_565),
.B1(n_496),
.B2(n_533),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_659),
.A2(n_671),
.B1(n_661),
.B2(n_613),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_694),
.B(n_600),
.Y(n_802)
);

O2A1O1Ixp5_ASAP7_75t_L g803 ( 
.A1(n_679),
.A2(n_533),
.B(n_548),
.C(n_519),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_649),
.B(n_600),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_645),
.B(n_533),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_638),
.A2(n_548),
.B(n_519),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_717),
.A2(n_548),
.B(n_519),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_638),
.A2(n_615),
.B(n_717),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_659),
.B(n_661),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_751),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_724),
.A2(n_548),
.B(n_519),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_724),
.A2(n_41),
.B(n_44),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_46),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_715),
.A2(n_46),
.B(n_47),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_752),
.A2(n_650),
.B(n_611),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_716),
.A2(n_718),
.B(n_627),
.Y(n_816)
);

OR2x4_ASAP7_75t_L g817 ( 
.A(n_696),
.B(n_737),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_682),
.B(n_608),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_711),
.A2(n_705),
.B(n_631),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_714),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_746),
.A2(n_727),
.B1(n_732),
.B2(n_722),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_670),
.B(n_687),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_745),
.A2(n_725),
.B(n_719),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_723),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_682),
.B(n_629),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_624),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_612),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_698),
.B(n_632),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_630),
.B(n_642),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_639),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_698),
.A2(n_750),
.B(n_753),
.C(n_651),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_730),
.A2(n_703),
.B(n_709),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_648),
.B(n_688),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_617),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_624),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_692),
.B(n_704),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_738),
.A2(n_647),
.B(n_693),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_616),
.B(n_741),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_607),
.Y(n_839)
);

INVx8_ASAP7_75t_L g840 ( 
.A(n_690),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_699),
.B(n_641),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_744),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_697),
.A2(n_712),
.B(n_728),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_SL g844 ( 
.A1(n_742),
.A2(n_739),
.B(n_702),
.C(n_754),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_694),
.B(n_733),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_612),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_736),
.B(n_740),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_694),
.B(n_733),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_672),
.B(n_678),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_739),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_664),
.Y(n_851)
);

AO21x2_ASAP7_75t_L g852 ( 
.A1(n_731),
.A2(n_668),
.B(n_686),
.Y(n_852)
);

AND2x2_ASAP7_75t_SL g853 ( 
.A(n_746),
.B(n_732),
.Y(n_853)
);

OA22x2_ASAP7_75t_L g854 ( 
.A1(n_666),
.A2(n_674),
.B1(n_742),
.B2(n_691),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_662),
.B(n_700),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_701),
.A2(n_726),
.B(n_706),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_727),
.A2(n_654),
.B1(n_754),
.B2(n_656),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_652),
.Y(n_858)
);

AO21x1_ASAP7_75t_L g859 ( 
.A1(n_654),
.A2(n_731),
.B(n_606),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_653),
.A2(n_735),
.B1(n_733),
.B2(n_694),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_720),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_610),
.A2(n_677),
.B(n_673),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_652),
.Y(n_863)
);

CKINVDCx6p67_ASAP7_75t_R g864 ( 
.A(n_626),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_660),
.A2(n_665),
.B(n_663),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_686),
.B(n_691),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_683),
.B(n_689),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_619),
.B(n_658),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_733),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_643),
.B(n_747),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_690),
.Y(n_871)
);

OAI321xp33_ASAP7_75t_L g872 ( 
.A1(n_644),
.A2(n_655),
.A3(n_729),
.B1(n_690),
.B2(n_748),
.C(n_684),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_675),
.B(n_695),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_657),
.A2(n_729),
.B(n_734),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_734),
.A2(n_536),
.B(n_713),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_734),
.A2(n_536),
.B(n_713),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_640),
.Y(n_877)
);

AOI22x1_ASAP7_75t_L g878 ( 
.A1(n_749),
.A2(n_707),
.B1(n_705),
.B2(n_654),
.Y(n_878)
);

AND2x6_ASAP7_75t_L g879 ( 
.A(n_614),
.B(n_509),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_609),
.A2(n_470),
.B(n_390),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_749),
.B(n_470),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_749),
.B(n_470),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_635),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_635),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_669),
.B(n_497),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_667),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_609),
.A2(n_634),
.B1(n_470),
.B2(n_749),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_609),
.A2(n_634),
.B1(n_470),
.B2(n_749),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_635),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_749),
.B(n_470),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_743),
.A2(n_470),
.B(n_680),
.C(n_462),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_749),
.B(n_470),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_895)
);

OA22x2_ASAP7_75t_L g896 ( 
.A1(n_609),
.A2(n_743),
.B1(n_680),
.B2(n_666),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_609),
.A2(n_470),
.B(n_722),
.C(n_710),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_614),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_609),
.B(n_470),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_614),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_609),
.A2(n_470),
.B1(n_708),
.B2(n_628),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_751),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_669),
.B(n_497),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_620),
.A2(n_633),
.B(n_536),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_635),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_749),
.B(n_470),
.Y(n_906)
);

NOR2xp67_ASAP7_75t_L g907 ( 
.A(n_610),
.B(n_564),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_635),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_749),
.B(n_470),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_SL g910 ( 
.A(n_751),
.B(n_510),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_609),
.A2(n_470),
.B(n_722),
.C(n_710),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_609),
.B(n_470),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_914)
);

AOI33xp33_ASAP7_75t_L g915 ( 
.A1(n_727),
.A2(n_529),
.A3(n_466),
.B1(n_534),
.B2(n_732),
.B3(n_502),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_749),
.B(n_470),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_609),
.A2(n_470),
.B1(n_708),
.B2(n_628),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_614),
.B(n_621),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_749),
.B(n_470),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_614),
.B(n_621),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_635),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_620),
.A2(n_633),
.B(n_536),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_713),
.A2(n_536),
.B(n_634),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_821),
.A2(n_853),
.B(n_913),
.C(n_899),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_815),
.A2(n_816),
.B(n_832),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_837),
.A2(n_887),
.B(n_882),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_886),
.B(n_903),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_895),
.A2(n_914),
.B(n_911),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_809),
.A2(n_800),
.B(n_797),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_821),
.A2(n_853),
.B(n_913),
.C(n_899),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_778),
.Y(n_933)
);

AOI21xp33_ASAP7_75t_L g934 ( 
.A1(n_880),
.A2(n_818),
.B(n_828),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_783),
.A2(n_781),
.B(n_818),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_901),
.B(n_917),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_881),
.B(n_883),
.Y(n_937)
);

AO21x1_ASAP7_75t_L g938 ( 
.A1(n_813),
.A2(n_890),
.B(n_889),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_765),
.A2(n_876),
.B(n_875),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_919),
.A2(n_924),
.B(n_904),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_828),
.A2(n_897),
.B1(n_912),
.B2(n_866),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_892),
.B(n_894),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_906),
.B(n_909),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_776),
.B(n_842),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_916),
.B(n_920),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_825),
.B(n_762),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_808),
.A2(n_769),
.B(n_755),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_840),
.B(n_858),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_897),
.A2(n_912),
.B(n_893),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_777),
.B(n_867),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_804),
.A2(n_787),
.B(n_784),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_842),
.B(n_839),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_877),
.B(n_830),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_878),
.A2(n_819),
.B(n_770),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_849),
.B(n_777),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_838),
.B(n_866),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_888),
.B(n_796),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_857),
.A2(n_870),
.B1(n_831),
.B2(n_850),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_798),
.A2(n_873),
.B(n_805),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_796),
.B(n_792),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_873),
.A2(n_918),
.B(n_921),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_824),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_855),
.B(n_846),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_859),
.A2(n_786),
.A3(n_764),
.B(n_756),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_898),
.B(n_900),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_829),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_850),
.B(n_756),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_SL g968 ( 
.A(n_915),
.B(n_795),
.C(n_794),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_785),
.B(n_833),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_817),
.B(n_896),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_918),
.A2(n_921),
.B(n_848),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_785),
.B(n_836),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_760),
.A2(n_772),
.B(n_757),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_885),
.B(n_891),
.Y(n_974)
);

AO31x2_ASAP7_75t_L g975 ( 
.A1(n_764),
.A2(n_771),
.A3(n_794),
.B(n_759),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_865),
.A2(n_788),
.B(n_793),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_SL g977 ( 
.A1(n_857),
.A2(n_814),
.B1(n_763),
.B2(n_812),
.C(n_768),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_789),
.A2(n_845),
.B(n_898),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_846),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_845),
.A2(n_766),
.B(n_767),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_862),
.B(n_834),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_774),
.A2(n_761),
.B(n_803),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_761),
.A2(n_844),
.B(n_847),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_872),
.A2(n_834),
.B(n_868),
.C(n_907),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_841),
.B(n_827),
.C(n_908),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_869),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_791),
.A2(n_922),
.B(n_905),
.C(n_884),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_SL g988 ( 
.A1(n_799),
.A2(n_852),
.B(n_874),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_900),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_766),
.A2(n_767),
.B(n_844),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_860),
.A2(n_773),
.B(n_775),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_896),
.B(n_820),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_807),
.A2(n_811),
.B(n_806),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_817),
.A2(n_854),
.B1(n_822),
.B2(n_879),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_869),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_822),
.B(n_801),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_779),
.A2(n_782),
.B(n_856),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_780),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_871),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_871),
.Y(n_1000)
);

AOI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_854),
.A2(n_851),
.B(n_861),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_802),
.A2(n_879),
.B(n_840),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_879),
.A2(n_840),
.B(n_758),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_864),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_879),
.B(n_910),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_879),
.A2(n_790),
.B(n_863),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_810),
.A2(n_902),
.B(n_826),
.Y(n_1007)
);

INVx5_ASAP7_75t_L g1008 ( 
.A(n_835),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_810),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_815),
.A2(n_621),
.B(n_614),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_882),
.A2(n_924),
.B(n_919),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_886),
.B(n_669),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_815),
.A2(n_621),
.B(n_614),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_815),
.A2(n_621),
.B(n_614),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_780),
.Y(n_1015)
);

OAI22x1_ASAP7_75t_L g1016 ( 
.A1(n_899),
.A2(n_609),
.B1(n_913),
.B2(n_901),
.Y(n_1016)
);

AO31x2_ASAP7_75t_L g1017 ( 
.A1(n_897),
.A2(n_912),
.A3(n_859),
.B(n_831),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_899),
.A2(n_609),
.B1(n_913),
.B2(n_809),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_776),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_843),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_778),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_840),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_818),
.B(n_809),
.Y(n_1025)
);

BUFx8_ASAP7_75t_L g1026 ( 
.A(n_858),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_818),
.B(n_809),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_815),
.A2(n_621),
.B(n_614),
.Y(n_1028)
);

INVx8_ASAP7_75t_L g1029 ( 
.A(n_840),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_809),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_818),
.B(n_809),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_810),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_882),
.A2(n_924),
.B(n_919),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_808),
.A2(n_819),
.B(n_897),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_886),
.B(n_669),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_899),
.B(n_609),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_840),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_SL g1041 ( 
.A1(n_899),
.A2(n_609),
.B(n_470),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_818),
.B(n_809),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_809),
.A2(n_800),
.B(n_797),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_809),
.A2(n_800),
.B(n_797),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_778),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_897),
.A2(n_912),
.A3(n_859),
.B(n_831),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_843),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_886),
.B(n_669),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_843),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_815),
.A2(n_621),
.B(n_614),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_776),
.Y(n_1052)
);

AND2x2_ASAP7_75t_SL g1053 ( 
.A(n_853),
.B(n_821),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_818),
.B(n_809),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_818),
.B(n_809),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_821),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_843),
.A2(n_823),
.B(n_923),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_886),
.B(n_669),
.Y(n_1060)
);

AO221x2_ASAP7_75t_L g1061 ( 
.A1(n_800),
.A2(n_666),
.B1(n_781),
.B2(n_809),
.C(n_890),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_877),
.B(n_651),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_962),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_1003),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_926),
.A2(n_976),
.B(n_940),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_988),
.A2(n_1013),
.B(n_1010),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_998),
.Y(n_1067)
);

INVxp33_ASAP7_75t_L g1068 ( 
.A(n_1020),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_1029),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_963),
.Y(n_1071)
);

AO32x2_ASAP7_75t_L g1072 ( 
.A1(n_958),
.A2(n_964),
.A3(n_1017),
.B1(n_1047),
.B2(n_949),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_1009),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_999),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1041),
.B(n_1038),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1038),
.B(n_1019),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1014),
.A2(n_1051),
.B(n_1028),
.Y(n_1078)
);

OAI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_1042),
.A2(n_1056),
.B(n_1054),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_950),
.B(n_955),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_950),
.B(n_946),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_937),
.B(n_942),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_927),
.A2(n_1055),
.B(n_1057),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1061),
.A2(n_1053),
.B1(n_1016),
.B2(n_968),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_929),
.B(n_1012),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_943),
.B(n_945),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_933),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_985),
.B(n_1015),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_925),
.B(n_932),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1037),
.B(n_1049),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_996),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1024),
.B(n_1040),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_956),
.B(n_1060),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_969),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_1023),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_931),
.A2(n_1045),
.B(n_1043),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_936),
.B(n_934),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_1009),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1029),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1046),
.B(n_957),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_925),
.B(n_932),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_960),
.B(n_944),
.Y(n_1102)
);

CKINVDCx8_ASAP7_75t_R g1103 ( 
.A(n_1008),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1053),
.B(n_1058),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_1029),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_952),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1058),
.B(n_941),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_972),
.Y(n_1109)
);

CKINVDCx11_ASAP7_75t_R g1110 ( 
.A(n_948),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1003),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_953),
.B(n_1020),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_939),
.A2(n_981),
.B(n_991),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_967),
.B(n_1061),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_948),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_970),
.B(n_1052),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_984),
.A2(n_970),
.B(n_1001),
.C(n_992),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1052),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1036),
.A2(n_984),
.B(n_982),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1061),
.B(n_935),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_994),
.A2(n_977),
.B(n_961),
.C(n_990),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1005),
.A2(n_1062),
.B1(n_971),
.B2(n_1002),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_986),
.B(n_995),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_948),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_979),
.B(n_1062),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_1062),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_SL g1127 ( 
.A(n_1026),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_986),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_938),
.A2(n_993),
.B(n_947),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_R g1130 ( 
.A(n_1033),
.B(n_1004),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_954),
.A2(n_928),
.B(n_978),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_975),
.B(n_1017),
.Y(n_1132)
);

INVx2_ASAP7_75t_R g1133 ( 
.A(n_1008),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1006),
.B(n_974),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_974),
.B(n_989),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_974),
.B(n_1017),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_L g1137 ( 
.A(n_1008),
.B(n_1033),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_995),
.B1(n_980),
.B2(n_1008),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_993),
.A2(n_973),
.B(n_959),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_927),
.A2(n_1039),
.B(n_1034),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_975),
.B(n_1047),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1017),
.B(n_1047),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_987),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1026),
.A2(n_1007),
.B1(n_975),
.B2(n_965),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1018),
.A2(n_1034),
.B(n_1059),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1026),
.Y(n_1146)
);

AO21x1_ASAP7_75t_L g1147 ( 
.A1(n_951),
.A2(n_930),
.B(n_1035),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_987),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_SL g1149 ( 
.A(n_1021),
.B(n_1050),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_975),
.B(n_1047),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_964),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_964),
.B(n_1011),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_997),
.Y(n_1153)
);

AO21x1_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_1048),
.B(n_1050),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_1018),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1022),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_1031),
.B(n_1044),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1044),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_1055),
.B(n_1057),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_929),
.B(n_1012),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_926),
.A2(n_976),
.B(n_816),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_934),
.A2(n_470),
.B(n_912),
.C(n_897),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1164)
);

OAI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_1038),
.A2(n_470),
.B(n_609),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1038),
.A2(n_917),
.B(n_901),
.C(n_913),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_963),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_934),
.A2(n_470),
.B(n_912),
.C(n_897),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_L g1169 ( 
.A(n_925),
.B(n_821),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_999),
.Y(n_1171)
);

O2A1O1Ixp5_ASAP7_75t_L g1172 ( 
.A1(n_931),
.A2(n_809),
.B(n_797),
.C(n_800),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_962),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_926),
.A2(n_976),
.B(n_816),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1019),
.A2(n_821),
.B1(n_853),
.B2(n_901),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_998),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_929),
.B(n_1012),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_933),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_962),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_999),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_SL g1183 ( 
.A(n_966),
.B(n_873),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_962),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1038),
.A2(n_917),
.B(n_901),
.C(n_913),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_963),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1003),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1020),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1024),
.B(n_1040),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1024),
.B(n_1040),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_933),
.Y(n_1193)
);

INVx3_ASAP7_75t_SL g1194 ( 
.A(n_1009),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_929),
.B(n_1012),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_963),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_R g1198 ( 
.A(n_1009),
.B(n_393),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1077),
.A2(n_1080),
.B1(n_1166),
.B2(n_1187),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1136),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1063),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1096),
.A2(n_1175),
.B(n_1161),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1118),
.Y(n_1203)
);

BUFx8_ASAP7_75t_L g1204 ( 
.A(n_1071),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_1106),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1082),
.A2(n_1086),
.B1(n_1081),
.B2(n_1165),
.Y(n_1206)
);

AO21x1_ASAP7_75t_L g1207 ( 
.A1(n_1162),
.A2(n_1168),
.B(n_1176),
.Y(n_1207)
);

BUFx8_ASAP7_75t_L g1208 ( 
.A(n_1167),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1176),
.A2(n_1169),
.B1(n_1089),
.B2(n_1076),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1090),
.A2(n_1097),
.B1(n_1179),
.B2(n_1160),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1174),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1181),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1101),
.A2(n_1120),
.B1(n_1114),
.B2(n_1081),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1083),
.A2(n_1145),
.B(n_1140),
.Y(n_1214)
);

BUFx8_ASAP7_75t_L g1215 ( 
.A(n_1188),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1084),
.A2(n_1101),
.B1(n_1114),
.B2(n_1108),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1108),
.A2(n_1079),
.B1(n_1196),
.B2(n_1085),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1185),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1106),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1103),
.Y(n_1220)
);

BUFx2_ASAP7_75t_R g1221 ( 
.A(n_1073),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1098),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1100),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1087),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1087),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1197),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1117),
.B(n_1141),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1194),
.Y(n_1228)
);

OAI21xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1082),
.A2(n_1086),
.B(n_1184),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1112),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1104),
.B(n_1135),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1163),
.A2(n_1186),
.B1(n_1164),
.B2(n_1184),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1070),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1104),
.B(n_1069),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1126),
.A2(n_1093),
.B1(n_1116),
.B2(n_1144),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1126),
.A2(n_1102),
.B1(n_1134),
.B2(n_1195),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1105),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1094),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1134),
.A2(n_1074),
.B1(n_1195),
.B2(n_1178),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1146),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1069),
.A2(n_1178),
.B1(n_1170),
.B2(n_1173),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1074),
.A2(n_1170),
.B1(n_1173),
.B2(n_1068),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1091),
.A2(n_1125),
.B1(n_1122),
.B2(n_1107),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1109),
.B(n_1107),
.Y(n_1244)
);

AO22x1_ASAP7_75t_L g1245 ( 
.A1(n_1124),
.A2(n_1148),
.B1(n_1143),
.B2(n_1115),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1111),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1088),
.A2(n_1137),
.B1(n_1124),
.B2(n_1180),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1131),
.A2(n_1066),
.B(n_1078),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1095),
.A2(n_1180),
.B1(n_1193),
.B2(n_1122),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1095),
.A2(n_1193),
.B1(n_1127),
.B2(n_1171),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1172),
.A2(n_1113),
.B(n_1121),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1189),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1151),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1119),
.A2(n_1065),
.B(n_1139),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1152),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1139),
.A2(n_1129),
.B(n_1147),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1190),
.B(n_1067),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1092),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1189),
.B(n_1153),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1075),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1198),
.A2(n_1183),
.B1(n_1130),
.B2(n_1182),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1138),
.A2(n_1177),
.B(n_1129),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1191),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1110),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1150),
.A2(n_1132),
.B1(n_1133),
.B2(n_1142),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1128),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1132),
.A2(n_1192),
.B1(n_1191),
.B2(n_1099),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1192),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1072),
.B(n_1123),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1154),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1072),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1149),
.A2(n_1099),
.B1(n_1158),
.B2(n_1156),
.Y(n_1272)
);

AOI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1157),
.A2(n_1159),
.B(n_1149),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1155),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_1159),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1157),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1087),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1106),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1064),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1165),
.A2(n_1061),
.B1(n_899),
.B2(n_913),
.Y(n_1280)
);

NOR2x1_ASAP7_75t_R g1281 ( 
.A(n_1073),
.B(n_622),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1098),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1080),
.B(n_1077),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1172),
.A2(n_609),
.B(n_809),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_SL g1285 ( 
.A1(n_1183),
.A2(n_935),
.B(n_983),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1077),
.A2(n_853),
.B1(n_470),
.B2(n_1038),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1106),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1106),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1165),
.A2(n_1061),
.B1(n_899),
.B2(n_913),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1087),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1106),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1063),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1198),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1080),
.B(n_1077),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1106),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1106),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1063),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_1194),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1203),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1202),
.A2(n_1251),
.B(n_1270),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1204),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1283),
.B(n_1294),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1273),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1203),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1232),
.B(n_1242),
.Y(n_1305)
);

BUFx2_ASAP7_75t_R g1306 ( 
.A(n_1293),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1200),
.B(n_1269),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1231),
.B(n_1227),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1225),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1226),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1231),
.B(n_1227),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1200),
.B(n_1269),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1253),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1274),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1234),
.B(n_1255),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1255),
.B(n_1275),
.Y(n_1316)
);

INVxp33_ASAP7_75t_L g1317 ( 
.A(n_1260),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1234),
.B(n_1209),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1273),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1204),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_1244),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1259),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1259),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1241),
.B(n_1286),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1259),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1276),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1204),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1208),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1240),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1271),
.B(n_1213),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1199),
.B(n_1216),
.Y(n_1331)
);

NAND4xp25_ASAP7_75t_L g1332 ( 
.A(n_1249),
.B(n_1289),
.C(n_1280),
.D(n_1217),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1201),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1223),
.B(n_1230),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1211),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1212),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1285),
.A2(n_1248),
.B(n_1207),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1214),
.A2(n_1284),
.B(n_1207),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1226),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1218),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1265),
.B(n_1210),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1277),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1248),
.A2(n_1262),
.B(n_1206),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1243),
.A2(n_1239),
.B(n_1236),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1290),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1245),
.B(n_1254),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1237),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1235),
.A2(n_1292),
.B(n_1297),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1229),
.B(n_1238),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1223),
.B(n_1224),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1208),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1208),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1246),
.A2(n_1252),
.B(n_1279),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1237),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1215),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1215),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1330),
.B(n_1338),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1330),
.B(n_1256),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1303),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1313),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1350),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1331),
.A2(n_1250),
.B1(n_1257),
.B2(n_1261),
.C(n_1245),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1321),
.B(n_1272),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1315),
.B(n_1314),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1337),
.B(n_1300),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1315),
.B(n_1247),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1346),
.A2(n_1266),
.B(n_1267),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1337),
.B(n_1300),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1346),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1305),
.B(n_1223),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1300),
.B(n_1307),
.Y(n_1373)
);

CKINVDCx6p67_ASAP7_75t_R g1374 ( 
.A(n_1301),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1316),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1346),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1307),
.B(n_1268),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1346),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1316),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1314),
.B(n_1215),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1349),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1349),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1312),
.B(n_1263),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1346),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1312),
.B(n_1258),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1354),
.Y(n_1386)
);

NOR2x1_ASAP7_75t_SL g1387 ( 
.A(n_1303),
.B(n_1205),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1355),
.B(n_1205),
.Y(n_1388)
);

OAI222xp33_ASAP7_75t_L g1389 ( 
.A1(n_1331),
.A2(n_1264),
.B1(n_1291),
.B2(n_1293),
.C1(n_1222),
.C2(n_1282),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1364),
.A2(n_1324),
.B1(n_1302),
.B2(n_1334),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1360),
.B(n_1326),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1360),
.B(n_1308),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1364),
.B(n_1332),
.C(n_1341),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1363),
.B(n_1304),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1363),
.B(n_1342),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1372),
.B(n_1341),
.C(n_1351),
.Y(n_1396)
);

AOI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1372),
.A2(n_1309),
.B1(n_1345),
.B2(n_1347),
.C(n_1356),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1365),
.A2(n_1358),
.B1(n_1328),
.B2(n_1352),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1375),
.B(n_1310),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1365),
.A2(n_1318),
.B1(n_1220),
.B2(n_1339),
.C(n_1308),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1375),
.B(n_1311),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1380),
.B(n_1299),
.C(n_1348),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1379),
.B(n_1311),
.Y(n_1403)
);

NOR3xp33_ASAP7_75t_L g1404 ( 
.A(n_1389),
.B(n_1291),
.C(n_1352),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1389),
.A2(n_1317),
.B(n_1318),
.Y(n_1405)
);

NAND2x1_ASAP7_75t_L g1406 ( 
.A(n_1388),
.B(n_1303),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1380),
.A2(n_1328),
.B1(n_1358),
.B2(n_1301),
.Y(n_1407)
);

AOI21xp33_ASAP7_75t_L g1408 ( 
.A1(n_1368),
.A2(n_1379),
.B(n_1348),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1359),
.B(n_1319),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1377),
.B(n_1299),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1367),
.B(n_1370),
.C(n_1368),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1359),
.B(n_1319),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1369),
.A2(n_1219),
.B(n_1295),
.Y(n_1413)
);

NOR3xp33_ASAP7_75t_L g1414 ( 
.A(n_1369),
.B(n_1233),
.C(n_1323),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1373),
.B(n_1319),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1377),
.B(n_1333),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1377),
.B(n_1333),
.Y(n_1417)
);

OAI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1371),
.A2(n_1220),
.B1(n_1288),
.B2(n_1287),
.C(n_1296),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1373),
.B(n_1319),
.Y(n_1420)
);

OAI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1371),
.A2(n_1288),
.B1(n_1287),
.B2(n_1296),
.C(n_1301),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1373),
.B(n_1371),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1367),
.B(n_1370),
.C(n_1348),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1383),
.A2(n_1344),
.B1(n_1329),
.B2(n_1353),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1388),
.B(n_1320),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1378),
.A2(n_1219),
.B(n_1278),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1387),
.A2(n_1344),
.B1(n_1343),
.B2(n_1327),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1384),
.B(n_1322),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1384),
.B(n_1322),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1383),
.B(n_1336),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1385),
.B(n_1340),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1385),
.B(n_1340),
.Y(n_1433)
);

NOR3xp33_ASAP7_75t_SL g1434 ( 
.A(n_1362),
.B(n_1323),
.C(n_1325),
.Y(n_1434)
);

AND4x1_ASAP7_75t_L g1435 ( 
.A(n_1374),
.B(n_1325),
.C(n_1306),
.D(n_1221),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1411),
.B(n_1381),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1415),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1393),
.A2(n_1370),
.B(n_1367),
.Y(n_1438)
);

NAND3x1_ASAP7_75t_SL g1439 ( 
.A(n_1405),
.B(n_1374),
.C(n_1387),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1422),
.B(n_1376),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1409),
.B(n_1376),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1406),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1411),
.B(n_1381),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1406),
.B(n_1376),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1420),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1423),
.B(n_1382),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1429),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1412),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1429),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1391),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1416),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1423),
.B(n_1382),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1392),
.B(n_1376),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1402),
.B(n_1382),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1430),
.B(n_1376),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1417),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1392),
.B(n_1376),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1391),
.B(n_1386),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1431),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1427),
.B(n_1386),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1402),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1425),
.B(n_1386),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1419),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1428),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1395),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1447),
.B(n_1414),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1436),
.B(n_1394),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1450),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1449),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1450),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1450),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1447),
.B(n_1426),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1444),
.B(n_1388),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1450),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1465),
.B(n_1329),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1447),
.B(n_1426),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1447),
.B(n_1401),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1465),
.B(n_1396),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1458),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1445),
.Y(n_1480)
);

NOR3xp33_ASAP7_75t_L g1481 ( 
.A(n_1438),
.B(n_1393),
.C(n_1396),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1436),
.B(n_1399),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1448),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1447),
.B(n_1403),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1463),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1447),
.B(n_1410),
.Y(n_1486)
);

INVx3_ASAP7_75t_SL g1487 ( 
.A(n_1444),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1443),
.B(n_1432),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1463),
.B(n_1397),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1438),
.A2(n_1413),
.B(n_1404),
.C(n_1400),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1464),
.B(n_1433),
.Y(n_1492)
);

CKINVDCx14_ASAP7_75t_R g1493 ( 
.A(n_1457),
.Y(n_1493)
);

NAND2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1442),
.B(n_1361),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1462),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1385),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1437),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1453),
.B(n_1388),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1444),
.B(n_1388),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1448),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1437),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1497),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1503)
);

NOR2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1478),
.B(n_1320),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1480),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1490),
.A2(n_1461),
.B(n_1413),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1485),
.Y(n_1507)
);

OAI32xp33_ASAP7_75t_L g1508 ( 
.A1(n_1489),
.A2(n_1446),
.A3(n_1452),
.B1(n_1454),
.B2(n_1443),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1467),
.B(n_1451),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1467),
.B(n_1451),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1469),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1483),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1483),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1482),
.B(n_1492),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1500),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1500),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1475),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1493),
.B(n_1472),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1482),
.B(n_1451),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1497),
.Y(n_1520)
);

AOI32xp33_ASAP7_75t_L g1521 ( 
.A1(n_1466),
.A2(n_1460),
.A3(n_1440),
.B1(n_1457),
.B2(n_1441),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_SL g1523 ( 
.A(n_1472),
.B(n_1421),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1469),
.A2(n_1390),
.B1(n_1418),
.B2(n_1374),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1496),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1494),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1488),
.B(n_1456),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1501),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1488),
.B(n_1437),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1501),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_L g1531 ( 
.A(n_1494),
.B(n_1434),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1468),
.Y(n_1532)
);

AND4x1_ASAP7_75t_L g1533 ( 
.A(n_1466),
.B(n_1424),
.C(n_1460),
.D(n_1439),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1494),
.B(n_1444),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1476),
.B(n_1487),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1495),
.B(n_1437),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1476),
.B(n_1453),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1486),
.A2(n_1398),
.B1(n_1407),
.B2(n_1455),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1468),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1470),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1470),
.A2(n_1442),
.B(n_1446),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1477),
.B(n_1456),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1477),
.B(n_1456),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1487),
.B(n_1459),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1503),
.B(n_1474),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1512),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1534),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1534),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1522),
.B(n_1471),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1505),
.B(n_1471),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1518),
.B(n_1535),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1535),
.B(n_1487),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1517),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1537),
.B(n_1498),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1513),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1516),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1511),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1511),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1507),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1514),
.B(n_1479),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1532),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1509),
.B(n_1446),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1539),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1504),
.B(n_1498),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1540),
.Y(n_1569)
);

INVx8_ASAP7_75t_L g1570 ( 
.A(n_1534),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_R g1571 ( 
.A(n_1523),
.B(n_1264),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1502),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1534),
.B(n_1473),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1502),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1520),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1506),
.A2(n_1499),
.B1(n_1473),
.B2(n_1455),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1526),
.B(n_1473),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1520),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1240),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1571),
.A2(n_1508),
.B1(n_1524),
.B2(n_1531),
.C(n_1521),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1545),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1563),
.B(n_1525),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1538),
.Y(n_1585)
);

NOR4xp25_ASAP7_75t_SL g1586 ( 
.A(n_1545),
.B(n_1533),
.C(n_1442),
.D(n_1531),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1546),
.B(n_1510),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1547),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1562),
.A2(n_1524),
.B(n_1526),
.C(n_1544),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1547),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1552),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1499),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1552),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1556),
.A2(n_1574),
.B(n_1573),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1519),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1546),
.A2(n_1544),
.B1(n_1527),
.B2(n_1542),
.C(n_1543),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

O2A1O1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1555),
.A2(n_1452),
.B(n_1454),
.C(n_1530),
.Y(n_1598)
);

AOI221x1_ASAP7_75t_L g1599 ( 
.A1(n_1555),
.A2(n_1528),
.B1(n_1460),
.B2(n_1455),
.C(n_1408),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1570),
.A2(n_1281),
.B(n_1452),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1578),
.A2(n_1435),
.B(n_1460),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1559),
.Y(n_1602)
);

AOI321xp33_ASAP7_75t_L g1603 ( 
.A1(n_1554),
.A2(n_1439),
.A3(n_1484),
.B1(n_1536),
.B2(n_1529),
.C(n_1454),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1561),
.B(n_1499),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1570),
.A2(n_1282),
.B(n_1222),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1559),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1605),
.B(n_1568),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1604),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1587),
.B(n_1551),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1594),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1597),
.B(n_1561),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1594),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1604),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1592),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1583),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_L g1617 ( 
.A(n_1582),
.B(n_1549),
.C(n_1548),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1586),
.B(n_1554),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1596),
.A2(n_1570),
.B1(n_1568),
.B2(n_1548),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1600),
.B(n_1548),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1558),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1601),
.A2(n_1570),
.B1(n_1549),
.B2(n_1575),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1590),
.B(n_1549),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

BUFx4f_ASAP7_75t_SL g1625 ( 
.A(n_1581),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1617),
.A2(n_1589),
.B1(n_1598),
.B2(n_1591),
.C(n_1593),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1616),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1613),
.B(n_1606),
.Y(n_1628)
);

OAI211xp5_ASAP7_75t_L g1629 ( 
.A1(n_1610),
.A2(n_1612),
.B(n_1619),
.C(n_1603),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1610),
.A2(n_1570),
.B(n_1595),
.C(n_1556),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1623),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1612),
.A2(n_1595),
.B1(n_1584),
.B2(n_1556),
.C(n_1574),
.Y(n_1632)
);

AND4x1_ASAP7_75t_SL g1633 ( 
.A(n_1622),
.B(n_1584),
.C(n_1551),
.D(n_1564),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1560),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1623),
.Y(n_1635)
);

AOI222xp33_ASAP7_75t_L g1636 ( 
.A1(n_1618),
.A2(n_1574),
.B1(n_1573),
.B2(n_1560),
.C1(n_1567),
.C2(n_1565),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1631),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1635),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1636),
.B(n_1618),
.C(n_1611),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1627),
.Y(n_1640)
);

AOI311xp33_ASAP7_75t_L g1641 ( 
.A1(n_1629),
.A2(n_1624),
.A3(n_1607),
.B(n_1621),
.C(n_1615),
.Y(n_1641)
);

AND4x1_ASAP7_75t_L g1642 ( 
.A(n_1636),
.B(n_1620),
.C(n_1625),
.D(n_1599),
.Y(n_1642)
);

AOI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1626),
.A2(n_1620),
.B(n_1609),
.C(n_1614),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1628),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1632),
.A2(n_1614),
.B1(n_1634),
.B2(n_1616),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1630),
.Y(n_1646)
);

OAI211xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1643),
.A2(n_1633),
.B(n_1609),
.C(n_1573),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1639),
.A2(n_1567),
.B(n_1565),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1646),
.B(n_1576),
.C(n_1572),
.Y(n_1649)
);

NOR4xp25_ASAP7_75t_L g1650 ( 
.A(n_1641),
.B(n_1577),
.C(n_1576),
.D(n_1580),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1637),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_L g1652 ( 
.A(n_1644),
.B(n_1580),
.C(n_1572),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1648),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1647),
.A2(n_1638),
.B1(n_1645),
.B2(n_1640),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1651),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1650),
.Y(n_1656)
);

OA22x2_ASAP7_75t_L g1657 ( 
.A1(n_1649),
.A2(n_1638),
.B1(n_1642),
.B2(n_1569),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1652),
.B(n_1575),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1651),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1658),
.B(n_1228),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_SL g1661 ( 
.A(n_1654),
.B(n_1435),
.C(n_1298),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1655),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1659),
.B(n_1579),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1657),
.A2(n_1569),
.B(n_1577),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1663),
.Y(n_1665)
);

XNOR2xp5_ASAP7_75t_L g1666 ( 
.A(n_1661),
.B(n_1653),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1662),
.Y(n_1667)
);

XOR2xp5_ASAP7_75t_L g1668 ( 
.A(n_1666),
.B(n_1653),
.Y(n_1668)
);

AND4x2_ASAP7_75t_L g1669 ( 
.A(n_1668),
.B(n_1664),
.C(n_1660),
.D(n_1656),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1669),
.B(n_1665),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1669),
.A2(n_1667),
.B1(n_1577),
.B2(n_1298),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1670),
.B(n_1564),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1670),
.Y(n_1673)
);

OA22x2_ASAP7_75t_L g1674 ( 
.A1(n_1672),
.A2(n_1579),
.B1(n_1550),
.B2(n_1233),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1673),
.B(n_1550),
.Y(n_1675)
);

OAI21xp33_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1566),
.B(n_1327),
.Y(n_1676)
);

XNOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1676),
.B(n_1674),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1566),
.B1(n_1357),
.B2(n_1353),
.Y(n_1678)
);

AOI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1320),
.B(n_1327),
.C(n_1353),
.Y(n_1679)
);


endmodule