module fake_jpeg_9532_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_33),
.Y(n_55)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_34),
.B1(n_24),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_52),
.B1(n_62),
.B2(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_34),
.B1(n_24),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_34),
.B1(n_24),
.B2(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_59),
.Y(n_89)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_30),
.B1(n_33),
.B2(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_30),
.B1(n_33),
.B2(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_81),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_39),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_27),
.B(n_29),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_22),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_32),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_86),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_41),
.C(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_41),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_32),
.Y(n_88)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_91),
.Y(n_123)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_22),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_96),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_103),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_23),
.Y(n_99)
);

NOR2x1_ASAP7_75t_R g119 ( 
.A(n_99),
.B(n_102),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_78),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_0),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_114),
.B(n_124),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_110),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_38),
.B1(n_37),
.B2(n_19),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_108),
.A2(n_122),
.B1(n_131),
.B2(n_98),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_0),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_1),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_134),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_85),
.B(n_99),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_141),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_140),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_80),
.B1(n_90),
.B2(n_74),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_129),
.B1(n_124),
.B2(n_96),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_120),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_70),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_160),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_84),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_114),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_79),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_125),
.B(n_105),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_165),
.B(n_173),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_131),
.B1(n_127),
.B2(n_130),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_176),
.B1(n_179),
.B2(n_185),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_131),
.B1(n_114),
.B2(n_122),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_181),
.B(n_196),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_148),
.B1(n_139),
.B2(n_163),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_114),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_186),
.B(n_111),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_105),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_104),
.A3(n_93),
.B1(n_80),
.B2(n_102),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_112),
.C(n_100),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_193),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_133),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_137),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_139),
.A2(n_83),
.B1(n_89),
.B2(n_91),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_153),
.B1(n_141),
.B2(n_134),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_78),
.B(n_100),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_199),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_145),
.C(n_142),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_162),
.C(n_158),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_201),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_132),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_210),
.B(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_212),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_159),
.B(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_136),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_223),
.B1(n_186),
.B2(n_183),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_159),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_172),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_89),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_89),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_222),
.A2(n_217),
.B1(n_201),
.B2(n_183),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_112),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_237),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_226),
.B(n_227),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_193),
.C(n_174),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_236),
.C(n_240),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_185),
.B1(n_187),
.B2(n_192),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_231),
.B1(n_206),
.B2(n_197),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_187),
.B1(n_175),
.B2(n_178),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_245),
.B1(n_222),
.B2(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_184),
.C(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_212),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_170),
.C(n_176),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_190),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_216),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_86),
.B1(n_113),
.B2(n_107),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_247),
.C(n_249),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_202),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_208),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_256),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_254),
.B1(n_244),
.B2(n_245),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_215),
.B(n_210),
.C(n_209),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_208),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_205),
.C(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_205),
.C(n_113),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_262),
.Y(n_276)
);

AOI32xp33_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_18),
.A3(n_16),
.B1(n_113),
.B2(n_27),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_107),
.B1(n_71),
.B2(n_82),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_269),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_238),
.B1(n_261),
.B2(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_230),
.B1(n_226),
.B2(n_229),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_275),
.C(n_16),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_243),
.B1(n_227),
.B2(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_107),
.B1(n_92),
.B2(n_3),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_9),
.B(n_15),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_9),
.B(n_11),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_275),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_247),
.B1(n_249),
.B2(n_256),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_287),
.B1(n_6),
.B2(n_12),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_8),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_27),
.C(n_7),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_289),
.B(n_291),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_1),
.B(n_2),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_8),
.B(n_13),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_276),
.B(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_274),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_288),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_277),
.B1(n_10),
.B2(n_4),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_27),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_300),
.C(n_291),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_301),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_6),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_289),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_4),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_292),
.A3(n_295),
.B1(n_296),
.B2(n_298),
.C1(n_6),
.C2(n_11),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_280),
.B(n_10),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_4),
.A3(n_5),
.B1(n_12),
.B2(n_13),
.C1(n_2),
.C2(n_3),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

AOI321xp33_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_308),
.A3(n_311),
.B1(n_302),
.B2(n_303),
.C(n_5),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_314),
.B(n_2),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_2),
.Y(n_317)
);


endmodule