module real_jpeg_18057_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AO22x1_ASAP7_75t_SL g10 ( 
.A1(n_0),
.A2(n_1),
.B1(n_11),
.B2(n_12),
.Y(n_10)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

OA22x2_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_4),
.B1(n_12),
.B2(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_18),
.Y(n_29)
);

OR2x4_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_10),
.Y(n_9)
);

INVx2_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

AOI221xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.C(n_27),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_8),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_13),
.Y(n_8)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_15),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

OR2x4_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);


endmodule