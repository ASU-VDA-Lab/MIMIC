module fake_jpeg_18793_n_227 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_10),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_20),
.B1(n_14),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_44),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_54),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_23),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_32),
.B1(n_25),
.B2(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_27),
.B1(n_26),
.B2(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_54),
.C(n_52),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_51),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_64),
.B1(n_70),
.B2(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_74),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_36),
.B1(n_38),
.B2(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_41),
.C(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_90),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_51),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_73),
.C(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_89),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_21),
.B(n_15),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_87),
.B(n_61),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_50),
.B(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_38),
.B1(n_50),
.B2(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_94),
.B1(n_76),
.B2(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_37),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_64),
.B1(n_69),
.B2(n_66),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_93),
.B1(n_84),
.B2(n_26),
.Y(n_124)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_69),
.B1(n_66),
.B2(n_68),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_69),
.B(n_67),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_115),
.B(n_81),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_67),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_99),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_72),
.B1(n_18),
.B2(n_11),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_11),
.B1(n_18),
.B2(n_19),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_72),
.B(n_2),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_119),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_95),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

XOR2x2_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_82),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_123),
.B(n_102),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_93),
.B1(n_87),
.B2(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_128),
.B1(n_112),
.B2(n_114),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_27),
.C(n_40),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_127),
.C(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_40),
.C(n_16),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_48),
.B1(n_22),
.B2(n_21),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_33),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_16),
.C(n_33),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_16),
.C(n_104),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_16),
.B(n_10),
.C(n_17),
.D(n_23),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_137),
.B(n_102),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_1),
.B(n_2),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_13),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_150),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_152),
.B1(n_158),
.B2(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_109),
.B(n_96),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_96),
.C(n_108),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_143),
.C(n_149),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_101),
.B(n_48),
.C(n_23),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_101),
.B1(n_48),
.B2(n_22),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_118),
.B1(n_121),
.B2(n_135),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_158),
.B1(n_120),
.B2(n_160),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_156),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_127),
.C(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

XOR2x2_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_119),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_152),
.B(n_141),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_131),
.C(n_128),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_185),
.Y(n_198)
);

OA21x2_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_175),
.B(n_2),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_141),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_174),
.C(n_162),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_142),
.B(n_150),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_19),
.B1(n_18),
.B2(n_11),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_144),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_154),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_19),
.C(n_21),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_192),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_163),
.B(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_163),
.A3(n_158),
.B1(n_101),
.B2(n_172),
.C1(n_175),
.C2(n_17),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_197),
.B1(n_21),
.B2(n_15),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_187),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_203),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_183),
.B1(n_180),
.B2(n_177),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_190),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_210),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_191),
.A3(n_198),
.B1(n_194),
.B2(n_197),
.C1(n_177),
.C2(n_4),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_9),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_5),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_200),
.A3(n_199),
.B(n_7),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_6),
.B(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_5),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_6),
.B(n_7),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_218),
.Y(n_220)
);

INVxp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.B1(n_221),
.B2(n_207),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_214),
.C(n_209),
.Y(n_224)
);

OAI321xp33_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_219),
.A3(n_216),
.B1(n_9),
.B2(n_8),
.C(n_7),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_9),
.Y(n_227)
);


endmodule