module fake_jpeg_30301_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_2),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_61),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_37),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_60),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_38),
.C(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_0),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_12),
.Y(n_80)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_34),
.B1(n_16),
.B2(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_63),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_74),
.C(n_14),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_3),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_13),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

AOI21x1_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_95),
.C(n_96),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_92),
.B1(n_83),
.B2(n_89),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_81),
.A3(n_88),
.B1(n_78),
.B2(n_20),
.C1(n_23),
.C2(n_24),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_15),
.C(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_19),
.Y(n_104)
);


endmodule