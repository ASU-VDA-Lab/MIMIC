module fake_ibex_1032_n_1917 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_414, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_428, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_1917);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_428;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_1917;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_557;
wire n_641;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_545;
wire n_887;
wire n_1162;
wire n_1894;
wire n_634;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_1349;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_934;
wire n_520;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1900;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_352),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_75),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_160),
.Y(n_432)
);

BUFx8_ASAP7_75t_SL g433 ( 
.A(n_340),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_279),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_393),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_308),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_346),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_271),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_353),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_409),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_336),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_109),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_321),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_206),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_56),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_215),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_199),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_149),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_114),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_373),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_294),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_5),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_174),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_249),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_72),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_45),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_382),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_73),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_61),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_32),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_404),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_300),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_402),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_88),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_376),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_408),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_239),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_158),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_35),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_423),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_357),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_334),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_344),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_391),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_43),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_67),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_276),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_91),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_327),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_288),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_284),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_395),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_295),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_129),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_181),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_144),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_85),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_230),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_405),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_263),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_24),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_216),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_368),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_320),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_285),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_351),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_53),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_289),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_400),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_109),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_150),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_264),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_75),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_231),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_341),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_84),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_16),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_332),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_380),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_203),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_122),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_157),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_267),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_153),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_333),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_303),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_369),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_14),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_416),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_140),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_265),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_233),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_36),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_127),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_57),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_245),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_413),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_38),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_184),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_397),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_48),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_66),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_337),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_309),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_392),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_338),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_137),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_387),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_377),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_244),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_48),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_401),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_88),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_383),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_21),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_19),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_49),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_154),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_318),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_192),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_195),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_394),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_354),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_403),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_68),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_253),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_290),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_74),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_421),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_128),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_429),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_317),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_40),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_274),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_350),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_378),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_235),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_371),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_343),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_201),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_364),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_61),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_94),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_360),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_412),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_359),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_45),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_207),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_291),
.Y(n_592)
);

BUFx5_ASAP7_75t_L g593 ( 
.A(n_311),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_319),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_133),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_26),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_42),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_330),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_415),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_26),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_70),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_209),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_44),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_83),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_365),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_348),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_374),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_85),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_427),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_347),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_407),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_305),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_281),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_83),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_362),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_342),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_390),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_349),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_426),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_178),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_272),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_379),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_72),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_367),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_240),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_261),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_76),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_292),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_118),
.Y(n_629)
);

CKINVDCx14_ASAP7_75t_R g630 ( 
.A(n_262),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_171),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_145),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_251),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_43),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_180),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_324),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_177),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_247),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_386),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_191),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_197),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_91),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_385),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_68),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_37),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_226),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_194),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_2),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_277),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_51),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_417),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_15),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_217),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_210),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_313),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_59),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_298),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_389),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_142),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_372),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_384),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_64),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_2),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_104),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_19),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_169),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_420),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_13),
.Y(n_668)
);

CKINVDCx16_ASAP7_75t_R g669 ( 
.A(n_293),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_126),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_14),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_0),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_335),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_356),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_81),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_5),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_363),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_381),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_361),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_411),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_38),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_399),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_111),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_8),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_183),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_345),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_419),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_42),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_8),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_76),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_355),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_98),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_325),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_69),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_296),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_339),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_168),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_553),
.Y(n_698)
);

INVxp33_ASAP7_75t_SL g699 ( 
.A(n_664),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_433),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_601),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_553),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_461),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_585),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_588),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_588),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_664),
.Y(n_707)
);

INVxp33_ASAP7_75t_SL g708 ( 
.A(n_603),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_432),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_623),
.Y(n_710)
);

BUFx2_ASAP7_75t_SL g711 ( 
.A(n_440),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_446),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_431),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_503),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_576),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_458),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_584),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_466),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_519),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_560),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_444),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_593),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_468),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_441),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_502),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_538),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_488),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_512),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_515),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_543),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_552),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_569),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_595),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_606),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_597),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_628),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_631),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_634),
.Y(n_740)
);

CKINVDCx16_ASAP7_75t_R g741 ( 
.A(n_669),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_650),
.Y(n_742)
);

INVxp67_ASAP7_75t_SL g743 ( 
.A(n_652),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_662),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_668),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_684),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_687),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_689),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_587),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_593),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_587),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_442),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_518),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_674),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_674),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_443),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_445),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_448),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_449),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_450),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_462),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_456),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_457),
.Y(n_763)
);

CKINVDCx14_ASAP7_75t_R g764 ( 
.A(n_459),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_465),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_581),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_518),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_460),
.Y(n_768)
);

BUFx6f_ASAP7_75t_SL g769 ( 
.A(n_447),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_464),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_469),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_470),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_518),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_471),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_518),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_593),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_593),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_478),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_485),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_486),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_593),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_509),
.Y(n_782)
);

CKINVDCx11_ASAP7_75t_R g783 ( 
.A(n_472),
.Y(n_783)
);

INVxp33_ASAP7_75t_SL g784 ( 
.A(n_530),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_721),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_721),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_713),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_698),
.B(n_474),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_716),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_702),
.B(n_630),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_719),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_710),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_750),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_776),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_713),
.Y(n_796)
);

BUFx6f_ASAP7_75t_SL g797 ( 
.A(n_749),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_720),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_769),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_722),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_777),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_705),
.B(n_483),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_707),
.B(n_472),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_773),
.Y(n_804)
);

OA21x2_ASAP7_75t_L g805 ( 
.A1(n_781),
.A2(n_493),
.B(n_487),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_766),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_773),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_721),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_721),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_766),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_753),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_753),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_724),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_706),
.B(n_535),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_728),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_765),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_729),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_730),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_731),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_R g821 ( 
.A(n_764),
.B(n_430),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_704),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_767),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_737),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_740),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_742),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_767),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_775),
.Y(n_828)
);

AND2x6_ASAP7_75t_L g829 ( 
.A(n_756),
.B(n_498),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_712),
.B(n_594),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_757),
.B(n_537),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_744),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_715),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_769),
.B(n_620),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_709),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_782),
.Y(n_836)
);

CKINVDCx11_ASAP7_75t_R g837 ( 
.A(n_783),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_745),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_758),
.B(n_540),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_741),
.B(n_497),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_748),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_778),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_SL g845 ( 
.A1(n_726),
.A2(n_556),
.B1(n_558),
.B2(n_545),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_760),
.B(n_559),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_718),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_762),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_763),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_751),
.B(n_434),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_768),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_770),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_701),
.B(n_497),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_718),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_725),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_771),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_743),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_764),
.B(n_671),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_743),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_772),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_774),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_733),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_754),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_733),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_727),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_755),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_779),
.B(n_499),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_699),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_708),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_784),
.B(n_568),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_703),
.B(n_624),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_505),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_759),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_571),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_761),
.B(n_586),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_700),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_780),
.B(n_590),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_717),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_736),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_739),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_747),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_732),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_734),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_735),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_738),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_716),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_707),
.B(n_671),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_710),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_766),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_723),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_716),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_713),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_766),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_704),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_725),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_710),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_698),
.B(n_596),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_765),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_704),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_698),
.B(n_600),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_766),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_766),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_716),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_766),
.Y(n_904)
);

CKINVDCx8_ASAP7_75t_R g905 ( 
.A(n_711),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_716),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_711),
.B(n_508),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_721),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_698),
.B(n_516),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_721),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_716),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_699),
.A2(n_608),
.B1(n_614),
.B2(n_604),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_766),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_721),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_710),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_766),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_716),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_710),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_766),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_716),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_710),
.Y(n_921)
);

BUFx8_ASAP7_75t_L g922 ( 
.A(n_769),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_716),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_698),
.B(n_517),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_766),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_710),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_723),
.A2(n_525),
.B(n_452),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_704),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_713),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_725),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_SL g931 ( 
.A1(n_704),
.A2(n_642),
.B1(n_644),
.B2(n_627),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_716),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_766),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_SL g934 ( 
.A1(n_704),
.A2(n_648),
.B1(n_663),
.B2(n_645),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_804),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_889),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_889),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_927),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_807),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_893),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_876),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_907),
.B(n_521),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_893),
.Y(n_943)
);

BUFx4f_ASAP7_75t_L g944 ( 
.A(n_876),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_901),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_836),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_L g947 ( 
.A(n_796),
.B(n_672),
.C(n_665),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_847),
.B(n_438),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_901),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_813),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_854),
.B(n_484),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_902),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_813),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_902),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_913),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_863),
.B(n_435),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_913),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_916),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_862),
.B(n_436),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_864),
.B(n_437),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_813),
.Y(n_961)
);

INVxp67_ASAP7_75t_SL g962 ( 
.A(n_787),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_916),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_863),
.B(n_439),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_919),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_919),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_857),
.B(n_451),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_789),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_819),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_819),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_791),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_922),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_819),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_798),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_803),
.B(n_675),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_820),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_892),
.B(n_676),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_820),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_820),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_826),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_922),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_800),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_886),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_822),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_891),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_859),
.B(n_453),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_826),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_816),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_826),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_842),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_816),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_842),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_799),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_842),
.Y(n_994)
);

CKINVDCx16_ASAP7_75t_R g995 ( 
.A(n_894),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_849),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_903),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_906),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_849),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_806),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_797),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_810),
.Y(n_1002)
);

INVx11_ASAP7_75t_L g1003 ( 
.A(n_905),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_861),
.B(n_454),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_790),
.B(n_572),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_817),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_929),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_887),
.Y(n_1008)
);

CKINVDCx6p67_ASAP7_75t_R g1009 ( 
.A(n_883),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_849),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_851),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_851),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_868),
.A2(n_683),
.B1(n_688),
.B2(n_681),
.Y(n_1013)
);

OAI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_868),
.A2(n_692),
.B1(n_694),
.B2(n_690),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_797),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_851),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_852),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_852),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_852),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_861),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_805),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_890),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_890),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_833),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_805),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_863),
.B(n_455),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_833),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_911),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_898),
.Y(n_1029)
);

AND3x2_ASAP7_75t_L g1030 ( 
.A(n_882),
.B(n_544),
.C(n_536),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_844),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_917),
.Y(n_1032)
);

NAND2xp33_ASAP7_75t_SL g1033 ( 
.A(n_821),
.B(n_463),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_811),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_812),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_866),
.B(n_693),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_904),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_SL g1038 ( 
.A(n_855),
.B(n_895),
.C(n_865),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_920),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_823),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_827),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_828),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_788),
.B(n_467),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_788),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_802),
.B(n_473),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_843),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_850),
.B(n_475),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_923),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_799),
.B(n_476),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_932),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_792),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_888),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_802),
.B(n_477),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_869),
.B(n_0),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_909),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_925),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_831),
.A2(n_567),
.B(n_562),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_814),
.B(n_479),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_933),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_896),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_848),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_856),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_915),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_918),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_909),
.B(n_480),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_860),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_921),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_815),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_926),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_818),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_912),
.B(n_577),
.C(n_573),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_824),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_837),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_793),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_876),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_L g1076 ( 
.A(n_829),
.B(n_593),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_873),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_924),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_SL g1079 ( 
.A(n_907),
.B(n_482),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_924),
.A2(n_583),
.B1(n_598),
.B2(n_579),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_794),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_795),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_853),
.B(n_489),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_801),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_829),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_825),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_867),
.B(n_491),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_867),
.B(n_492),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_897),
.B(n_900),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_832),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_838),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_899),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_841),
.B(n_494),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_SL g1094 ( 
.A(n_885),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_928),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_839),
.B(n_495),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_829),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_829),
.Y(n_1098)
);

AOI22x1_ASAP7_75t_L g1099 ( 
.A1(n_785),
.A2(n_570),
.B1(n_574),
.B2(n_555),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_785),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_785),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_786),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_846),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_870),
.B(n_496),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_830),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_834),
.B(n_500),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_786),
.Y(n_1107)
);

OAI22xp33_ASAP7_75t_SL g1108 ( 
.A1(n_930),
.A2(n_610),
.B1(n_611),
.B2(n_607),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_875),
.B(n_1),
.Y(n_1109)
);

CKINVDCx16_ASAP7_75t_R g1110 ( 
.A(n_835),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_786),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_858),
.B(n_501),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_872),
.A2(n_615),
.B1(n_619),
.B2(n_613),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_840),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_808),
.Y(n_1115)
);

AND2x6_ASAP7_75t_L g1116 ( 
.A(n_878),
.B(n_629),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_874),
.B(n_506),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_877),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_L g1119 ( 
.A(n_880),
.B(n_507),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_808),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_808),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_809),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_809),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_872),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_879),
.B(n_633),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_809),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_908),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_883),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_908),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_908),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_910),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_871),
.B(n_510),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_910),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_910),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_914),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_914),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_883),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_914),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_881),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_845),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_884),
.B(n_637),
.C(n_636),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_931),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_934),
.B(n_511),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_847),
.A2(n_639),
.B1(n_670),
.B2(n_667),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_817),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_836),
.B(n_513),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_889),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_804),
.Y(n_1148)
);

AO22x2_ASAP7_75t_L g1149 ( 
.A1(n_884),
.A2(n_679),
.B1(n_680),
.B2(n_678),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_862),
.B(n_514),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_836),
.B(n_520),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_889),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_862),
.B(n_522),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_889),
.Y(n_1154)
);

AND2x6_ASAP7_75t_L g1155 ( 
.A(n_803),
.B(n_686),
.Y(n_1155)
);

NAND2xp33_ASAP7_75t_L g1156 ( 
.A(n_829),
.B(n_523),
.Y(n_1156)
);

OAI21xp33_ASAP7_75t_SL g1157 ( 
.A1(n_862),
.A2(n_640),
.B(n_605),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_836),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_847),
.B(n_526),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1158),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1072),
.B(n_527),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1020),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1140),
.A2(n_697),
.B1(n_661),
.B2(n_695),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_988),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1089),
.B(n_528),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1029),
.B(n_1),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1007),
.A2(n_531),
.B1(n_533),
.B2(n_529),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1097),
.A2(n_539),
.B1(n_542),
.B2(n_534),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_988),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1097),
.B(n_696),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1145),
.B(n_3),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1020),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1085),
.B(n_546),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1085),
.B(n_691),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1118),
.B(n_547),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_975),
.B(n_548),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1103),
.B(n_549),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1085),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1077),
.B(n_3),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_935),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1068),
.B(n_550),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_935),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_991),
.Y(n_1183)
);

INVx8_ASAP7_75t_L g1184 ( 
.A(n_942),
.Y(n_1184)
);

BUFx5_ASAP7_75t_L g1185 ( 
.A(n_1025),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1079),
.B(n_685),
.Y(n_1186)
);

NAND2xp33_ASAP7_75t_L g1187 ( 
.A(n_1021),
.B(n_551),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_939),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_939),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_L g1190 ( 
.A(n_1021),
.B(n_557),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_991),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1148),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1044),
.A2(n_563),
.B1(n_564),
.B2(n_561),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_975),
.B(n_565),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1148),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1031),
.B(n_4),
.Y(n_1196)
);

AND2x6_ASAP7_75t_SL g1197 ( 
.A(n_1073),
.B(n_4),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1068),
.B(n_566),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1006),
.A2(n_578),
.B1(n_580),
.B2(n_575),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1024),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_968),
.B(n_582),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_971),
.B(n_589),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_946),
.B(n_6),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1070),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1086),
.Y(n_1205)
);

AO221x1_ASAP7_75t_L g1206 ( 
.A1(n_1149),
.A2(n_490),
.B1(n_504),
.B2(n_481),
.C(n_444),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1055),
.B(n_682),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1078),
.B(n_591),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_L g1209 ( 
.A(n_1114),
.B(n_1038),
.C(n_995),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_974),
.B(n_599),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1091),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1008),
.B(n_602),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_972),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1021),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1098),
.B(n_677),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_982),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_947),
.B(n_612),
.C(n_609),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1024),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1098),
.B(n_616),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_962),
.B(n_6),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_977),
.B(n_7),
.Y(n_1221)
);

NAND2xp33_ASAP7_75t_L g1222 ( 
.A(n_1025),
.B(n_617),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1125),
.B(n_7),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1125),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_993),
.B(n_9),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_L g1226 ( 
.A(n_1116),
.B(n_618),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1139),
.B(n_673),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1155),
.A2(n_1124),
.B1(n_1113),
.B2(n_1083),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_983),
.B(n_622),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1114),
.B(n_9),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_981),
.B(n_625),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_993),
.B(n_10),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_985),
.B(n_626),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_997),
.Y(n_1234)
);

INVx5_ASAP7_75t_L g1235 ( 
.A(n_1001),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_L g1236 ( 
.A(n_1128),
.B(n_10),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1155),
.A2(n_635),
.B1(n_638),
.B2(n_632),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_998),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_L g1239 ( 
.A(n_1116),
.B(n_643),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1028),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1110),
.B(n_11),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1124),
.B(n_646),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_R g1243 ( 
.A(n_1095),
.B(n_647),
.Y(n_1243)
);

AND2x6_ASAP7_75t_SL g1244 ( 
.A(n_942),
.B(n_11),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1032),
.B(n_649),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1155),
.A2(n_641),
.B1(n_653),
.B2(n_651),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1039),
.B(n_654),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1139),
.B(n_666),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1048),
.B(n_655),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1087),
.B(n_657),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1050),
.Y(n_1251)
);

NAND2x1_ASAP7_75t_L g1252 ( 
.A(n_1022),
.B(n_444),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1080),
.A2(n_659),
.B1(n_660),
.B2(n_658),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1090),
.B(n_12),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1128),
.B(n_12),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1061),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1155),
.A2(n_481),
.B1(n_490),
.B2(n_444),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1105),
.B(n_1043),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1109),
.B(n_481),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1096),
.B(n_481),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1053),
.B(n_490),
.Y(n_1261)
);

NOR2xp67_ASAP7_75t_SL g1262 ( 
.A(n_1059),
.B(n_490),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1149),
.A2(n_524),
.B1(n_532),
.B2(n_504),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1088),
.B(n_13),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1061),
.B(n_15),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_948),
.A2(n_524),
.B1(n_532),
.B2(n_504),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1062),
.B(n_16),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1062),
.B(n_17),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1001),
.B(n_17),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1066),
.B(n_18),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1066),
.B(n_18),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1022),
.A2(n_524),
.B(n_532),
.C(n_504),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_958),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1027),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_951),
.B(n_20),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1054),
.B(n_20),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_958),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_959),
.B(n_524),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_L g1279 ( 
.A(n_1116),
.B(n_532),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1036),
.B(n_1005),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1023),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_984),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_L g1283 ( 
.A(n_1108),
.B(n_21),
.C(n_22),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_960),
.B(n_541),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1092),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1045),
.B(n_22),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1023),
.Y(n_1287)
);

AND2x6_ASAP7_75t_SL g1288 ( 
.A(n_1143),
.B(n_23),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_965),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1159),
.B(n_23),
.Y(n_1290)
);

OR2x6_ASAP7_75t_L g1291 ( 
.A(n_1142),
.B(n_541),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1065),
.B(n_24),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1013),
.B(n_25),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1150),
.B(n_541),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1058),
.B(n_25),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1071),
.B(n_27),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1153),
.B(n_1015),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1116),
.B(n_27),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1003),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1137),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1027),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1057),
.B(n_967),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1051),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1075),
.B(n_541),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1157),
.A2(n_621),
.B(n_592),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1057),
.B(n_28),
.Y(n_1306)
);

OAI22x1_ASAP7_75t_SL g1307 ( 
.A1(n_1009),
.A2(n_1015),
.B1(n_1094),
.B2(n_1030),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_986),
.B(n_28),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1052),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1112),
.B(n_29),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_941),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_965),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1144),
.B(n_29),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1004),
.B(n_30),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1093),
.B(n_30),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1141),
.A2(n_621),
.B1(n_592),
.B2(n_33),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1060),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1014),
.B(n_592),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1063),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1034),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1067),
.B(n_31),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1067),
.B(n_31),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1037),
.B(n_32),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1064),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1074),
.A2(n_621),
.B(n_592),
.Y(n_1325)
);

NOR3xp33_ASAP7_75t_L g1326 ( 
.A(n_1146),
.B(n_33),
.C(n_34),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1151),
.B(n_34),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1069),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1037),
.B(n_35),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1049),
.B(n_36),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1035),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1040),
.Y(n_1332)
);

NAND2xp33_ASAP7_75t_SL g1333 ( 
.A(n_1132),
.B(n_621),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1119),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1152),
.B(n_39),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1000),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1152),
.B(n_41),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1002),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1041),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1056),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1056),
.B(n_41),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1106),
.B(n_44),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1042),
.Y(n_1343)
);

NAND2xp33_ASAP7_75t_L g1344 ( 
.A(n_999),
.B(n_112),
.Y(n_1344)
);

OR2x2_ASAP7_75t_SL g1345 ( 
.A(n_1094),
.B(n_46),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_SL g1346 ( 
.A(n_941),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1204),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1160),
.B(n_1282),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1199),
.B(n_1224),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1258),
.B(n_1104),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1231),
.B(n_944),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1235),
.B(n_1185),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1235),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1285),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1225),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1184),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1185),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1185),
.Y(n_1358)
);

INVxp33_ASAP7_75t_SL g1359 ( 
.A(n_1243),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1185),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1205),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1223),
.B(n_944),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1235),
.B(n_936),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1185),
.B(n_1033),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1293),
.A2(n_940),
.B1(n_943),
.B2(n_937),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1211),
.B(n_945),
.Y(n_1366)
);

OR2x2_ASAP7_75t_SL g1367 ( 
.A(n_1241),
.B(n_949),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1216),
.Y(n_1368)
);

AND2x2_ASAP7_75t_SL g1369 ( 
.A(n_1279),
.B(n_1156),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1180),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1182),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1184),
.B(n_999),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1234),
.B(n_952),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1238),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1184),
.B(n_1117),
.Y(n_1375)
);

BUFx5_ASAP7_75t_L g1376 ( 
.A(n_1162),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1307),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1213),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1225),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1188),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1189),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1307),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1178),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1283),
.A2(n_955),
.B1(n_957),
.B2(n_954),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1228),
.B(n_1047),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1240),
.B(n_1251),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1192),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1297),
.B(n_963),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1195),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1346),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1320),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1232),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1280),
.B(n_966),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1167),
.B(n_999),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1281),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1287),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1221),
.B(n_1046),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1172),
.B(n_1147),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1220),
.B(n_1154),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1301),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1176),
.B(n_956),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1165),
.B(n_1081),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1237),
.B(n_1016),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1196),
.B(n_1082),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1291),
.B(n_964),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1232),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1291),
.A2(n_1084),
.B1(n_1026),
.B2(n_1076),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1304),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1331),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1299),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1203),
.B(n_950),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1230),
.B(n_950),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1256),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_R g1414 ( 
.A(n_1346),
.B(n_46),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1166),
.B(n_47),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1171),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1343),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1244),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1332),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1323),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1179),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1274),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1175),
.B(n_1016),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1276),
.B(n_953),
.Y(n_1424)
);

INVx5_ASAP7_75t_L g1425 ( 
.A(n_1304),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1339),
.Y(n_1426)
);

BUFx4f_ASAP7_75t_L g1427 ( 
.A(n_1269),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1329),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1265),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1300),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1178),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1323),
.A2(n_953),
.B1(n_978),
.B2(n_961),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1311),
.B(n_1016),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1303),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1309),
.Y(n_1435)
);

INVx5_ASAP7_75t_L g1436 ( 
.A(n_1178),
.Y(n_1436)
);

NAND2xp33_ASAP7_75t_L g1437 ( 
.A(n_1302),
.B(n_938),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1340),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1267),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1194),
.B(n_1212),
.Y(n_1440)
);

INVx5_ASAP7_75t_L g1441 ( 
.A(n_1197),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1177),
.B(n_961),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1214),
.A2(n_938),
.B(n_978),
.Y(n_1443)
);

AND3x1_ASAP7_75t_SL g1444 ( 
.A(n_1345),
.B(n_47),
.C(n_49),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1250),
.B(n_989),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1286),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1340),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1209),
.A2(n_989),
.B1(n_996),
.B2(n_990),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1292),
.B(n_1310),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_L g1450 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1207),
.B(n_990),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1324),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1208),
.B(n_996),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1264),
.B(n_1010),
.Y(n_1454)
);

NAND2xp33_ASAP7_75t_L g1455 ( 
.A(n_1328),
.B(n_938),
.Y(n_1455)
);

NOR2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1298),
.B(n_1010),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1336),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1161),
.B(n_1017),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1268),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1270),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1273),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_L g1462 ( 
.A(n_1263),
.B(n_1017),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1168),
.B(n_1018),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1334),
.A2(n_1018),
.B1(n_970),
.B2(n_973),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1338),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1341),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1313),
.A2(n_976),
.B1(n_979),
.B2(n_969),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1271),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1181),
.B(n_980),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1186),
.Y(n_1470)
);

NAND2xp33_ASAP7_75t_L g1471 ( 
.A(n_1198),
.B(n_987),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1327),
.B(n_992),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1254),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1164),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1273),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1201),
.B(n_994),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1277),
.B(n_1011),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1277),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1169),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1202),
.B(n_1210),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1229),
.B(n_1012),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1233),
.B(n_1019),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1321),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1289),
.B(n_1126),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1245),
.B(n_50),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1253),
.B(n_50),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1247),
.B(n_51),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1249),
.B(n_52),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1193),
.B(n_1122),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1183),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1385),
.A2(n_1326),
.B1(n_1318),
.B2(n_1296),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1383),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1437),
.A2(n_1259),
.B(n_1222),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_R g1494 ( 
.A(n_1354),
.B(n_1226),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1359),
.A2(n_1242),
.B1(n_1239),
.B2(n_1275),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1377),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1440),
.A2(n_1290),
.B1(n_1308),
.B2(n_1315),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1430),
.Y(n_1498)
);

NOR2x1_ASAP7_75t_L g1499 ( 
.A(n_1356),
.B(n_1236),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1348),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1386),
.B(n_1246),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1347),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1356),
.B(n_1191),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1421),
.A2(n_1342),
.B1(n_1295),
.B2(n_1314),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1386),
.B(n_1163),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1355),
.B(n_1305),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1361),
.B(n_1330),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1449),
.A2(n_1306),
.B(n_1322),
.C(n_1335),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1368),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1480),
.A2(n_1316),
.B(n_1266),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_SL g1511 ( 
.A(n_1382),
.B(n_1410),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1379),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1446),
.A2(n_1255),
.B1(n_1227),
.B2(n_1248),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1353),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1393),
.A2(n_1337),
.B(n_1325),
.C(n_1333),
.Y(n_1515)
);

OR2x6_ASAP7_75t_L g1516 ( 
.A(n_1390),
.B(n_1405),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1416),
.A2(n_1206),
.B1(n_1217),
.B2(n_1289),
.Y(n_1517)
);

O2A1O1Ixp5_ASAP7_75t_SL g1518 ( 
.A1(n_1489),
.A2(n_1278),
.B(n_1294),
.C(n_1284),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1408),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1455),
.A2(n_1260),
.B(n_1261),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1486),
.A2(n_1312),
.B1(n_1218),
.B2(n_1200),
.Y(n_1521)
);

BUFx12f_ASAP7_75t_L g1522 ( 
.A(n_1390),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1471),
.A2(n_1443),
.B(n_1439),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1370),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1392),
.B(n_1312),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1357),
.A2(n_1252),
.B(n_1257),
.Y(n_1526)
);

O2A1O1Ixp5_ASAP7_75t_L g1527 ( 
.A1(n_1364),
.A2(n_1272),
.B(n_1173),
.C(n_1174),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1420),
.B(n_52),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1429),
.A2(n_1190),
.B(n_1187),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1414),
.Y(n_1530)
);

AO22x1_ASAP7_75t_L g1531 ( 
.A1(n_1441),
.A2(n_1288),
.B1(n_55),
.B2(n_53),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1415),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1358),
.A2(n_1099),
.B(n_1126),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1374),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1378),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1371),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1387),
.B(n_1170),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1408),
.B(n_1215),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1380),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1418),
.B(n_54),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1384),
.A2(n_1219),
.B1(n_1099),
.B2(n_1344),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1459),
.A2(n_1111),
.B(n_1107),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1408),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1460),
.A2(n_1111),
.B(n_1115),
.C(n_1107),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1441),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1391),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1349),
.B(n_54),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1406),
.B(n_1362),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1425),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1441),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1427),
.B(n_55),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1367),
.B(n_56),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1363),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1389),
.B(n_57),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1350),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1381),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1468),
.A2(n_1127),
.B1(n_1134),
.B2(n_1115),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1450),
.A2(n_1134),
.B(n_1127),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1432),
.A2(n_1133),
.B1(n_1138),
.B2(n_1122),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1397),
.A2(n_1133),
.B1(n_1138),
.B2(n_1122),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1383),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1425),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1473),
.A2(n_1262),
.B(n_1101),
.C(n_1102),
.Y(n_1563)
);

NAND2x1p5_ASAP7_75t_L g1564 ( 
.A(n_1425),
.B(n_1133),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1376),
.B(n_1138),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1413),
.B(n_58),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1376),
.B(n_1100),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1442),
.A2(n_1136),
.B(n_1121),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1375),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1405),
.B(n_58),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1485),
.A2(n_1487),
.B(n_1488),
.C(n_1483),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1404),
.A2(n_1123),
.B1(n_1129),
.B2(n_1120),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1403),
.A2(n_1135),
.B(n_1131),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1409),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1419),
.B(n_59),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1375),
.B(n_60),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1401),
.B(n_60),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1395),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1470),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1428),
.B(n_62),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1352),
.Y(n_1581)
);

O2A1O1Ixp33_ASAP7_75t_SL g1582 ( 
.A1(n_1538),
.A2(n_1372),
.B(n_1351),
.C(n_1394),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1508),
.A2(n_1571),
.B(n_1523),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1500),
.B(n_1426),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1555),
.B(n_1422),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1498),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1533),
.A2(n_1431),
.B(n_1360),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1570),
.B(n_1388),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1577),
.A2(n_1552),
.B(n_1532),
.C(n_1505),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1515),
.A2(n_1493),
.B(n_1369),
.Y(n_1590)
);

AOI31xp67_ASAP7_75t_L g1591 ( 
.A1(n_1504),
.A2(n_1565),
.A3(n_1423),
.B(n_1567),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1502),
.B(n_1366),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1509),
.Y(n_1593)
);

O2A1O1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1547),
.A2(n_1402),
.B(n_1399),
.C(n_1466),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1510),
.A2(n_1464),
.B(n_1365),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1579),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1556),
.B(n_1457),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1569),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1576),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1534),
.B(n_1366),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1546),
.B(n_1373),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1373),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1560),
.A2(n_1462),
.B(n_1412),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1524),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1526),
.A2(n_1431),
.B(n_1433),
.Y(n_1605)
);

AOI31xp67_ASAP7_75t_L g1606 ( 
.A1(n_1513),
.A2(n_1463),
.A3(n_1396),
.B(n_1467),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1518),
.A2(n_1438),
.B(n_1456),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1551),
.A2(n_1499),
.B(n_1495),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1559),
.A2(n_1573),
.B(n_1520),
.Y(n_1609)
);

AO31x2_ASAP7_75t_L g1610 ( 
.A1(n_1544),
.A2(n_1454),
.A3(n_1458),
.B(n_1469),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1558),
.A2(n_1568),
.B(n_1527),
.Y(n_1611)
);

AO31x2_ASAP7_75t_L g1612 ( 
.A1(n_1529),
.A2(n_1563),
.A3(n_1507),
.B(n_1566),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1564),
.A2(n_1438),
.B(n_1400),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1497),
.A2(n_1445),
.B(n_1453),
.C(n_1451),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1536),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1517),
.A2(n_1407),
.B(n_1444),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1539),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1519),
.B(n_1376),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1501),
.B(n_1465),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1570),
.A2(n_1424),
.B1(n_1411),
.B2(n_1448),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1553),
.B(n_1461),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1576),
.A2(n_1521),
.B1(n_1548),
.B2(n_1506),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1542),
.A2(n_1398),
.B(n_1476),
.Y(n_1623)
);

OAI22x1_ASAP7_75t_L g1624 ( 
.A1(n_1530),
.A2(n_1363),
.B1(n_1478),
.B2(n_1461),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1543),
.A2(n_1482),
.B(n_1481),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1512),
.B(n_1417),
.Y(n_1626)
);

O2A1O1Ixp5_ASAP7_75t_SL g1627 ( 
.A1(n_1543),
.A2(n_1472),
.B(n_1376),
.C(n_115),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1491),
.A2(n_1388),
.B(n_1434),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1580),
.B(n_1435),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1622),
.A2(n_1516),
.B1(n_1554),
.B2(n_1562),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1583),
.A2(n_1575),
.B(n_1541),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1586),
.Y(n_1633)
);

AO21x2_ASAP7_75t_L g1634 ( 
.A1(n_1590),
.A2(n_1537),
.B(n_1572),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1616),
.B(n_1516),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1599),
.A2(n_1519),
.B1(n_1549),
.B2(n_1511),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1611),
.A2(n_1557),
.B(n_1578),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1609),
.A2(n_1549),
.B(n_1452),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1587),
.A2(n_1605),
.B(n_1625),
.Y(n_1639)
);

CKINVDCx11_ASAP7_75t_R g1640 ( 
.A(n_1596),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_1525),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1436),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1584),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1608),
.B(n_1531),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1618),
.B(n_1522),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1604),
.B(n_1492),
.Y(n_1646)
);

CKINVDCx9p33_ASAP7_75t_R g1647 ( 
.A(n_1598),
.Y(n_1647)
);

AND2x6_ASAP7_75t_L g1648 ( 
.A(n_1581),
.B(n_1492),
.Y(n_1648)
);

BUFx2_ASAP7_75t_SL g1649 ( 
.A(n_1621),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1595),
.A2(n_1528),
.B(n_1479),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1620),
.A2(n_1514),
.B1(n_1503),
.B2(n_1447),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1603),
.A2(n_1490),
.B(n_1474),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1615),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1617),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1588),
.B(n_1535),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1503),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1627),
.A2(n_1561),
.B(n_1492),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1597),
.B(n_62),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1607),
.A2(n_1561),
.B(n_1130),
.Y(n_1659)
);

INVx5_ASAP7_75t_L g1660 ( 
.A(n_1581),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1613),
.A2(n_1561),
.B(n_1436),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1623),
.A2(n_1436),
.B(n_1383),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1614),
.A2(n_1478),
.B1(n_1550),
.B2(n_1545),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1644),
.A2(n_1589),
.B(n_1594),
.C(n_1585),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1643),
.B(n_1619),
.Y(n_1665)
);

O2A1O1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1644),
.A2(n_1600),
.B(n_1601),
.C(n_1592),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1656),
.B(n_1602),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1653),
.B(n_1628),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1644),
.A2(n_1629),
.B1(n_1475),
.B2(n_1496),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1632),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1633),
.B(n_1658),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1635),
.B(n_1612),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1646),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1635),
.B(n_1612),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1654),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1649),
.B(n_1612),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_SL g1680 ( 
.A(n_1645),
.B(n_1624),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1635),
.B(n_1610),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1663),
.A2(n_1540),
.B(n_1591),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1663),
.A2(n_1475),
.B(n_1484),
.C(n_1477),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1651),
.A2(n_1475),
.B1(n_1484),
.B2(n_1477),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1630),
.A2(n_1494),
.B1(n_1582),
.B2(n_1606),
.Y(n_1685)
);

O2A1O1Ixp5_ASAP7_75t_L g1686 ( 
.A1(n_1631),
.A2(n_116),
.B(n_117),
.C(n_113),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1655),
.B(n_63),
.Y(n_1687)
);

AOI21x1_ASAP7_75t_SL g1688 ( 
.A1(n_1647),
.A2(n_63),
.B(n_64),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1645),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1631),
.A2(n_65),
.B(n_66),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1630),
.A2(n_69),
.B1(n_65),
.B2(n_67),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1662),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1665),
.B(n_1660),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1692),
.A2(n_1659),
.B(n_1639),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1677),
.B(n_1676),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1675),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1672),
.B(n_1645),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1678),
.B(n_1650),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1673),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1670),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1679),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1672),
.Y(n_1702)
);

AO21x2_ASAP7_75t_L g1703 ( 
.A1(n_1692),
.A2(n_1652),
.B(n_1638),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1673),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1668),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1674),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1691),
.A2(n_1634),
.B1(n_1636),
.B2(n_1648),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1674),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1681),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1683),
.A2(n_1657),
.B(n_1661),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1669),
.A2(n_1634),
.B1(n_1648),
.B2(n_1650),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1689),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1667),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1664),
.B(n_1640),
.C(n_70),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1705),
.B(n_1671),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1700),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1666),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1713),
.B(n_1652),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1700),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1699),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1697),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1704),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1680),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1683),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1713),
.B(n_1660),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1714),
.A2(n_1682),
.B1(n_1690),
.B2(n_1685),
.C(n_1687),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1699),
.Y(n_1727)
);

NOR4xp25_ASAP7_75t_SL g1728 ( 
.A(n_1704),
.B(n_1688),
.C(n_1648),
.D(n_1684),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_SL g1729 ( 
.A(n_1697),
.B(n_1642),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1696),
.Y(n_1730)
);

OAI21xp33_ASAP7_75t_L g1731 ( 
.A1(n_1709),
.A2(n_1642),
.B(n_1688),
.Y(n_1731)
);

OAI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1729),
.A2(n_1697),
.B1(n_1702),
.B2(n_1693),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1717),
.B(n_1712),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1722),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1731),
.A2(n_1697),
.B(n_1709),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1715),
.B(n_1712),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1723),
.B(n_1702),
.Y(n_1737)
);

NAND4xp25_ASAP7_75t_L g1738 ( 
.A(n_1726),
.B(n_1707),
.C(n_1711),
.D(n_1702),
.Y(n_1738)
);

OAI31xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1725),
.A2(n_1706),
.A3(n_1708),
.B(n_1698),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1724),
.A2(n_1708),
.B1(n_1706),
.B2(n_1698),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1720),
.B(n_1701),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1721),
.A2(n_1727),
.B1(n_1720),
.B2(n_1719),
.Y(n_1742)
);

NOR4xp25_ASAP7_75t_SL g1743 ( 
.A(n_1728),
.B(n_1696),
.C(n_1710),
.D(n_1648),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1716),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1721),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1718),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1721),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1727),
.B(n_1701),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1730),
.B(n_1710),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_R g1750 ( 
.A(n_1729),
.B(n_71),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1726),
.A2(n_1686),
.B(n_74),
.C(n_71),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1720),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1737),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1733),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1734),
.B(n_1703),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1736),
.B(n_1703),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1746),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1750),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1738),
.B(n_73),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1752),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1751),
.A2(n_1686),
.B(n_1710),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1745),
.B(n_1660),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1739),
.B(n_1710),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1758),
.B(n_1735),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1754),
.B(n_1740),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1753),
.B(n_1745),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1760),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1759),
.B(n_1747),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1757),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1767),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1764),
.B(n_1763),
.Y(n_1771)
);

OAI21xp33_ASAP7_75t_L g1772 ( 
.A1(n_1764),
.A2(n_1742),
.B(n_1756),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1765),
.B(n_1755),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1770),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1771),
.B(n_1768),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1773),
.B(n_1749),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1772),
.B(n_1766),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1774),
.A2(n_1751),
.B(n_1761),
.C(n_1732),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1777),
.B(n_1769),
.Y(n_1779)
);

OAI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1775),
.A2(n_1747),
.B1(n_1761),
.B2(n_1762),
.C1(n_1755),
.C2(n_1744),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1776),
.B(n_1746),
.Y(n_1781)
);

A2O1A1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1775),
.A2(n_1746),
.B(n_1748),
.C(n_1741),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1777),
.B(n_1743),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1778),
.B(n_1779),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1781),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1782),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1783),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1780),
.B(n_77),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1781),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1779),
.A2(n_1660),
.B1(n_1703),
.B2(n_1694),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1779),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1779),
.Y(n_1792)
);

INVxp67_ASAP7_75t_L g1793 ( 
.A(n_1779),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1779),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1794),
.B(n_1743),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1786),
.A2(n_1694),
.B1(n_1637),
.B2(n_79),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1788),
.A2(n_1694),
.B1(n_1637),
.B2(n_79),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1784),
.A2(n_1694),
.B1(n_78),
.B2(n_80),
.C(n_81),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1794),
.A2(n_80),
.B1(n_77),
.B2(n_78),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_1793),
.B(n_82),
.C(n_84),
.Y(n_1800)
);

O2A1O1Ixp5_ASAP7_75t_L g1801 ( 
.A1(n_1787),
.A2(n_87),
.B(n_82),
.C(n_86),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1785),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1789),
.B(n_86),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1791),
.A2(n_87),
.B(n_89),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1792),
.B(n_89),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1790),
.B(n_90),
.Y(n_1806)
);

AOI211xp5_ASAP7_75t_L g1807 ( 
.A1(n_1788),
.A2(n_93),
.B(n_90),
.C(n_92),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1785),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1794),
.B(n_92),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1794),
.B(n_93),
.Y(n_1810)
);

NOR2x1_ASAP7_75t_L g1811 ( 
.A(n_1788),
.B(n_94),
.Y(n_1811)
);

AOI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1810),
.A2(n_1811),
.B(n_1803),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1809),
.Y(n_1813)
);

OAI21xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1802),
.A2(n_95),
.B(n_96),
.Y(n_1814)
);

AOI21xp33_ASAP7_75t_L g1815 ( 
.A1(n_1808),
.A2(n_1806),
.B(n_1807),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1801),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1799),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1797),
.B(n_97),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1795),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1798),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1805),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1800),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1804),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.C1(n_104),
.C2(n_105),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1796),
.A2(n_102),
.B(n_103),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1809),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1811),
.B(n_105),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1807),
.B(n_106),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1803),
.A2(n_106),
.B(n_107),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1818),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1819),
.B(n_107),
.C(n_108),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1814),
.B(n_108),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1813),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1817),
.B(n_110),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1826),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1824),
.B(n_110),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1822),
.B(n_111),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1827),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1825),
.B(n_428),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1823),
.B(n_119),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1822),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1820),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.C(n_124),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1821),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1828),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1816),
.B(n_1815),
.Y(n_1844)
);

NOR2xp67_ASAP7_75t_SL g1845 ( 
.A(n_1812),
.B(n_125),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1818),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1827),
.Y(n_1847)
);

OAI211xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1843),
.A2(n_1844),
.B(n_1846),
.C(n_1832),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1840),
.Y(n_1849)
);

OAI321xp33_ASAP7_75t_L g1850 ( 
.A1(n_1829),
.A2(n_130),
.A3(n_131),
.B1(n_132),
.B2(n_134),
.C(n_135),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1834),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1833),
.B(n_136),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1835),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1831),
.A2(n_141),
.B(n_138),
.C(n_139),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1842),
.Y(n_1855)
);

AOI322xp5_ASAP7_75t_L g1856 ( 
.A1(n_1847),
.A2(n_143),
.A3(n_146),
.B1(n_147),
.B2(n_148),
.C1(n_151),
.C2(n_152),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1830),
.A2(n_155),
.B1(n_156),
.B2(n_159),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1836),
.Y(n_1858)
);

OAI211xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1847),
.A2(n_161),
.B(n_162),
.C(n_163),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_L g1860 ( 
.A(n_1841),
.B(n_164),
.C(n_165),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1839),
.A2(n_166),
.B1(n_167),
.B2(n_170),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1838),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1849),
.B(n_1837),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1848),
.B(n_1845),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1851),
.B(n_172),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1855),
.B(n_1858),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1854),
.A2(n_173),
.B(n_175),
.C(n_176),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1858),
.Y(n_1868)
);

XOR2x1_ASAP7_75t_L g1869 ( 
.A(n_1852),
.B(n_179),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1862),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1853),
.Y(n_1871)
);

NOR4xp25_ASAP7_75t_L g1872 ( 
.A(n_1850),
.B(n_182),
.C(n_185),
.D(n_186),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1861),
.B(n_187),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1857),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1860),
.B(n_188),
.Y(n_1875)
);

NAND4xp25_ASAP7_75t_L g1876 ( 
.A(n_1859),
.B(n_189),
.C(n_190),
.D(n_193),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1863),
.A2(n_1856),
.B(n_196),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1875),
.A2(n_198),
.B1(n_200),
.B2(n_202),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1864),
.B(n_204),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1865),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1872),
.B(n_205),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1866),
.A2(n_425),
.B1(n_211),
.B2(n_212),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1868),
.Y(n_1883)
);

AND4x1_ASAP7_75t_L g1884 ( 
.A(n_1867),
.B(n_1870),
.C(n_1869),
.D(n_1876),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_SL g1885 ( 
.A(n_1874),
.B(n_208),
.C(n_213),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1883),
.B(n_1871),
.Y(n_1886)
);

AOI322xp5_ASAP7_75t_L g1887 ( 
.A1(n_1880),
.A2(n_1873),
.A3(n_218),
.B1(n_219),
.B2(n_220),
.C1(n_221),
.C2(n_222),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1881),
.A2(n_214),
.B1(n_223),
.B2(n_224),
.Y(n_1888)
);

OAI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1878),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.C(n_229),
.Y(n_1889)
);

AOI322xp5_ASAP7_75t_L g1890 ( 
.A1(n_1879),
.A2(n_232),
.A3(n_234),
.B1(n_236),
.B2(n_237),
.C1(n_238),
.C2(n_241),
.Y(n_1890)
);

AOI322xp5_ASAP7_75t_L g1891 ( 
.A1(n_1885),
.A2(n_242),
.A3(n_243),
.B1(n_246),
.B2(n_248),
.C1(n_250),
.C2(n_252),
.Y(n_1891)
);

OAI211xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1877),
.A2(n_254),
.B(n_255),
.C(n_256),
.Y(n_1892)
);

AOI322xp5_ASAP7_75t_L g1893 ( 
.A1(n_1884),
.A2(n_257),
.A3(n_258),
.B1(n_259),
.B2(n_260),
.C1(n_266),
.C2(n_268),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1886),
.Y(n_1894)
);

NOR4xp25_ASAP7_75t_SL g1895 ( 
.A(n_1892),
.B(n_1882),
.C(n_270),
.D(n_273),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1888),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1889),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1894),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1897),
.A2(n_1887),
.B1(n_1893),
.B2(n_1891),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1896),
.A2(n_1890),
.B1(n_275),
.B2(n_278),
.Y(n_1900)
);

AOI211x1_ASAP7_75t_L g1901 ( 
.A1(n_1895),
.A2(n_269),
.B(n_280),
.C(n_282),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1894),
.Y(n_1902)
);

OAI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1898),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1899),
.A2(n_297),
.B1(n_299),
.B2(n_301),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1900),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1901),
.Y(n_1907)
);

AOI21xp33_ASAP7_75t_L g1908 ( 
.A1(n_1904),
.A2(n_302),
.B(n_304),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1905),
.A2(n_306),
.B1(n_307),
.B2(n_310),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1906),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1910),
.A2(n_1907),
.B(n_1903),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1909),
.A2(n_312),
.B(n_314),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1908),
.A2(n_315),
.B(n_316),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1911),
.B(n_322),
.Y(n_1914)
);

AND2x2_ASAP7_75t_SL g1915 ( 
.A(n_1914),
.B(n_1912),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1913),
.B1(n_326),
.B2(n_328),
.Y(n_1916)
);

AOI211xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_323),
.B(n_329),
.C(n_331),
.Y(n_1917)
);


endmodule