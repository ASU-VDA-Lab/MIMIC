module fake_jpeg_25495_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_62),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

CKINVDCx11_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_47),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_48),
.C(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_19),
.B1(n_21),
.B2(n_28),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_51),
.B1(n_29),
.B2(n_34),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_19),
.B1(n_21),
.B2(n_28),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_82),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_26),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_89),
.B1(n_98),
.B2(n_59),
.Y(n_105)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_99),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_45),
.B1(n_49),
.B2(n_18),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_65),
.B1(n_52),
.B2(n_45),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_101),
.A2(n_104),
.B1(n_91),
.B2(n_87),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_65),
.B1(n_49),
.B2(n_52),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_92),
.B(n_99),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_48),
.C(n_47),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_119),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_70),
.B1(n_86),
.B2(n_85),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_36),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_35),
.B1(n_34),
.B2(n_23),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_70),
.B(n_86),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_121),
.B1(n_123),
.B2(n_127),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_130),
.B(n_55),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_73),
.B1(n_79),
.B2(n_94),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_132),
.B1(n_139),
.B2(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_93),
.B1(n_90),
.B2(n_86),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_143),
.Y(n_164)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_84),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_151),
.Y(n_167)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_141),
.Y(n_160)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_150),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_69),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_151),
.B(n_152),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_80),
.B1(n_90),
.B2(n_76),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_155),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_75),
.B1(n_76),
.B2(n_83),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_120),
.B1(n_108),
.B2(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_77),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_66),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_156),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_68),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_121),
.B1(n_117),
.B2(n_119),
.Y(n_158)
);

NAND2x1_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_163),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_162),
.B(n_166),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_118),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_118),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_172),
.B(n_180),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_183),
.B1(n_172),
.B2(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_134),
.B(n_153),
.C(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_190),
.B(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

O2A1O1Ixp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_102),
.B(n_109),
.C(n_36),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_102),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_95),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_95),
.B1(n_78),
.B2(n_48),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_191),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_192),
.B(n_193),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_193),
.B(n_218),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_170),
.B(n_162),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_194),
.A2(n_207),
.B(n_50),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_174),
.A2(n_157),
.B1(n_136),
.B2(n_140),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g242 ( 
.A1(n_197),
.A2(n_199),
.B(n_50),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_136),
.B(n_112),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_220),
.B(n_40),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_124),
.B1(n_137),
.B2(n_123),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_206),
.B1(n_212),
.B2(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_168),
.B1(n_158),
.B2(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_33),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_23),
.B1(n_35),
.B2(n_29),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_179),
.B1(n_184),
.B2(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_173),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_218)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_158),
.B(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_47),
.C(n_40),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_201),
.C(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_161),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_167),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_226),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_166),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_194),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_185),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_161),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_207),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_171),
.B1(n_17),
.B2(n_36),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_239),
.B1(n_205),
.B2(n_217),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_204),
.B1(n_220),
.B2(n_203),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_243),
.B1(n_216),
.B2(n_205),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_171),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_238),
.B(n_241),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_24),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_244),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_247),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_10),
.B(n_16),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_228),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_249),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_221),
.C(n_196),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.C(n_267),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_196),
.C(n_209),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_256),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_202),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_199),
.B(n_215),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_0),
.B(n_1),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_202),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_225),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_247),
.B1(n_232),
.B2(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_214),
.C(n_219),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_9),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_268),
.B(n_11),
.Y(n_284)
);

OA21x2_ASAP7_75t_SL g270 ( 
.A1(n_262),
.A2(n_240),
.B(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_273),
.B1(n_278),
.B2(n_276),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_245),
.B1(n_232),
.B2(n_227),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_280),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_227),
.B1(n_236),
.B2(n_239),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_279),
.A2(n_287),
.B1(n_257),
.B2(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_222),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_244),
.C(n_31),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_254),
.C(n_256),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_258),
.B(n_263),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_259),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_288),
.A2(n_303),
.B1(n_1),
.B2(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_302),
.C(n_12),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_264),
.C(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

AO221x1_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_248),
.B1(n_258),
.B2(n_269),
.C(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_298),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_253),
.C(n_269),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_274),
.C(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_8),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_300),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_9),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_50),
.C(n_9),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_272),
.B1(n_273),
.B2(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_7),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_7),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_50),
.B(n_2),
.C(n_3),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_3),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_310),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_12),
.CI(n_14),
.CON(n_311),
.SN(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_294),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_293),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_6),
.C(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_6),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_317),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_297),
.B(n_293),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_323),
.C(n_324),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_322),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_306),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_6),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_305),
.B(n_13),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_315),
.B1(n_313),
.B2(n_311),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_316),
.C(n_307),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.C(n_321),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_307),
.C(n_13),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_330),
.B1(n_326),
.B2(n_327),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_330),
.C(n_333),
.Y(n_338)
);

AOI321xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_4),
.A3(n_14),
.B1(n_16),
.B2(n_330),
.C(n_335),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_16),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_4),
.Y(n_342)
);


endmodule