module fake_jpeg_2206_n_211 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_211);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_60),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_64),
.Y(n_95)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_73),
.B1(n_64),
.B2(n_71),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_57),
.B1(n_54),
.B2(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_81),
.B1(n_53),
.B2(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_104),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_63),
.B1(n_71),
.B2(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_102),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_69),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_70),
.B1(n_59),
.B2(n_58),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_72),
.B1(n_62),
.B2(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_121),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_120),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_98),
.B1(n_106),
.B2(n_4),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_59),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_52),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_126),
.Y(n_143)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_1),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_120),
.B(n_123),
.C(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_146),
.B1(n_155),
.B2(n_8),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_2),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_106),
.B1(n_22),
.B2(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_19),
.B1(n_46),
.B2(n_45),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_3),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_116),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_49),
.B1(n_44),
.B2(n_42),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_41),
.B(n_40),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_37),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_170),
.C(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_5),
.B(n_6),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_155),
.B1(n_138),
.B2(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_9),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_35),
.C(n_34),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_31),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_30),
.B(n_28),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_174),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_144),
.B1(n_138),
.B2(n_11),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_27),
.B(n_10),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_185),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_161),
.B1(n_162),
.B2(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_167),
.B1(n_174),
.B2(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_10),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_158),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_179),
.B(n_180),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_11),
.B(n_12),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_163),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_171),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.C(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_170),
.C(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_198),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_186),
.A3(n_184),
.B1(n_178),
.B2(n_177),
.C1(n_15),
.C2(n_16),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_190),
.C(n_198),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_192),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_204),
.Y(n_206)
);

AOI211xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_201),
.B(n_205),
.C(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_13),
.C(n_14),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

OAI311xp33_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_18),
.A3(n_14),
.B1(n_15),
.C1(n_17),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_13),
.Y(n_211)
);


endmodule