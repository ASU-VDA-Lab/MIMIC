module fake_jpeg_1815_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_69),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_17),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_72),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_15),
.B(n_8),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_80),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_26),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_85),
.B(n_0),
.Y(n_121)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_16),
.B1(n_20),
.B2(n_42),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_88),
.A2(n_100),
.B1(n_105),
.B2(n_114),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_42),
.B1(n_20),
.B2(n_41),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_126),
.B1(n_74),
.B2(n_52),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_42),
.B1(n_20),
.B2(n_16),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_54),
.B1(n_83),
.B2(n_56),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_36),
.B1(n_24),
.B2(n_33),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_128),
.B1(n_51),
.B2(n_61),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_99),
.B(n_122),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_36),
.B1(n_32),
.B2(n_30),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_32),
.B1(n_28),
.B2(n_25),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_39),
.B1(n_35),
.B2(n_18),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_39),
.B1(n_35),
.B2(n_2),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_9),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_35),
.B1(n_39),
.B2(n_10),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_86),
.B1(n_82),
.B2(n_79),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_53),
.A2(n_39),
.B1(n_35),
.B2(n_3),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_75),
.A2(n_39),
.B1(n_35),
.B2(n_0),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_135),
.B1(n_1),
.B2(n_8),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_55),
.A2(n_39),
.B1(n_35),
.B2(n_0),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_140),
.Y(n_193)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g190 ( 
.A(n_139),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_49),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_179),
.Y(n_195)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_49),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_146),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_66),
.B1(n_64),
.B2(n_54),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_171),
.B1(n_118),
.B2(n_102),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_48),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_147),
.B(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_56),
.B(n_5),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_149),
.B(n_182),
.Y(n_216)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_91),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_163),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_169),
.B1(n_128),
.B2(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_5),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_170),
.Y(n_215)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_8),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_92),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_110),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_93),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_103),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_94),
.Y(n_197)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_103),
.B(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_142),
.A2(n_115),
.B1(n_108),
.B2(n_97),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_121),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_214),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_198),
.B1(n_155),
.B2(n_137),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_94),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_217),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_152),
.A2(n_127),
.B(n_118),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_201),
.A2(n_160),
.B(n_174),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_183),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_90),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_140),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_102),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_148),
.Y(n_229)
);

INVx2_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_224),
.B(n_198),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_151),
.A2(n_111),
.B(n_116),
.C(n_155),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_140),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_161),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_230),
.B(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_164),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_234),
.A2(n_238),
.B1(n_253),
.B2(n_190),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_235),
.A2(n_236),
.B(n_243),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_181),
.B(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_111),
.B1(n_116),
.B2(n_153),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_165),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_162),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_178),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_188),
.A2(n_143),
.B(n_150),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_178),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_246),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_251),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_154),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_193),
.A2(n_177),
.B1(n_178),
.B2(n_139),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_193),
.C(n_200),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_246),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_282),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_193),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_262),
.B(n_282),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_225),
.A2(n_195),
.B1(n_224),
.B2(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_280),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_195),
.B(n_186),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_267),
.A2(n_272),
.B(n_277),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_223),
.B(n_222),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_204),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_284),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_222),
.B(n_204),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_232),
.B(n_257),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_226),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_213),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_194),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_194),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_237),
.Y(n_303)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_244),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_190),
.Y(n_295)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_184),
.C(n_208),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_235),
.C(n_250),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_296),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_228),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_236),
.B(n_243),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_297),
.B(n_300),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_227),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_302),
.C(n_309),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_258),
.C(n_231),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_306),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_291),
.Y(n_306)
);

XOR2x2_ASAP7_75t_SL g307 ( 
.A(n_287),
.B(n_257),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_313),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_310),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_256),
.C(n_255),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_238),
.B(n_249),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_270),
.A2(n_248),
.B(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_247),
.Y(n_315)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_315),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_244),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_316),
.Y(n_323)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_267),
.B1(n_277),
.B2(n_283),
.Y(n_322)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_315),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_327),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_292),
.C(n_279),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_330),
.C(n_338),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_295),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_298),
.B(n_265),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_331),
.C(n_337),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_269),
.C(n_280),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_271),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_271),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_263),
.C(n_272),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_299),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_330),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_311),
.A2(n_286),
.B1(n_272),
.B2(n_290),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_340),
.A2(n_311),
.B1(n_310),
.B2(n_304),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_312),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_309),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_294),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_344),
.Y(n_368)
);

BUFx12_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_328),
.B(n_318),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_352),
.Y(n_365)
);

NOR3xp33_ASAP7_75t_SL g346 ( 
.A(n_332),
.B(n_312),
.C(n_317),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_346),
.B(n_350),
.Y(n_370)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_321),
.B(n_264),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_313),
.Y(n_352)
);

BUFx12_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_353),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_358),
.Y(n_363)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_326),
.A2(n_300),
.B(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_320),
.A2(n_316),
.B1(n_268),
.B2(n_266),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g359 ( 
.A1(n_331),
.A2(n_307),
.B(n_268),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_359),
.A2(n_341),
.B(n_335),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_364),
.A2(n_345),
.B(n_353),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_360),
.Y(n_366)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_321),
.C(n_336),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_373),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_338),
.C(n_335),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_342),
.C(n_349),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_376),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_348),
.C(n_337),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_348),
.Y(n_377)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_377),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_364),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_383),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_366),
.A2(n_323),
.B1(n_346),
.B2(n_333),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_385),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_365),
.Y(n_391)
);

XOR2x2_ASAP7_75t_SL g383 ( 
.A(n_363),
.B(n_353),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_266),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g388 ( 
.A(n_377),
.B(n_363),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_394),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_382),
.A2(n_375),
.B(n_373),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_390),
.A2(n_391),
.B(n_389),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_396),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_371),
.C(n_383),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_362),
.C(n_376),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_399),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_367),
.Y(n_399)
);

A2O1A1O1Ixp25_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_378),
.B(n_343),
.C(n_369),
.D(n_372),
.Y(n_400)
);

A2O1A1Ixp33_ASAP7_75t_L g405 ( 
.A1(n_400),
.A2(n_401),
.B(n_273),
.C(n_289),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_369),
.Y(n_401)
);

AOI322xp5_ASAP7_75t_L g403 ( 
.A1(n_397),
.A2(n_343),
.A3(n_393),
.B1(n_289),
.B2(n_273),
.C1(n_288),
.C2(n_203),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_403),
.A2(n_405),
.B(n_401),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_406),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_288),
.B(n_190),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_402),
.B(n_407),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_208),
.Y(n_410)
);


endmodule