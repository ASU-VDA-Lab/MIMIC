module fake_netlist_5_1362_n_1685 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1685);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1685;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_35),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_35),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_84),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_45),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_85),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_61),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_16),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_54),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_56),
.Y(n_165)
);

BUFx8_ASAP7_75t_SL g166 ( 
.A(n_3),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_37),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_33),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_80),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_115),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_12),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_95),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_68),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_112),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_69),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_20),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_7),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_98),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_36),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_113),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_75),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_78),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_109),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_52),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_33),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_62),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_7),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_141),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_106),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_5),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_71),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_1),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_42),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_65),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_39),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_31),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_139),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_17),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_47),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_6),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_51),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_67),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_128),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_140),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_104),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_79),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_101),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

HB1xp67_ASAP7_75t_SL g245 ( 
.A(n_40),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_81),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_29),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_24),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_70),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_57),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_137),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_31),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_93),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_108),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_0),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_25),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_48),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_1),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_38),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_45),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_138),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_26),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_11),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_44),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_100),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_19),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_15),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_146),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_114),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_29),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_131),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_77),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_124),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_24),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_13),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_74),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_30),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_20),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_88),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_53),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_25),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_90),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_39),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_166),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_174),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_160),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_160),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_176),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_174),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_174),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_256),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_174),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_166),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_219),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_225),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_204),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_175),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_175),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_154),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_219),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_219),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_230),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_176),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_183),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_185),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_168),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_181),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_193),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_208),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_245),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_217),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_254),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_202),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_213),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_230),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_176),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_163),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_157),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_157),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_191),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_242),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_196),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_215),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_260),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_197),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_197),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_207),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_196),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_203),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_203),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_159),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_195),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_221),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_234),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_224),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_207),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_274),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_164),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_170),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_163),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_195),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_367),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_324),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_311),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_231),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_306),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_231),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_195),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_169),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_329),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_308),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_324),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_167),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_374),
.B(n_370),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_315),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_331),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_180),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_178),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_318),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_319),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_312),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_330),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_310),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_331),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_178),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_189),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_322),
.A2(n_209),
.B1(n_223),
.B2(n_264),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_334),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_307),
.B(n_189),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_323),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_357),
.A2(n_210),
.B(n_192),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_327),
.A2(n_278),
.B1(n_153),
.B2(n_209),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_309),
.B(n_210),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_334),
.B(n_184),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_353),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_377),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_336),
.B(n_167),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_378),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_321),
.A2(n_328),
.B1(n_381),
.B2(n_355),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_341),
.B(n_222),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_340),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_339),
.B(n_194),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_337),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_407),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_419),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_384),
.B(n_392),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_385),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_453),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_339),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_399),
.B(n_346),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g469 ( 
.A(n_396),
.B(n_255),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_346),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_453),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_404),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_423),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_406),
.B(n_342),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g480 ( 
.A1(n_450),
.A2(n_274),
.B1(n_297),
.B2(n_188),
.Y(n_480)
);

NOR2x1p5_ASAP7_75t_L g481 ( 
.A(n_405),
.B(n_305),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_398),
.B(n_328),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

AO22x2_ASAP7_75t_L g487 ( 
.A1(n_397),
.A2(n_227),
.B1(n_257),
.B2(n_198),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_413),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_406),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_410),
.B(n_349),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_427),
.A2(n_351),
.B1(n_347),
.B2(n_343),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_437),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_413),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_415),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_438),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_389),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_425),
.B(n_349),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_393),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_444),
.B(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_414),
.B(n_395),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_448),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_394),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_455),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_433),
.B(n_345),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_440),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_448),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_427),
.A2(n_363),
.B1(n_350),
.B2(n_352),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_429),
.B(n_271),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_414),
.B(n_373),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_417),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_SL g526 ( 
.A(n_451),
.B(n_255),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_425),
.A2(n_373),
.B1(n_375),
.B2(n_266),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_425),
.B(n_375),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_424),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_408),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_414),
.B(n_237),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_393),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_394),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_425),
.B(n_305),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_425),
.B(n_316),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_414),
.B(n_286),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_427),
.A2(n_368),
.B1(n_348),
.B2(n_271),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_425),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_420),
.B(n_155),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_400),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_400),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_400),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_422),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_401),
.Y(n_554)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_411),
.A2(n_229),
.B(n_200),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_386),
.B(n_156),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_394),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_394),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_431),
.B(n_316),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_433),
.B(n_241),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_401),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_401),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_441),
.A2(n_294),
.B1(n_282),
.B2(n_284),
.Y(n_565)
);

BUFx6f_ASAP7_75t_SL g566 ( 
.A(n_433),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_426),
.B(n_442),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_432),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_432),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_432),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_441),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_443),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_443),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_427),
.B(n_344),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_443),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_446),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_433),
.B(n_271),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_386),
.B(n_158),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_434),
.B(n_232),
.C(n_228),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_394),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_L g586 ( 
.A(n_383),
.B(n_176),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_402),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_446),
.Y(n_588)
);

INVx6_ASAP7_75t_L g589 ( 
.A(n_402),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_402),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_402),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_435),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_402),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_428),
.B(n_290),
.C(n_268),
.Y(n_594)
);

INVx8_ASAP7_75t_L g595 ( 
.A(n_383),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_446),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_402),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_387),
.B(n_161),
.Y(n_598)
);

NOR2x1p5_ASAP7_75t_L g599 ( 
.A(n_434),
.B(n_244),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_567),
.B(n_435),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_489),
.B(n_435),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_489),
.B(n_435),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_483),
.B(n_492),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_512),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_544),
.B(n_449),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_508),
.B(n_338),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_471),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_592),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_462),
.A2(n_452),
.B(n_447),
.C(n_439),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_504),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_510),
.A2(n_281),
.B1(n_243),
.B2(n_246),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_459),
.B(n_358),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_502),
.B(n_449),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_518),
.B(n_465),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_502),
.B(n_449),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_599),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_479),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_592),
.B(n_449),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_474),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_491),
.B(n_364),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_510),
.B(n_520),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_507),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_466),
.B(n_365),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_520),
.B(n_446),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_L g629 ( 
.A1(n_491),
.A2(n_280),
.B1(n_265),
.B2(n_376),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_507),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_522),
.B(n_468),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_471),
.B(n_446),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_507),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_460),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_472),
.A2(n_387),
.B(n_388),
.Y(n_635)
);

BUFx8_ASAP7_75t_L g636 ( 
.A(n_457),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_523),
.B(n_176),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_461),
.Y(n_638)
);

NAND2x1_ASAP7_75t_L g639 ( 
.A(n_471),
.B(n_383),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_514),
.B(n_446),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_457),
.B(n_428),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_469),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_514),
.B(n_412),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_518),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_463),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_479),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_522),
.B(n_366),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_500),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_529),
.B(n_265),
.Y(n_649)
);

AND2x6_ASAP7_75t_SL g650 ( 
.A(n_562),
.B(n_153),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_527),
.B(n_412),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_469),
.B(n_280),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_527),
.B(n_412),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_532),
.B(n_163),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_505),
.B(n_239),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_482),
.B(n_388),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_516),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_480),
.A2(n_487),
.B1(n_536),
.B2(n_531),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_526),
.A2(n_211),
.B1(n_171),
.B2(n_165),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_539),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_482),
.B(n_388),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_476),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_530),
.B(n_239),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_541),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_486),
.B(n_490),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_595),
.Y(n_667)
);

NOR2xp67_ASAP7_75t_L g668 ( 
.A(n_463),
.B(n_436),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_541),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_486),
.B(n_412),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_562),
.B(n_452),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_556),
.A2(n_416),
.B(n_412),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_549),
.B(n_304),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_584),
.B(n_304),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_548),
.B(n_176),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_569),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_566),
.A2(n_205),
.B1(n_162),
.B2(n_302),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_573),
.B(n_287),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_498),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_490),
.B(n_412),
.Y(n_683)
);

NOR2x1p5_ASAP7_75t_L g684 ( 
.A(n_533),
.B(n_249),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_571),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_562),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_586),
.A2(n_447),
.B(n_439),
.C(n_436),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_498),
.Y(n_688)
);

NAND2x1p5_ASAP7_75t_L g689 ( 
.A(n_548),
.B(n_250),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_566),
.A2(n_190),
.B1(n_172),
.B2(n_173),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_571),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_493),
.B(n_416),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_572),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_538),
.B(n_177),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_566),
.A2(n_201),
.B1(n_179),
.B2(n_182),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_550),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_572),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_493),
.B(n_416),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_550),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_574),
.B(n_458),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_546),
.B(n_186),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_565),
.B(n_187),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_545),
.B(n_533),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_590),
.B(n_261),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_467),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_477),
.B(n_258),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_532),
.B(n_199),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_495),
.B(n_416),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_495),
.B(n_416),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_467),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_496),
.B(n_416),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_574),
.A2(n_562),
.B1(n_285),
.B2(n_277),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_496),
.B(n_176),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_595),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_238),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_551),
.B(n_238),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_532),
.B(n_206),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_470),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_552),
.B(n_238),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_595),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_515),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_470),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_552),
.B(n_238),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_583),
.B(n_269),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_475),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_475),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_554),
.B(n_238),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_547),
.B(n_212),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_554),
.A2(n_214),
.B(n_216),
.C(n_235),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_598),
.B(n_594),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_480),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_550),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_480),
.A2(n_238),
.B1(n_287),
.B2(n_383),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_590),
.B(n_473),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_595),
.Y(n_735)
);

BUFx5_ASAP7_75t_L g736 ( 
.A(n_563),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_573),
.A2(n_430),
.B(n_287),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_563),
.B(n_238),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_480),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_458),
.B(n_296),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_557),
.B(n_296),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_564),
.B(n_383),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_487),
.A2(n_481),
.B1(n_582),
.B2(n_292),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_557),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_487),
.A2(n_223),
.B1(n_264),
.B2(n_278),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_590),
.B(n_383),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_485),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_487),
.B(n_296),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_586),
.B(n_303),
.C(n_273),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_494),
.B(n_218),
.Y(n_750)
);

INVx5_ASAP7_75t_L g751 ( 
.A(n_456),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_488),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_488),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_585),
.B(n_300),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_521),
.B(n_299),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_575),
.B(n_259),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_676),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_604),
.B(n_576),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_607),
.B(n_275),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_739),
.A2(n_582),
.B1(n_499),
.B2(n_501),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_679),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_685),
.Y(n_762)
);

AND2x4_ASAP7_75t_SL g763 ( 
.A(n_619),
.B(n_519),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_620),
.B(n_576),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_608),
.B(n_577),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_646),
.B(n_577),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_691),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_618),
.B(n_464),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_663),
.Y(n_769)
);

AOI21x1_ASAP7_75t_L g770 ( 
.A1(n_606),
.A2(n_597),
.B(n_587),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_609),
.Y(n_771)
);

INVx6_ASAP7_75t_L g772 ( 
.A(n_636),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_731),
.A2(n_582),
.B1(n_499),
.B2(n_501),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_688),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_624),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_693),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_721),
.B(n_519),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_675),
.B(n_478),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_697),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_631),
.A2(n_730),
.B1(n_627),
.B2(n_642),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_601),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_724),
.A2(n_591),
.B1(n_593),
.B2(n_596),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_667),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_600),
.B(n_478),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_682),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_648),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_608),
.B(n_579),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_654),
.Y(n_788)
);

AND2x2_ASAP7_75t_SL g789 ( 
.A(n_733),
.B(n_580),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_753),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_667),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_740),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_741),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_705),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_621),
.B(n_497),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_710),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_614),
.B(n_291),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_625),
.B(n_497),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_609),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_609),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_657),
.B(n_497),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_722),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_660),
.B(n_503),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_645),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_725),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_726),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_605),
.B(n_668),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_623),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_644),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_672),
.A2(n_580),
.B1(n_588),
.B2(n_581),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_747),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_752),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_616),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_602),
.A2(n_581),
.B1(n_226),
.B2(n_252),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_671),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_616),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_638),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_744),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_700),
.Y(n_821)
);

BUFx8_ASAP7_75t_L g822 ( 
.A(n_647),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_666),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_671),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_666),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_745),
.A2(n_582),
.B1(n_517),
.B2(n_524),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_665),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_628),
.B(n_503),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_745),
.A2(n_582),
.B1(n_517),
.B2(n_524),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_652),
.B(n_473),
.Y(n_830)
);

BUFx12f_ASAP7_75t_SL g831 ( 
.A(n_641),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_636),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_706),
.B(n_748),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_686),
.B(n_473),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_714),
.B(n_456),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_665),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_656),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_749),
.B(n_714),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_649),
.A2(n_582),
.B1(n_525),
.B2(n_528),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_703),
.A2(n_589),
.B1(n_233),
.B2(n_240),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_658),
.A2(n_525),
.B(n_553),
.C(n_542),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_714),
.B(n_456),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_SL g843 ( 
.A(n_629),
.B(n_262),
.C(n_247),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_656),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_602),
.Y(n_845)
);

AO22x1_ASAP7_75t_L g846 ( 
.A1(n_655),
.A2(n_289),
.B1(n_267),
.B2(n_253),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_661),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_720),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_687),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_603),
.B(n_615),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_SL g851 ( 
.A(n_702),
.B(n_251),
.C(n_293),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_736),
.Y(n_852)
);

NOR2x1p5_ASAP7_75t_L g853 ( 
.A(n_650),
.B(n_298),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_603),
.B(n_528),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_736),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_622),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_641),
.B(n_555),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_615),
.A2(n_540),
.B1(n_534),
.B2(n_535),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_736),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_SL g860 ( 
.A(n_677),
.B(n_222),
.C(n_4),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_617),
.B(n_540),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_611),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_720),
.B(n_484),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_735),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_712),
.B(n_570),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_612),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_617),
.B(n_537),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_626),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_735),
.B(n_684),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_630),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_707),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_735),
.B(n_484),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_664),
.A2(n_589),
.B1(n_570),
.B2(n_568),
.Y(n_873)
);

AND2x6_ASAP7_75t_SL g874 ( 
.A(n_641),
.B(n_222),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_633),
.Y(n_875)
);

NOR2x1p5_ASAP7_75t_L g876 ( 
.A(n_756),
.B(n_542),
.Y(n_876)
);

BUFx4f_ASAP7_75t_L g877 ( 
.A(n_689),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_736),
.B(n_456),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_734),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_756),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_640),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_610),
.B(n_537),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_717),
.B(n_534),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_736),
.B(n_456),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_743),
.B(n_513),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_674),
.B(n_570),
.Y(n_886)
);

AND2x4_ASAP7_75t_SL g887 ( 
.A(n_659),
.B(n_484),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_750),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_662),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_637),
.A2(n_589),
.B1(n_568),
.B2(n_513),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_SL g891 ( 
.A1(n_689),
.A2(n_0),
.B1(n_10),
.B2(n_11),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_680),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_643),
.A2(n_560),
.B(n_535),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_690),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_694),
.B(n_701),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_734),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_755),
.B(n_568),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_651),
.B(n_484),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_669),
.Y(n_899)
);

BUFx12f_ASAP7_75t_L g900 ( 
.A(n_704),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_653),
.B(n_560),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_754),
.B(n_553),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_696),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_699),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_732),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_728),
.A2(n_559),
.B1(n_558),
.B2(n_543),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_613),
.B(n_484),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_670),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_632),
.B(n_559),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_695),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_670),
.B(n_559),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_683),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_683),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_692),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_692),
.B(n_559),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_742),
.B(n_751),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_R g917 ( 
.A(n_678),
.B(n_76),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_698),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_713),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_698),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_708),
.B(n_559),
.Y(n_921)
);

BUFx4f_ASAP7_75t_SL g922 ( 
.A(n_681),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_729),
.A2(n_746),
.B1(n_639),
.B2(n_742),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_708),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_709),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_709),
.B(n_558),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_713),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_711),
.B(n_558),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_751),
.B(n_543),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_711),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_751),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_715),
.B(n_558),
.C(n_543),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_715),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_791),
.B(n_864),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_823),
.A2(n_825),
.B1(n_780),
.B2(n_773),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_757),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_850),
.A2(n_635),
.B(n_673),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_SL g938 ( 
.A(n_759),
.B(n_833),
.C(n_894),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_845),
.B(n_704),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_818),
.B(n_719),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_931),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_779),
.Y(n_942)
);

BUFx8_ASAP7_75t_L g943 ( 
.A(n_775),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_881),
.A2(n_506),
.B(n_511),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_841),
.A2(n_719),
.B(n_738),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_781),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_781),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_797),
.B(n_716),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_895),
.A2(n_738),
.B(n_716),
.C(n_727),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_802),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_881),
.A2(n_506),
.B(n_511),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_879),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_815),
.B(n_723),
.Y(n_953)
);

AO21x2_ASAP7_75t_L g954 ( 
.A1(n_882),
.A2(n_758),
.B(n_932),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_845),
.B(n_558),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_773),
.A2(n_543),
.B1(n_737),
.B2(n_13),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_786),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_808),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_909),
.A2(n_681),
.B(n_59),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_792),
.B(n_10),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_802),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_841),
.A2(n_927),
.B(n_861),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_933),
.B(n_681),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_810),
.B(n_14),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_880),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_933),
.B(n_681),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_821),
.B(n_92),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_772),
.B(n_91),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_803),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_927),
.B(n_19),
.Y(n_970)
);

AO21x1_ASAP7_75t_L g971 ( 
.A1(n_830),
.A2(n_22),
.B(n_23),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_783),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_769),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_821),
.B(n_97),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_839),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_783),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_809),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_837),
.B(n_27),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_810),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.C(n_38),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_785),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_805),
.B(n_32),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_SL g982 ( 
.A(n_843),
.B(n_41),
.C(n_43),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_803),
.Y(n_983)
);

OR2x6_ASAP7_75t_L g984 ( 
.A(n_772),
.B(n_50),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_793),
.B(n_73),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_877),
.B(n_96),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_931),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_785),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_818),
.B(n_102),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_770),
.A2(n_105),
.B(n_116),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_854),
.A2(n_150),
.B(n_120),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_761),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_879),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_871),
.B(n_117),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_824),
.B(n_122),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_795),
.A2(n_134),
.B(n_147),
.C(n_148),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_769),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_839),
.A2(n_760),
.B1(n_847),
.B2(n_844),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_783),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_762),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_789),
.A2(n_849),
.B1(n_844),
.B2(n_847),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_832),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_912),
.B(n_914),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_774),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_830),
.A2(n_865),
.B(n_888),
.C(n_886),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_791),
.A2(n_864),
.B(n_878),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_791),
.A2(n_864),
.B(n_878),
.Y(n_1007)
);

CKINVDCx16_ASAP7_75t_R g1008 ( 
.A(n_777),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_767),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_776),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_893),
.A2(n_867),
.B(n_787),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_879),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_820),
.B(n_788),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_864),
.A2(n_884),
.B(n_901),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_817),
.B(n_892),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_931),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_843),
.A2(n_768),
.B(n_860),
.C(n_814),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_777),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_910),
.B(n_819),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_806),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_865),
.A2(n_886),
.B(n_919),
.C(n_877),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_L g1022 ( 
.A(n_840),
.B(n_869),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_831),
.B(n_900),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_920),
.B(n_925),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_930),
.B(n_908),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_789),
.A2(n_859),
.B1(n_855),
.B2(n_852),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_869),
.B(n_903),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_764),
.B(n_766),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_806),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_851),
.B(n_860),
.C(n_891),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_879),
.B(n_764),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_SL g1032 ( 
.A1(n_916),
.A2(n_835),
.B(n_872),
.C(n_863),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_908),
.B(n_913),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_857),
.A2(n_856),
.B(n_811),
.C(n_904),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_913),
.B(n_918),
.Y(n_1035)
);

OR2x6_ASAP7_75t_SL g1036 ( 
.A(n_816),
.B(n_794),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_883),
.A2(n_851),
.B(n_876),
.C(n_885),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_918),
.B(n_924),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_766),
.B(n_771),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_924),
.B(n_771),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_874),
.B(n_853),
.C(n_875),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_915),
.A2(n_928),
.B(n_921),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_777),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_826),
.A2(n_829),
.B1(n_891),
.B2(n_907),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_807),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_799),
.B(n_800),
.Y(n_1046)
);

AO22x1_ASAP7_75t_L g1047 ( 
.A1(n_822),
.A2(n_885),
.B1(n_838),
.B2(n_834),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_826),
.A2(n_829),
.B1(n_857),
.B2(n_858),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_765),
.A2(n_898),
.B(n_916),
.Y(n_1049)
);

INVx3_ASAP7_75t_SL g1050 ( 
.A(n_772),
.Y(n_1050)
);

CKINVDCx14_ASAP7_75t_R g1051 ( 
.A(n_857),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_838),
.B(n_848),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_799),
.B(n_800),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_904),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_902),
.B(n_798),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_796),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_783),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_905),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_763),
.B(n_813),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_887),
.A2(n_911),
.B(n_897),
.C(n_923),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_812),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_822),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_SL g1063 ( 
.A(n_917),
.B(n_782),
.C(n_873),
.Y(n_1063)
);

NOR2x1_ASAP7_75t_SL g1064 ( 
.A(n_848),
.B(n_931),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_887),
.A2(n_911),
.B(n_897),
.C(n_889),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_868),
.B(n_929),
.C(n_801),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_827),
.B(n_836),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_834),
.B(n_784),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_905),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_848),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1019),
.B(n_763),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_941),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_1060),
.A2(n_926),
.A3(n_828),
.B(n_778),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_1049),
.A2(n_765),
.B(n_858),
.Y(n_1074)
);

INVx8_ASAP7_75t_L g1075 ( 
.A(n_941),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_942),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_946),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_979),
.A2(n_846),
.B1(n_917),
.B2(n_804),
.C(n_790),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_950),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1003),
.B(n_1024),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_1005),
.A2(n_866),
.A3(n_870),
.B(n_862),
.Y(n_1081)
);

NAND2xp33_ASAP7_75t_L g1082 ( 
.A(n_1021),
.B(n_848),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1055),
.A2(n_842),
.B(n_835),
.Y(n_1083)
);

INVx3_ASAP7_75t_SL g1084 ( 
.A(n_1050),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1011),
.A2(n_1014),
.B(n_951),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1025),
.B(n_896),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1065),
.A2(n_1048),
.B(n_935),
.Y(n_1087)
);

OAI22x1_ASAP7_75t_L g1088 ( 
.A1(n_1030),
.A2(n_906),
.B1(n_899),
.B2(n_929),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_948),
.B(n_899),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_981),
.B(n_890),
.C(n_922),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_944),
.A2(n_945),
.B(n_990),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_945),
.A2(n_962),
.B(n_991),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1027),
.B(n_1052),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_962),
.A2(n_1044),
.B(n_935),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_961),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1033),
.B(n_1035),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1038),
.B(n_1001),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1006),
.A2(n_1007),
.B(n_1026),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_973),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_938),
.A2(n_1022),
.B1(n_1015),
.B2(n_958),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_943),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1044),
.A2(n_1034),
.B(n_998),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_941),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_977),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_998),
.A2(n_1063),
.B(n_1037),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1017),
.A2(n_956),
.B(n_978),
.Y(n_1106)
);

OA21x2_ASAP7_75t_L g1107 ( 
.A1(n_1066),
.A2(n_953),
.B(n_1068),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_955),
.A2(n_1040),
.B(n_1045),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_969),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_994),
.A2(n_1059),
.B1(n_1043),
.B2(n_1051),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_946),
.B(n_947),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1032),
.A2(n_954),
.B(n_939),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_971),
.A2(n_956),
.A3(n_975),
.B(n_965),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_985),
.A2(n_974),
.B1(n_967),
.B2(n_1018),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_940),
.B(n_936),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1052),
.B(n_989),
.Y(n_1116)
);

BUFx4f_ASAP7_75t_SL g1117 ( 
.A(n_947),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_964),
.B(n_970),
.C(n_975),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_997),
.B(n_1004),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1028),
.B(n_1054),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_983),
.A2(n_1029),
.B(n_1020),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1058),
.A2(n_1069),
.B(n_959),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_954),
.A2(n_1031),
.B(n_934),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_988),
.Y(n_1124)
);

OA21x2_ASAP7_75t_L g1125 ( 
.A1(n_963),
.A2(n_966),
.B(n_1056),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_960),
.B(n_995),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1053),
.A2(n_993),
.B(n_1012),
.Y(n_1127)
);

O2A1O1Ixp5_ASAP7_75t_L g1128 ( 
.A1(n_1047),
.A2(n_986),
.B(n_1039),
.C(n_940),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_943),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_SL g1130 ( 
.A1(n_1064),
.A2(n_934),
.B(n_989),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_996),
.A2(n_1061),
.B(n_1009),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_992),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1000),
.B(n_1010),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_952),
.A2(n_1012),
.B(n_993),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_972),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1008),
.B(n_1013),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_1002),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1067),
.Y(n_1138)
);

OA21x2_ASAP7_75t_L g1139 ( 
.A1(n_1036),
.A2(n_1041),
.B(n_982),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1057),
.A2(n_1046),
.A3(n_1016),
.B(n_987),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1057),
.A2(n_1016),
.A3(n_987),
.B(n_976),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1062),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_968),
.A2(n_984),
.B(n_976),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_968),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_968),
.B(n_984),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_999),
.A2(n_1070),
.B(n_984),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_999),
.A2(n_1070),
.B(n_1023),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_957),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1019),
.B(n_607),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1027),
.B(n_818),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1060),
.A2(n_608),
.B(n_937),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_973),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_957),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_SL g1154 ( 
.A1(n_1021),
.A2(n_1037),
.B(n_1005),
.C(n_1065),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1019),
.B(n_604),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_948),
.A2(n_604),
.B(n_759),
.C(n_780),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_943),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1003),
.B(n_823),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_938),
.B(n_721),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1060),
.A2(n_949),
.B(n_1005),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_946),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_980),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1060),
.A2(n_1005),
.A3(n_1048),
.B(n_1044),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1060),
.A2(n_608),
.B(n_1042),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1019),
.B(n_607),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_942),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1027),
.B(n_818),
.Y(n_1174)
);

INVx6_ASAP7_75t_SL g1175 ( 
.A(n_968),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_957),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_980),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1003),
.B(n_823),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_979),
.A2(n_604),
.B1(n_483),
.B2(n_745),
.C(n_607),
.Y(n_1179)
);

AO21x2_ASAP7_75t_L g1180 ( 
.A1(n_1060),
.A2(n_1005),
.B(n_1063),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_948),
.A2(n_604),
.B(n_759),
.C(n_780),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1003),
.B(n_823),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_957),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1002),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1003),
.B(n_823),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_938),
.A2(n_604),
.B1(n_607),
.B2(n_483),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1060),
.A2(n_1005),
.A3(n_1048),
.B(n_1044),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1002),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1060),
.A2(n_949),
.B(n_1005),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1060),
.A2(n_949),
.B(n_1005),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_988),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1027),
.B(n_818),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1060),
.A2(n_608),
.B(n_1042),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1049),
.A2(n_937),
.B(n_770),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_941),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1060),
.A2(n_608),
.B(n_1042),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_941),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_988),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1060),
.A2(n_608),
.B(n_937),
.Y(n_1202)
);

AOI221x1_ASAP7_75t_L g1203 ( 
.A1(n_1030),
.A2(n_604),
.B1(n_1044),
.B2(n_1005),
.C(n_1048),
.Y(n_1203)
);

AO21x2_ASAP7_75t_L g1204 ( 
.A1(n_1151),
.A2(n_1202),
.B(n_1112),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1156),
.B(n_1149),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1117),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1077),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1179),
.A2(n_1188),
.B1(n_1169),
.B2(n_1071),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1080),
.A2(n_1100),
.B1(n_1184),
.B2(n_1178),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1165),
.A2(n_1171),
.B(n_1170),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1166),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1133),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1133),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1080),
.B(n_1161),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1161),
.B(n_1178),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1172),
.A2(n_1183),
.B(n_1181),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1190),
.A2(n_1197),
.B(n_1085),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1202),
.A2(n_1168),
.B(n_1196),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1075),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1199),
.A2(n_1091),
.B(n_1098),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_SL g1221 ( 
.A1(n_1106),
.A2(n_1143),
.B(n_1105),
.Y(n_1221)
);

AND2x2_ASAP7_75t_SL g1222 ( 
.A(n_1092),
.B(n_1145),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1118),
.B(n_1114),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1074),
.A2(n_1122),
.B(n_1127),
.Y(n_1224)
);

OAI211xp5_ASAP7_75t_L g1225 ( 
.A1(n_1203),
.A2(n_1162),
.B(n_1087),
.C(n_1193),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1177),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1075),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1145),
.B(n_1146),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1163),
.A2(n_1192),
.B(n_1108),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1163),
.A2(n_1192),
.B(n_1123),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1083),
.A2(n_1102),
.B(n_1094),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1184),
.A2(n_1187),
.B1(n_1110),
.B2(n_1138),
.Y(n_1232)
);

CKINVDCx8_ASAP7_75t_R g1233 ( 
.A(n_1186),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1077),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1102),
.A2(n_1189),
.A3(n_1167),
.B1(n_1092),
.B2(n_1113),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_1078),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1126),
.B(n_1120),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1134),
.A2(n_1125),
.B(n_1097),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1130),
.B(n_1116),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1099),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1125),
.A2(n_1097),
.B(n_1086),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1187),
.A2(n_1082),
.B(n_1154),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1180),
.A2(n_1139),
.B1(n_1175),
.B2(n_1090),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1107),
.A2(n_1089),
.B(n_1115),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1136),
.A2(n_1093),
.B1(n_1195),
.B2(n_1150),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1084),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1075),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1081),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1115),
.A2(n_1096),
.B(n_1147),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1175),
.A2(n_1176),
.B1(n_1153),
.B2(n_1185),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1164),
.A2(n_1119),
.B1(n_1132),
.B2(n_1148),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1104),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1137),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1076),
.A2(n_1109),
.B(n_1173),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1079),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1095),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1081),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1194),
.B(n_1201),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1073),
.A2(n_1189),
.B(n_1167),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1124),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1073),
.A2(n_1167),
.B(n_1189),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1141),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1072),
.A2(n_1200),
.B(n_1198),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1174),
.B(n_1195),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1174),
.A2(n_1072),
.B(n_1198),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1159),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1103),
.A2(n_1200),
.B(n_1113),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1103),
.A2(n_1141),
.B(n_1140),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1101),
.A2(n_1129),
.B(n_1152),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1142),
.A2(n_1191),
.B1(n_1135),
.B2(n_1144),
.Y(n_1270)
);

AND2x2_ASAP7_75t_SL g1271 ( 
.A(n_1144),
.B(n_1135),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1158),
.A2(n_604),
.B(n_1182),
.C(n_483),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1192),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1133),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1145),
.B(n_1146),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1156),
.B(n_604),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1179),
.A2(n_604),
.B1(n_483),
.B2(n_1156),
.C(n_492),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1156),
.B(n_1149),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1077),
.B(n_1164),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1156),
.A2(n_604),
.B1(n_1188),
.B2(n_1182),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1077),
.B(n_1164),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1155),
.A2(n_1160),
.B(n_1157),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1117),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1192),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1133),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1179),
.A2(n_604),
.B1(n_1156),
.B2(n_1118),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1156),
.A2(n_604),
.B1(n_1188),
.B2(n_1182),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1121),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1155),
.A2(n_1160),
.B(n_1157),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1158),
.A2(n_604),
.B(n_1182),
.C(n_1179),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1158),
.A2(n_604),
.B(n_1182),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1111),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1156),
.A2(n_604),
.B1(n_1188),
.B2(n_1182),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1145),
.B(n_1146),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1179),
.A2(n_604),
.B1(n_1156),
.B2(n_1118),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1133),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1192),
.Y(n_1297)
);

BUFx8_ASAP7_75t_L g1298 ( 
.A(n_1159),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_1160),
.B(n_1157),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1151),
.A2(n_1202),
.B(n_1112),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1159),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1156),
.B(n_1149),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1117),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1203),
.A2(n_1112),
.A3(n_1088),
.B(n_1151),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1133),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1117),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1133),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1155),
.A2(n_1160),
.B(n_1157),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1192),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1117),
.Y(n_1310)
);

NOR2x1_ASAP7_75t_L g1311 ( 
.A(n_1080),
.B(n_1130),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1149),
.B(n_1169),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1291),
.A2(n_1272),
.B(n_1242),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1277),
.A2(n_1276),
.B1(n_1295),
.B2(n_1286),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1214),
.B(n_1276),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1215),
.B(n_1232),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1209),
.B(n_1286),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1290),
.A2(n_1287),
.B(n_1280),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1295),
.A2(n_1208),
.B1(n_1293),
.B2(n_1205),
.Y(n_1319)
);

O2A1O1Ixp5_ASAP7_75t_L g1320 ( 
.A1(n_1223),
.A2(n_1236),
.B(n_1290),
.C(n_1225),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1273),
.A2(n_1297),
.B(n_1284),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1233),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1278),
.B(n_1302),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1250),
.A2(n_1292),
.B1(n_1243),
.B2(n_1245),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1239),
.B(n_1263),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1207),
.B(n_1234),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1311),
.A2(n_1271),
.B1(n_1260),
.B2(n_1307),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1279),
.B(n_1281),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1273),
.A2(n_1284),
.B(n_1309),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1274),
.B(n_1285),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1221),
.A2(n_1251),
.B(n_1258),
.C(n_1270),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1273),
.A2(n_1297),
.B(n_1309),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1252),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1264),
.B(n_1296),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1305),
.B(n_1211),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1266),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1284),
.A2(n_1297),
.B(n_1309),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1218),
.A2(n_1229),
.B(n_1230),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1255),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1239),
.B(n_1263),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1226),
.B(n_1256),
.Y(n_1342)
);

NOR2xp67_ASAP7_75t_L g1343 ( 
.A(n_1246),
.B(n_1219),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1222),
.B(n_1228),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1222),
.B(n_1228),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1227),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1206),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1239),
.B(n_1267),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1269),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1257),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1258),
.B(n_1249),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1262),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1269),
.A2(n_1265),
.B(n_1240),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1266),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1275),
.B(n_1294),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1253),
.A2(n_1310),
.B1(n_1306),
.B2(n_1240),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1231),
.B(n_1244),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1253),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1238),
.A2(n_1220),
.B(n_1241),
.Y(n_1361)
);

OAI31xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1268),
.A2(n_1235),
.A3(n_1254),
.B(n_1248),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1261),
.B(n_1247),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1235),
.B(n_1303),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1235),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1283),
.A2(n_1204),
.B(n_1300),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1304),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1304),
.B(n_1288),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1235),
.B(n_1304),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1224),
.A2(n_1308),
.B(n_1210),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1282),
.A2(n_1289),
.B(n_1216),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1217),
.A2(n_1299),
.B(n_1298),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1298),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1301),
.B(n_1237),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1214),
.B(n_1156),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1279),
.B(n_1281),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1291),
.A2(n_1182),
.B(n_1158),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1237),
.B(n_1312),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1276),
.A2(n_604),
.B1(n_1156),
.B2(n_1188),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1292),
.B(n_958),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1277),
.A2(n_604),
.B1(n_1276),
.B2(n_1156),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1277),
.A2(n_604),
.B1(n_1276),
.B2(n_1156),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1291),
.A2(n_1182),
.B(n_1158),
.Y(n_1383)
);

OA22x2_ASAP7_75t_L g1384 ( 
.A1(n_1208),
.A2(n_1188),
.B1(n_1100),
.B2(n_1110),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1364),
.B(n_1369),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1349),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1352),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1333),
.B(n_1365),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1314),
.A2(n_1379),
.B1(n_1319),
.B2(n_1384),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1321),
.B(n_1330),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1377),
.A2(n_1383),
.B(n_1313),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1316),
.B(n_1351),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1350),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1366),
.B(n_1318),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_1367),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1349),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1368),
.B(n_1358),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1350),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1317),
.B(n_1315),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1362),
.B(n_1339),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1363),
.B(n_1339),
.Y(n_1403)
);

BUFx4f_ASAP7_75t_SL g1404 ( 
.A(n_1373),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1326),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1348),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1320),
.A2(n_1372),
.B(n_1334),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1326),
.B(n_1341),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1344),
.B(n_1345),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1348),
.A2(n_1331),
.B(n_1324),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1353),
.A2(n_1325),
.B(n_1341),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1340),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1370),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1341),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1355),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1375),
.B(n_1329),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1332),
.B(n_1328),
.C(n_1323),
.Y(n_1417)
);

OR2x2_ASAP7_75t_SL g1418 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1370),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1371),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1361),
.B(n_1371),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1342),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1371),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1335),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1413),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1397),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1401),
.B(n_1327),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1387),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1397),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1356),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1413),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1388),
.B(n_1378),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1391),
.B(n_1384),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1386),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1410),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1386),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1403),
.B(n_1360),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1395),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1389),
.A2(n_1390),
.B1(n_1417),
.B2(n_1400),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1400),
.B(n_1347),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1410),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1385),
.B(n_1374),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1408),
.B(n_1346),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1385),
.B(n_1408),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1393),
.B(n_1380),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1408),
.B(n_1402),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1394),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1410),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_R g1450 ( 
.A(n_1410),
.B(n_1354),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1449),
.A2(n_1420),
.B(n_1419),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1435),
.Y(n_1452)
);

OAI21xp33_ASAP7_75t_L g1453 ( 
.A1(n_1440),
.A2(n_1390),
.B(n_1389),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1447),
.B(n_1405),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1438),
.B(n_1418),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1426),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1440),
.A2(n_1417),
.B1(n_1392),
.B2(n_1418),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1434),
.A2(n_1422),
.B1(n_1402),
.B2(n_1416),
.C(n_1424),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1438),
.B(n_1418),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1446),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1425),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1428),
.B(n_1414),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1426),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1437),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1428),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1447),
.B(n_1405),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1450),
.A2(n_1395),
.B1(n_1416),
.B2(n_1422),
.C(n_1343),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1446),
.A2(n_1395),
.B1(n_1373),
.B2(n_1414),
.C(n_1354),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_R g1469 ( 
.A(n_1441),
.B(n_1322),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1429),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1438),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1427),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1447),
.B(n_1406),
.Y(n_1473)
);

OAI31xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1434),
.A2(n_1424),
.A3(n_1409),
.B(n_1395),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1429),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1430),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1431),
.B(n_1398),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1431),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1449),
.A2(n_1420),
.B(n_1423),
.Y(n_1479)
);

AOI33xp33_ASAP7_75t_L g1480 ( 
.A1(n_1434),
.A2(n_1412),
.A3(n_1396),
.B1(n_1394),
.B2(n_1399),
.B3(n_1415),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1445),
.B(n_1406),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_R g1482 ( 
.A(n_1444),
.B(n_1322),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1439),
.A2(n_1395),
.B1(n_1411),
.B2(n_1407),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1463),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1470),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1470),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1475),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1465),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1478),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1478),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1453),
.B(n_1337),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1428),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1462),
.B(n_1436),
.Y(n_1493)
);

INVx4_ASAP7_75t_SL g1494 ( 
.A(n_1452),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1453),
.A2(n_1442),
.B(n_1436),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1479),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1457),
.B(n_1439),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1464),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1452),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1464),
.Y(n_1500)
);

AO21x1_ASAP7_75t_L g1501 ( 
.A1(n_1457),
.A2(n_1431),
.B(n_1448),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1456),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1461),
.A2(n_1421),
.B(n_1432),
.Y(n_1503)
);

INVx4_ASAP7_75t_SL g1504 ( 
.A(n_1452),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1476),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1479),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1451),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1494),
.B(n_1466),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1494),
.B(n_1466),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1497),
.B(n_1439),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1503),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1491),
.B(n_1337),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1485),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1460),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1499),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1494),
.B(n_1436),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1442),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1495),
.B(n_1480),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1485),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1503),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1486),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1477),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1502),
.B(n_1477),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1499),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1507),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1495),
.B(n_1483),
.C(n_1458),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1504),
.B(n_1462),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1504),
.B(n_1462),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1503),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1504),
.B(n_1462),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1504),
.B(n_1442),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1507),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1497),
.A2(n_1467),
.B1(n_1468),
.B2(n_1459),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1486),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1487),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1505),
.B(n_1472),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1501),
.A2(n_1507),
.B(n_1506),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1497),
.B(n_1471),
.Y(n_1543)
);

NOR2x1_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1487),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1481),
.Y(n_1546)
);

OAI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1505),
.A2(n_1474),
.B(n_1469),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1511),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1513),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1533),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1527),
.A2(n_1482),
.B1(n_1455),
.B2(n_1459),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1513),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1533),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1519),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1484),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1518),
.B(n_1443),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1516),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1493),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1523),
.B(n_1484),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1540),
.B(n_1443),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1522),
.B(n_1498),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1508),
.B(n_1493),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1519),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1511),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1512),
.B(n_1404),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1522),
.B(n_1498),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1511),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1509),
.B(n_1493),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1521),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1520),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1521),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1547),
.B(n_1443),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1509),
.B(n_1493),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1529),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1538),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1526),
.B(n_1492),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1515),
.B(n_1433),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1544),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1500),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.B(n_1492),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1538),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1575),
.B(n_1524),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1544),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1558),
.B(n_1528),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1583),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1583),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1549),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1550),
.B(n_1571),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1549),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1553),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1582),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1548),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1557),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1524),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1579),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1555),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1530),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1539),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1562),
.B(n_1530),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1552),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1559),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1531),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1531),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1568),
.B(n_1534),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1559),
.B(n_1539),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1609)
);

OAI21xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1586),
.A2(n_1573),
.B(n_1574),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1598),
.B(n_1580),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1592),
.Y(n_1612)
);

OAI322xp33_ASAP7_75t_L g1613 ( 
.A1(n_1597),
.A2(n_1551),
.A3(n_1527),
.B1(n_1580),
.B2(n_1576),
.C1(n_1552),
.C2(n_1554),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1586),
.B(n_1574),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1603),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1593),
.B(n_1577),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1599),
.B(n_1582),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1590),
.A2(n_1537),
.B(n_1517),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1563),
.C(n_1554),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1592),
.Y(n_1620)
);

OAI311xp33_ASAP7_75t_L g1621 ( 
.A1(n_1596),
.A2(n_1557),
.A3(n_1543),
.B1(n_1561),
.C1(n_1566),
.Y(n_1621)
);

OAI322xp33_ASAP7_75t_L g1622 ( 
.A1(n_1600),
.A2(n_1569),
.A3(n_1563),
.B1(n_1572),
.B2(n_1576),
.C1(n_1517),
.C2(n_1566),
.Y(n_1622)
);

NAND2xp67_ASAP7_75t_L g1623 ( 
.A(n_1594),
.B(n_1543),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1594),
.A2(n_1564),
.B(n_1548),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1595),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1585),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1585),
.A2(n_1565),
.B(n_1517),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1585),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1585),
.A2(n_1557),
.B(n_1514),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1577),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1616),
.B(n_1600),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1612),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1626),
.B(n_1620),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

AOI222xp33_ASAP7_75t_L g1635 ( 
.A1(n_1615),
.A2(n_1588),
.B1(n_1589),
.B2(n_1591),
.C1(n_1587),
.C2(n_1602),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1625),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1614),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1611),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1617),
.B(n_1601),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1611),
.Y(n_1641)
);

AOI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1639),
.A2(n_1627),
.B(n_1628),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1632),
.A2(n_1621),
.B(n_1613),
.C(n_1622),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1637),
.B(n_1617),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1631),
.B(n_1610),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1635),
.B(n_1629),
.C(n_1628),
.Y(n_1646)
);

AOI211xp5_ASAP7_75t_L g1647 ( 
.A1(n_1632),
.A2(n_1618),
.B(n_1619),
.C(n_1630),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1641),
.Y(n_1648)
);

AOI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1638),
.A2(n_1601),
.B(n_1604),
.C(n_1605),
.Y(n_1649)
);

OAI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1640),
.A2(n_1510),
.B1(n_1595),
.B2(n_1608),
.C(n_1604),
.Y(n_1650)
);

AOI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1633),
.A2(n_1636),
.B(n_1634),
.C(n_1605),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1642),
.B(n_1606),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1648),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1643),
.A2(n_1635),
.B(n_1624),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1644),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1651),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1652),
.B(n_1649),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1654),
.B(n_1646),
.C(n_1647),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1653),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1656),
.A2(n_1650),
.B1(n_1645),
.B2(n_1588),
.C(n_1587),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1655),
.Y(n_1661)
);

OAI32xp33_ASAP7_75t_L g1662 ( 
.A1(n_1656),
.A2(n_1602),
.A3(n_1589),
.B1(n_1591),
.B2(n_1608),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1658),
.A2(n_1607),
.B1(n_1606),
.B2(n_1510),
.Y(n_1663)
);

NOR2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1661),
.B(n_1607),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1657),
.B(n_1623),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_R g1666 ( 
.A(n_1659),
.B(n_1404),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1660),
.B(n_1624),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1662),
.B(n_1594),
.C(n_1624),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1664),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1665),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1669),
.Y(n_1671)
);

OAI322xp33_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1668),
.A3(n_1670),
.B1(n_1663),
.B2(n_1666),
.C1(n_1609),
.C2(n_1570),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1672),
.B(n_1623),
.Y(n_1673)
);

OAI222xp33_ASAP7_75t_L g1674 ( 
.A1(n_1672),
.A2(n_1607),
.B1(n_1609),
.B2(n_1564),
.C1(n_1548),
.C2(n_1567),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1673),
.A2(n_1607),
.B1(n_1569),
.B2(n_1572),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1674),
.A2(n_1570),
.B1(n_1567),
.B2(n_1564),
.Y(n_1676)
);

AO22x1_ASAP7_75t_L g1677 ( 
.A1(n_1675),
.A2(n_1535),
.B1(n_1516),
.B2(n_1570),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_SL g1678 ( 
.A(n_1676),
.B(n_1560),
.C(n_1578),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1677),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1678),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1567),
.B1(n_1536),
.B2(n_1525),
.Y(n_1681)
);

OAI222xp33_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1679),
.B1(n_1525),
.B2(n_1536),
.C1(n_1510),
.C2(n_1535),
.Y(n_1682)
);

AOI322xp5_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1535),
.A3(n_1516),
.B1(n_1581),
.B2(n_1546),
.C1(n_1532),
.C2(n_1520),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1542),
.B1(n_1545),
.B2(n_1535),
.C(n_1516),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1581),
.B(n_1546),
.C(n_1496),
.Y(n_1685)
);


endmodule