module fake_jpeg_16947_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_17),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_14),
.C(n_15),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_42),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_25),
.B1(n_15),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_55),
.B1(n_24),
.B2(n_12),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_20),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_61),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_15),
.B1(n_25),
.B2(n_17),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_59),
.B(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_12),
.B1(n_24),
.B2(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_51),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_37),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_76),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_74),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_2),
.B(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_56),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_82),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_84),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_47),
.B(n_54),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_67),
.B(n_66),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_79),
.B(n_67),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_66),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_55),
.B1(n_56),
.B2(n_34),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_69),
.B1(n_78),
.B2(n_77),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_63),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_101),
.A3(n_106),
.B1(n_86),
.B2(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_75),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_65),
.B(n_69),
.C(n_71),
.D(n_64),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_19),
.C(n_22),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_18),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_21),
.C(n_22),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_115),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_89),
.C(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_30),
.C(n_40),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_104),
.B1(n_105),
.B2(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_97),
.B1(n_103),
.B2(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_126),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_109),
.B(n_114),
.Y(n_125)
);

OAI31xp33_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_122),
.A3(n_117),
.B(n_7),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_93),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_4),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_40),
.C(n_14),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_5),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_125),
.A3(n_61),
.B1(n_34),
.B2(n_40),
.C1(n_7),
.C2(n_6),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_16),
.A3(n_107),
.B1(n_113),
.B2(n_88),
.C(n_137),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_61),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_135),
.C(n_16),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_140),
.Y(n_142)
);


endmodule