module real_aes_6782_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_693;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_0), .A2(n_201), .B1(n_360), .B2(n_362), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_1), .A2(n_87), .B1(n_364), .B2(n_367), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_2), .A2(n_210), .B1(n_407), .B2(n_472), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_3), .A2(n_218), .B1(n_396), .B2(n_524), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_4), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_5), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_6), .B(n_393), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_7), .Y(n_658) );
AOI22xp5_ASAP7_75t_SL g408 ( .A1(n_8), .A2(n_51), .B1(n_409), .B2(n_411), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_9), .A2(n_20), .B1(n_302), .B2(n_305), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_10), .A2(n_147), .B1(n_481), .B2(n_507), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_11), .B(n_444), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_12), .A2(n_59), .B1(n_567), .B2(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_13), .A2(n_108), .B1(n_282), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_14), .A2(n_103), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_15), .A2(n_190), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_16), .A2(n_126), .B1(n_343), .B2(n_387), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_17), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g610 ( .A1(n_18), .A2(n_91), .B1(n_114), .B2(n_309), .C1(n_316), .C2(n_494), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_19), .A2(n_166), .B1(n_269), .B2(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_21), .A2(n_30), .B1(n_290), .B2(n_318), .Y(n_529) );
INVx1_ASAP7_75t_L g448 ( .A(n_22), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_23), .A2(n_157), .B1(n_360), .B2(n_373), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_24), .Y(n_675) );
AOI22xp5_ASAP7_75t_SL g405 ( .A1(n_25), .A2(n_221), .B1(n_406), .B2(n_407), .Y(n_405) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_26), .A2(n_67), .B1(n_249), .B2(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g648 ( .A(n_26), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_27), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_28), .A2(n_32), .B1(n_318), .B2(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_29), .A2(n_53), .B1(n_480), .B2(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_31), .B(n_391), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_33), .A2(n_142), .B1(n_361), .B2(n_370), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_34), .A2(n_64), .B1(n_476), .B2(n_570), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_35), .A2(n_175), .B1(n_259), .B2(n_376), .Y(n_701) );
AOI22xp5_ASAP7_75t_SL g399 ( .A1(n_36), .A2(n_123), .B1(n_299), .B2(n_400), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g308 ( .A1(n_37), .A2(n_109), .B1(n_173), .B2(n_309), .C1(n_311), .C2(n_316), .Y(n_308) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_38), .A2(n_69), .B1(n_249), .B2(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g649 ( .A(n_38), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_39), .A2(n_167), .B1(n_376), .B2(n_409), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_40), .A2(n_81), .B1(n_569), .B2(n_570), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_41), .A2(n_55), .B1(n_290), .B2(n_446), .Y(n_587) );
AOI222xp33_ASAP7_75t_L g588 ( .A1(n_42), .A2(n_141), .B1(n_184), .B2(n_439), .C1(n_589), .C2(n_590), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_43), .A2(n_143), .B1(n_305), .B2(n_377), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_44), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_45), .A2(n_200), .B1(n_360), .B2(n_483), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_46), .Y(n_334) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_47), .A2(n_66), .B1(n_467), .B2(n_468), .Y(n_466) );
XOR2xp5_ASAP7_75t_L g596 ( .A(n_48), .B(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_49), .A2(n_202), .B1(n_296), .B2(n_299), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_50), .A2(n_455), .B1(n_456), .B2(n_484), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_50), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g285 ( .A1(n_52), .A2(n_120), .B1(n_286), .B2(n_290), .Y(n_285) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_54), .A2(n_111), .B1(n_299), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_56), .A2(n_132), .B1(n_524), .B2(n_525), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_57), .A2(n_99), .B1(n_403), .B2(n_508), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_58), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_60), .A2(n_212), .B1(n_396), .B2(n_397), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_61), .B(n_556), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_62), .A2(n_139), .B1(n_474), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_63), .A2(n_68), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_65), .A2(n_73), .B1(n_704), .B2(n_705), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_70), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_71), .B(n_281), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_72), .A2(n_160), .B1(n_423), .B2(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g230 ( .A(n_74), .Y(n_230) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_75), .A2(n_137), .B1(n_406), .B2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_76), .A2(n_96), .B1(n_259), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_77), .A2(n_125), .B1(n_312), .B2(n_318), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_78), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_79), .A2(n_95), .B1(n_242), .B2(n_259), .Y(n_241) );
INVx1_ASAP7_75t_L g228 ( .A(n_80), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_82), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_83), .A2(n_93), .B1(n_403), .B2(n_422), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_84), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_85), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_86), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_88), .A2(n_128), .B1(n_302), .B2(n_570), .Y(n_580) );
OA22x2_ASAP7_75t_L g611 ( .A1(n_89), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_89), .Y(n_612) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_90), .A2(n_92), .B1(n_367), .B2(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_94), .A2(n_113), .B1(n_286), .B2(n_338), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_97), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_98), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_100), .A2(n_107), .B1(n_259), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_101), .A2(n_153), .B1(n_318), .B2(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_102), .A2(n_145), .B1(n_266), .B2(n_269), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_104), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_105), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_106), .A2(n_223), .B(n_232), .C(n_650), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_110), .A2(n_652), .B1(n_685), .B2(n_686), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_110), .Y(n_685) );
XOR2x2_ASAP7_75t_L g543 ( .A(n_112), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_115), .A2(n_187), .B1(n_373), .B2(n_376), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_116), .Y(n_350) );
XNOR2x2_ASAP7_75t_L g575 ( .A(n_117), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_118), .A2(n_138), .B1(n_411), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_119), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_121), .Y(n_385) );
INVx2_ASAP7_75t_L g231 ( .A(n_122), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_124), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_127), .A2(n_151), .B1(n_569), .B2(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_129), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_130), .A2(n_186), .B1(n_422), .B2(n_423), .Y(n_421) );
OA22x2_ASAP7_75t_L g516 ( .A1(n_131), .A2(n_517), .B1(n_518), .B2(n_539), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_131), .Y(n_517) );
INVx1_ASAP7_75t_L g511 ( .A(n_133), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_134), .B(n_589), .Y(n_622) );
AND2x6_ASAP7_75t_L g227 ( .A(n_135), .B(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_135), .Y(n_642) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_136), .A2(n_196), .B1(n_249), .B2(n_253), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_140), .Y(n_550) );
AOI22xp5_ASAP7_75t_SL g401 ( .A1(n_144), .A2(n_194), .B1(n_402), .B2(n_403), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_146), .A2(n_203), .B1(n_406), .B2(n_632), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_148), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_149), .A2(n_211), .B1(n_397), .B2(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_150), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_152), .B(n_281), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_154), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_155), .A2(n_208), .B1(n_306), .B2(n_364), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_156), .B(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_158), .A2(n_162), .B1(n_483), .B2(n_599), .Y(n_633) );
AO22x2_ASAP7_75t_L g258 ( .A1(n_159), .A2(n_204), .B1(n_249), .B2(n_250), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_161), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_163), .A2(n_181), .B1(n_312), .B2(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_164), .B(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_192), .B1(n_361), .B2(n_370), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_168), .A2(n_185), .B1(n_400), .B2(n_407), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_169), .Y(n_274) );
INVx1_ASAP7_75t_L g412 ( .A(n_170), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_171), .A2(n_188), .B1(n_411), .B2(n_533), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_172), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_174), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_176), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_177), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_178), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_179), .A2(n_180), .B1(n_411), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_182), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_183), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_183), .A2(n_694), .B1(n_697), .B2(n_724), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_189), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_191), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_193), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_195), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_196), .B(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_197), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_198), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_199), .Y(n_671) );
INVx1_ASAP7_75t_L g645 ( .A(n_204), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_205), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_206), .B(n_312), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_207), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_209), .B(n_281), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_213), .Y(n_332) );
INVx1_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
INVx1_ASAP7_75t_L g251 ( .A(n_214), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_215), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_216), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_217), .A2(n_220), .B1(n_302), .B2(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_219), .B(n_391), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_228), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_229), .A2(n_640), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_513), .B1(n_635), .B2(n_636), .C(n_637), .Y(n_232) );
INVx1_ASAP7_75t_L g635 ( .A(n_233), .Y(n_635) );
XOR2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_414), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B1(n_322), .B2(n_323), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
XOR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_321), .Y(n_238) );
NAND4xp75_ASAP7_75t_L g239 ( .A(n_240), .B(n_273), .C(n_294), .D(n_308), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_265), .Y(n_240) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx5_ASAP7_75t_SL g370 ( .A(n_243), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_243), .A2(n_297), .B1(n_426), .B2(n_427), .Y(n_425) );
INVx4_ASAP7_75t_L g533 ( .A(n_243), .Y(n_533) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_243), .Y(n_655) );
INVx11_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx11_ASAP7_75t_L g410 ( .A(n_244), .Y(n_410) );
AND2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_254), .Y(n_244) );
AND2x4_ASAP7_75t_L g284 ( .A(n_245), .B(n_279), .Y(n_284) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g330 ( .A(n_246), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
AND2x2_ASAP7_75t_L g263 ( .A(n_247), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g278 ( .A(n_247), .B(n_252), .Y(n_278) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g289 ( .A(n_248), .B(n_256), .Y(n_289) );
AND2x2_ASAP7_75t_L g293 ( .A(n_248), .B(n_252), .Y(n_293) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g253 ( .A(n_251), .Y(n_253) );
INVx2_ASAP7_75t_L g264 ( .A(n_252), .Y(n_264) );
INVx1_ASAP7_75t_L g288 ( .A(n_252), .Y(n_288) );
AND2x2_ASAP7_75t_L g268 ( .A(n_254), .B(n_263), .Y(n_268) );
AND2x4_ASAP7_75t_L g298 ( .A(n_254), .B(n_278), .Y(n_298) );
AND2x6_ASAP7_75t_L g310 ( .A(n_254), .B(n_293), .Y(n_310) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
AND2x2_ASAP7_75t_L g279 ( .A(n_255), .B(n_258), .Y(n_279) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_256), .B(n_258), .Y(n_262) );
AND2x2_ASAP7_75t_L g271 ( .A(n_256), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
INVx1_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
BUFx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_SL g371 ( .A(n_260), .Y(n_371) );
BUFx2_ASAP7_75t_L g407 ( .A(n_260), .Y(n_407) );
BUFx2_ASAP7_75t_SL g423 ( .A(n_260), .Y(n_423) );
BUFx3_ASAP7_75t_L g503 ( .A(n_260), .Y(n_503) );
BUFx3_ASAP7_75t_L g632 ( .A(n_260), .Y(n_632) );
INVx1_ASAP7_75t_L g664 ( .A(n_260), .Y(n_664) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x2_ASAP7_75t_L g510 ( .A(n_261), .B(n_349), .Y(n_510) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x6_ASAP7_75t_L g307 ( .A(n_262), .B(n_288), .Y(n_307) );
AND2x2_ASAP7_75t_L g270 ( .A(n_263), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g300 ( .A(n_263), .B(n_279), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_263), .B(n_271), .Y(n_434) );
AND2x2_ASAP7_75t_L g314 ( .A(n_264), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g349 ( .A(n_264), .Y(n_349) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g628 ( .A(n_267), .Y(n_628) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_268), .Y(n_361) );
BUFx2_ASAP7_75t_SL g400 ( .A(n_268), .Y(n_400) );
BUFx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx3_ASAP7_75t_L g375 ( .A(n_270), .Y(n_375) );
BUFx3_ASAP7_75t_L g406 ( .A(n_270), .Y(n_406) );
BUFx3_ASAP7_75t_L g608 ( .A(n_270), .Y(n_608) );
AND2x2_ASAP7_75t_L g304 ( .A(n_271), .B(n_278), .Y(n_304) );
INVx1_ASAP7_75t_L g292 ( .A(n_272), .Y(n_292) );
OA211x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B(n_280), .C(n_285), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx3_ASAP7_75t_L g333 ( .A(n_277), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x6_ASAP7_75t_L g393 ( .A(n_278), .B(n_279), .Y(n_393) );
INVx1_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g444 ( .A(n_283), .Y(n_444) );
INVx2_ASAP7_75t_L g497 ( .A(n_283), .Y(n_497) );
INVx2_ASAP7_75t_L g603 ( .A(n_283), .Y(n_603) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g396 ( .A(n_286), .Y(n_396) );
INVx1_ASAP7_75t_L g447 ( .A(n_286), .Y(n_447) );
BUFx2_ASAP7_75t_L g525 ( .A(n_286), .Y(n_525) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g313 ( .A(n_289), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g319 ( .A(n_289), .B(n_320), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_289), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g469 ( .A(n_290), .Y(n_469) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_SL g397 ( .A(n_291), .Y(n_397) );
BUFx3_ASAP7_75t_L g494 ( .A(n_291), .Y(n_494) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g355 ( .A(n_292), .Y(n_355) );
INVx1_ASAP7_75t_L g354 ( .A(n_293), .Y(n_354) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_301), .Y(n_294) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g411 ( .A(n_297), .Y(n_411) );
INVx2_ASAP7_75t_L g704 ( .A(n_297), .Y(n_704) );
INVx6_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx3_ASAP7_75t_L g362 ( .A(n_298), .Y(n_362) );
BUFx3_ASAP7_75t_L g507 ( .A(n_298), .Y(n_507) );
BUFx3_ASAP7_75t_L g599 ( .A(n_298), .Y(n_599) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx3_ASAP7_75t_L g377 ( .A(n_300), .Y(n_377) );
BUFx3_ASAP7_75t_L g422 ( .A(n_300), .Y(n_422) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_300), .Y(n_474) );
INVx2_ASAP7_75t_L g662 ( .A(n_300), .Y(n_662) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx4_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
BUFx3_ASAP7_75t_L g477 ( .A(n_303), .Y(n_477) );
INVx5_ASAP7_75t_L g508 ( .A(n_303), .Y(n_508) );
INVx1_ASAP7_75t_L g537 ( .A(n_303), .Y(n_537) );
INVx8_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g403 ( .A(n_306), .Y(n_403) );
BUFx4f_ASAP7_75t_SL g708 ( .A(n_306), .Y(n_708) );
INVx6_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g367 ( .A(n_307), .Y(n_367) );
INVx1_ASAP7_75t_L g570 ( .A(n_307), .Y(n_570) );
INVx2_ASAP7_75t_L g459 ( .A(n_309), .Y(n_459) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_SL g340 ( .A(n_310), .Y(n_340) );
INVx4_ASAP7_75t_L g384 ( .A(n_310), .Y(n_384) );
INVx2_ASAP7_75t_L g492 ( .A(n_310), .Y(n_492) );
BUFx3_ASAP7_75t_L g589 ( .A(n_310), .Y(n_589) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx4_ASAP7_75t_L g388 ( .A(n_312), .Y(n_388) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_313), .Y(n_524) );
BUFx2_ASAP7_75t_L g590 ( .A(n_313), .Y(n_590) );
BUFx4f_ASAP7_75t_SL g674 ( .A(n_313), .Y(n_674) );
INVx1_ASAP7_75t_L g320 ( .A(n_315), .Y(n_320) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx4f_ASAP7_75t_SL g439 ( .A(n_318), .Y(n_439) );
BUFx12f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_319), .Y(n_344) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_319), .Y(n_557) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_378), .B1(n_379), .B2(n_413), .Y(n_323) );
INVx2_ASAP7_75t_L g413 ( .A(n_324), .Y(n_413) );
XNOR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_357), .Y(n_326) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_335), .C(n_346), .Y(n_327) );
OAI22xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_332), .B1(n_333), .B2(n_334), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g549 ( .A(n_330), .Y(n_549) );
BUFx3_ASAP7_75t_L g618 ( .A(n_330), .Y(n_618) );
INVx2_ASAP7_75t_L g552 ( .A(n_333), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_333), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_333), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
BUFx3_ASAP7_75t_L g723 ( .A(n_333), .Y(n_723) );
OAI222xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B1(n_340), .B2(n_341), .C1(n_342), .C2(n_345), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx4f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI22xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_350), .B1(n_351), .B2(n_356), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_348), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_348), .A2(n_353), .B1(n_624), .B2(n_625), .Y(n_623) );
INVx4_ASAP7_75t_L g678 ( .A(n_348), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_351), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g714 ( .A(n_352), .Y(n_714) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g684 ( .A(n_353), .Y(n_684) );
OR2x6_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_368), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_363), .Y(n_358) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g430 ( .A(n_361), .Y(n_430) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_361), .Y(n_480) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_366), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx4f_ASAP7_75t_SL g481 ( .A(n_375), .Y(n_481) );
BUFx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
XOR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_412), .Y(n_380) );
NAND3x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_398), .C(n_404), .Y(n_381) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_383), .B(n_389), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_386), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g436 ( .A1(n_384), .A2(n_437), .B(n_438), .Y(n_436) );
BUFx2_ASAP7_75t_L g527 ( .A(n_384), .Y(n_527) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_394), .C(n_395), .Y(n_389) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g586 ( .A(n_392), .Y(n_586) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
BUFx2_ASAP7_75t_L g464 ( .A(n_393), .Y(n_464) );
BUFx4f_ASAP7_75t_L g604 ( .A(n_393), .Y(n_604) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g706 ( .A(n_406), .Y(n_706) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx4_ASAP7_75t_L g483 ( .A(n_410), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_449), .B2(n_450), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
XOR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_448), .Y(n_417) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_419), .B(n_435), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_425), .C(n_428), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_428) );
INVx2_ASAP7_75t_L g567 ( .A(n_430), .Y(n_567) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_440), .Y(n_435) );
INVx1_ASAP7_75t_L g682 ( .A(n_439), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .C(n_445), .Y(n_440) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g467 ( .A(n_447), .Y(n_467) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_452), .B1(n_485), .B2(n_512), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g484 ( .A(n_456), .Y(n_484) );
NAND3x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_470), .C(n_478), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_460), .B(n_461), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .C(n_466), .Y(n_462) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g579 ( .A(n_473), .Y(n_579) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g512 ( .A(n_485), .Y(n_512) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
XOR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_511), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_493), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_492), .A2(n_554), .B1(n_555), .B2(n_558), .C(n_559), .Y(n_553) );
OAI222xp33_ASAP7_75t_L g672 ( .A1(n_492), .A2(n_673), .B1(n_675), .B2(n_676), .C1(n_677), .C2(n_679), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g715 ( .A1(n_492), .A2(n_716), .B1(n_717), .B2(n_718), .C(n_719), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .C(n_499), .Y(n_495) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_509), .Y(n_505) );
INVx3_ASAP7_75t_L g657 ( .A(n_507), .Y(n_657) );
INVx1_ASAP7_75t_L g636 ( .A(n_513), .Y(n_636) );
XOR2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_593), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_540), .B1(n_591), .B2(n_592), .Y(n_514) );
INVx1_ASAP7_75t_L g591 ( .A(n_515), .Y(n_591) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g539 ( .A(n_518), .Y(n_539) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
NOR2xp67_ASAP7_75t_SL g519 ( .A(n_520), .B(n_526), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .C(n_523), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g592 ( .A(n_540), .Y(n_592) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_543), .B1(n_574), .B2(n_575), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_564), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_553), .C(n_560), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_550), .B2(n_551), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_SL g670 ( .A(n_549), .Y(n_670) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_571), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND4xp75_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .C(n_584), .D(n_588), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_SL g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g717 ( .A(n_590), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_611), .B2(n_634), .Y(n_593) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_595), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND5xp2_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .C(n_601), .D(n_606), .E(n_610), .Y(n_597) );
AND2x2_ASAP7_75t_SL g601 ( .A(n_602), .B(n_605), .Y(n_601) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
BUFx3_ASAP7_75t_L g660 ( .A(n_608), .Y(n_660) );
INVx2_ASAP7_75t_SL g634 ( .A(n_611), .Y(n_634) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND3x1_ASAP7_75t_L g614 ( .A(n_615), .B(n_626), .C(n_630), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .C(n_623), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_643), .Y(n_638) );
OR2x2_ASAP7_75t_SL g727 ( .A(n_639), .B(n_644), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_641), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_641), .B(n_690), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g690 ( .A(n_642), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OAI322xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_687), .A3(n_688), .B1(n_691), .B2(n_694), .C1(n_695), .C2(n_725), .Y(n_650) );
INVx1_ASAP7_75t_L g686 ( .A(n_652), .Y(n_686) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_653), .B(n_667), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_661), .Y(n_653) );
OAI221xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_656), .B1(n_657), .B2(n_658), .C(n_659), .Y(n_654) );
OAI221xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_663), .B1(n_664), .B2(n_665), .C(n_666), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_672), .C(n_680), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_670), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_SL g712 ( .A(n_678), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_680) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g724 ( .A(n_697), .Y(n_724) );
AND2x2_ASAP7_75t_SL g697 ( .A(n_698), .B(n_709), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .Y(n_702) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR3xp33_ASAP7_75t_SL g709 ( .A(n_710), .B(n_715), .C(n_720), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
endmodule