module fake_jpeg_14852_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_20),
.Y(n_79)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_17),
.B1(n_21),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_70)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_28),
.B1(n_17),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_64),
.B1(n_73),
.B2(n_25),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_40),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_70),
.B1(n_34),
.B2(n_53),
.Y(n_88)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_40),
.B1(n_25),
.B2(n_23),
.Y(n_95)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_38),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_24),
.B1(n_23),
.B2(n_27),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_22),
.Y(n_105)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_36),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_83),
.C(n_85),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_14),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_95),
.B1(n_101),
.B2(n_90),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_0),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_20),
.B1(n_30),
.B2(n_16),
.Y(n_136)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_32),
.C(n_66),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_75),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_33),
.B1(n_26),
.B2(n_19),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_24),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_33),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_116),
.B1(n_123),
.B2(n_127),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_91),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_0),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_121),
.B1(n_92),
.B2(n_14),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_76),
.B1(n_81),
.B2(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_92),
.Y(n_124)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_104),
.B1(n_87),
.B2(n_68),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_60),
.B1(n_30),
.B2(n_27),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_106),
.Y(n_146)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_20),
.B(n_16),
.Y(n_155)
);

AO21x2_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_97),
.B(n_102),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_153),
.B(n_156),
.C(n_110),
.Y(n_169)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_154),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_83),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_149),
.C(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_150),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_94),
.B1(n_90),
.B2(n_86),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_152),
.B1(n_165),
.B2(n_136),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_86),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_116),
.B1(n_111),
.B2(n_125),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_75),
.B(n_32),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_87),
.B1(n_12),
.B2(n_13),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_32),
.C(n_55),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_11),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_15),
.B(n_1),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_110),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_165)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_185),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_169),
.A2(n_184),
.B(n_194),
.C(n_167),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_68),
.B1(n_71),
.B2(n_59),
.Y(n_201)
);

CKINVDCx10_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_173),
.B(n_179),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_117),
.B1(n_122),
.B2(n_131),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_180),
.B1(n_183),
.B2(n_62),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_117),
.B1(n_131),
.B2(n_126),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_187),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_134),
.B1(n_128),
.B2(n_114),
.Y(n_183)
);

NAND2x1p5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_129),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_68),
.B(n_59),
.C(n_55),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_62),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_195),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_15),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_32),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_159),
.C(n_144),
.Y(n_198)
);

CKINVDCx10_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_15),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_146),
.B(n_152),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_204),
.B(n_214),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_208),
.C(n_213),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_147),
.B1(n_155),
.B2(n_161),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_218),
.B1(n_219),
.B2(n_168),
.Y(n_228)
);

NOR4xp25_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_162),
.C(n_32),
.D(n_55),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_212),
.B1(n_202),
.B2(n_215),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_55),
.C(n_62),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_193),
.C(n_189),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_186),
.B1(n_182),
.B2(n_176),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_13),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_183),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_12),
.B(n_11),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_169),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_177),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_226),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_169),
.B1(n_174),
.B2(n_167),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_171),
.B1(n_180),
.B2(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_217),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_231),
.B1(n_232),
.B2(n_218),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_175),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_236),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_214),
.B(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_176),
.B1(n_182),
.B2(n_196),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_196),
.B1(n_188),
.B2(n_2),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_188),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_214),
.B1(n_2),
.B2(n_3),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_199),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_0),
.Y(n_251)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_245),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_209),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_229),
.A2(n_207),
.B1(n_205),
.B2(n_208),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_224),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_205),
.C(n_207),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_223),
.C(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_256),
.C(n_265),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_223),
.C(n_220),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_230),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_258),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_253),
.B1(n_247),
.B2(n_248),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_233),
.B(n_236),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_243),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_227),
.C(n_237),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_237),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_240),
.C(n_4),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_272),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_276),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_242),
.B1(n_246),
.B2(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.C(n_277),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_3),
.C(n_4),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_5),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_263),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_256),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.C(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_271),
.B(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_286),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_264),
.B1(n_255),
.B2(n_8),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_255),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_287),
.B(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_290),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_277),
.B(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_264),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_276),
.B(n_7),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_284),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_295),
.C(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_285),
.B(n_292),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_294),
.B(n_6),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_6),
.B(n_8),
.Y(n_304)
);


endmodule