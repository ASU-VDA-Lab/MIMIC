module fake_jpeg_26576_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_4),
.B(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_53),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_18),
.B1(n_16),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_51),
.B1(n_23),
.B2(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_25),
.B1(n_16),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_55),
.B1(n_56),
.B2(n_41),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_22),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_17),
.C(n_20),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_39),
.C(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_72),
.Y(n_94)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_36),
.B1(n_22),
.B2(n_28),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_75),
.B1(n_23),
.B2(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_36),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_39),
.B(n_50),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_28),
.B1(n_33),
.B2(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_30),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_27),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_46),
.Y(n_91)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_96),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_48),
.B(n_2),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_80),
.B(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_45),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_100),
.Y(n_119)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_45),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_104),
.B1(n_19),
.B2(n_4),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_45),
.B1(n_37),
.B2(n_39),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_50),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_39),
.C(n_20),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_39),
.C(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_2),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_78),
.B1(n_84),
.B2(n_74),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_118),
.B1(n_136),
.B2(n_111),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_135),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_130),
.B(n_110),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_20),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_131),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_66),
.B(n_62),
.C(n_23),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_62),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_110),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_50),
.B(n_19),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_107),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_19),
.C(n_4),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_112),
.C(n_108),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_147),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_151),
.B(n_158),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_156),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_102),
.B(n_90),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_162),
.B1(n_122),
.B2(n_120),
.Y(n_171)
);

XOR2x2_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_90),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_96),
.C(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_123),
.C(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_132),
.B1(n_87),
.B2(n_6),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_3),
.C(n_5),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_170),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_152),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_135),
.C(n_116),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_118),
.C(n_117),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_127),
.B1(n_136),
.B2(n_134),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_101),
.C(n_134),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_180),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_101),
.C(n_87),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_143),
.B1(n_139),
.B2(n_159),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_3),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_5),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_185),
.C(n_164),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_150),
.B(n_151),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_189),
.A2(n_190),
.B1(n_196),
.B2(n_201),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_175),
.B(n_140),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_167),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_163),
.B1(n_162),
.B2(n_157),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_142),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_139),
.B(n_150),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_173),
.C(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_210),
.C(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_169),
.C(n_165),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_208),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_207),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_174),
.C(n_179),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_183),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_183),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_193),
.C(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_191),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_200),
.B1(n_201),
.B2(n_194),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_216),
.B1(n_144),
.B2(n_223),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_225),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_200),
.B1(n_168),
.B2(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_222),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

AOI31xp33_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_210),
.A3(n_211),
.B(n_161),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_142),
.Y(n_232)
);

AOI31xp33_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_6),
.B(n_7),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_235),
.B(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_8),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_8),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_229),
.B1(n_228),
.B2(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_9),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_9),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_12),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_241),
.B(n_234),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_246),
.B(n_12),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_248),
.Y(n_250)
);


endmodule