module fake_jpeg_7499_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_30),
.B1(n_23),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_67),
.B1(n_22),
.B2(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_60),
.B1(n_63),
.B2(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_32),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_59),
.CON(n_82),
.SN(n_82)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_33),
.B(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_31),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_32),
.Y(n_67)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_74),
.B1(n_79),
.B2(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_30),
.B1(n_33),
.B2(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_38),
.B1(n_33),
.B2(n_37),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_84),
.B1(n_36),
.B2(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_81)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_84)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_22),
.B1(n_28),
.B2(n_25),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_91),
.B1(n_51),
.B2(n_44),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_14),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_63),
.B(n_61),
.C(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_83),
.B1(n_62),
.B2(n_53),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_107),
.B(n_114),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_45),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_44),
.B1(n_26),
.B2(n_17),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_118),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_73),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_39),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_17),
.B1(n_26),
.B2(n_16),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_135),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_112),
.B1(n_95),
.B2(n_116),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_127),
.B1(n_128),
.B2(n_132),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_134),
.B1(n_94),
.B2(n_117),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_85),
.B1(n_75),
.B2(n_71),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_123),
.A2(n_125),
.B1(n_137),
.B2(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_114),
.B1(n_107),
.B2(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_90),
.B1(n_71),
.B2(n_64),
.Y(n_127)
);

OAI22x1_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_39),
.B1(n_42),
.B2(n_34),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_57),
.B1(n_77),
.B2(n_83),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_70),
.B(n_24),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_140),
.B(n_146),
.Y(n_160)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_92),
.B1(n_88),
.B2(n_76),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_70),
.B(n_24),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_88),
.B1(n_92),
.B2(n_76),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_42),
.B(n_76),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_156),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_94),
.B1(n_99),
.B2(n_96),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_170),
.B1(n_50),
.B2(n_42),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_39),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_164),
.Y(n_177)
);

OAI22x1_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_19),
.B1(n_16),
.B2(n_24),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_128),
.B1(n_136),
.B2(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_157),
.B(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_41),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_17),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_39),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_166),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_34),
.C(n_41),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_73),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_73),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_39),
.C(n_34),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_42),
.C(n_41),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_86),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_122),
.B(n_26),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_136),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_176),
.A2(n_183),
.B1(n_185),
.B2(n_188),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_142),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_164),
.C(n_174),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_154),
.Y(n_209)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_54),
.B1(n_68),
.B2(n_78),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_158),
.A2(n_154),
.B1(n_148),
.B2(n_149),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_161),
.B(n_171),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_130),
.B1(n_138),
.B2(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_130),
.B1(n_138),
.B2(n_129),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_200),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_117),
.B1(n_78),
.B2(n_54),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_190),
.A2(n_19),
.B1(n_16),
.B2(n_42),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_68),
.B1(n_86),
.B2(n_50),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_192),
.B1(n_148),
.B2(n_155),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_68),
.B1(n_50),
.B2(n_40),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_19),
.B1(n_42),
.B2(n_40),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_159),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_203),
.C(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_165),
.C(n_166),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_160),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_177),
.C(n_181),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_221),
.C(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_214),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_219),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_163),
.B1(n_153),
.B2(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_185),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_160),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_42),
.CI(n_41),
.CON(n_218),
.SN(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_220),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_41),
.C(n_40),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_40),
.C(n_42),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_40),
.C(n_31),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_203),
.C(n_221),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_225),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_239),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_206),
.B(n_204),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_31),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_237),
.C(n_245),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_188),
.B(n_176),
.C(n_183),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_242),
.B1(n_219),
.B2(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_186),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_180),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_241),
.B(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_191),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_202),
.A2(n_192),
.B(n_190),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_246),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_216),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_15),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_263),
.B1(n_229),
.B2(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_256),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_206),
.B1(n_218),
.B2(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_253),
.B1(n_258),
.B2(n_13),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_218),
.B1(n_223),
.B2(n_19),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_31),
.C(n_1),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_257),
.C(n_260),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_31),
.C(n_1),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_227),
.C(n_245),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_230),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_0),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_247),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_229),
.B1(n_238),
.B2(n_237),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_246),
.B1(n_241),
.B2(n_226),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_227),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_272),
.B(n_274),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_12),
.C(n_11),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_11),
.C(n_2),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_2),
.C(n_3),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_282),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_257),
.B1(n_255),
.B2(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_3),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_258),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_252),
.B(n_253),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_276),
.B(n_4),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_266),
.B(n_263),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_3),
.C(n_4),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_0),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_5),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_288),
.C(n_5),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_3),
.C(n_4),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_289),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_294),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_7),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_298),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_5),
.B(n_6),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_287),
.B(n_8),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_10),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_285),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_7),
.B(n_8),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_294),
.C(n_292),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_304),
.B(n_305),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_311),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_300),
.B(n_310),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.C(n_303),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_10),
.B(n_7),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.Y(n_318)
);


endmodule