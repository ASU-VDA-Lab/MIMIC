module real_jpeg_26795_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_0),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_256)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_1),
.Y(n_114)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_146),
.B(n_160),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_34),
.B1(n_63),
.B2(n_64),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_3),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_32),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_32),
.B(n_172),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_129),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_11),
.B(n_63),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_3),
.B(n_87),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_3),
.A2(n_108),
.B1(n_109),
.B2(n_223),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_126),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_126),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_126),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_8),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_10),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_124),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_124),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_124),
.Y(n_215)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_12),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_131),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_131),
.Y(n_223)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_79),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_69),
.C(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_20),
.A2(n_21),
.B1(n_69),
.B2(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_23),
.A2(n_37),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_23),
.A2(n_37),
.B1(n_137),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_23),
.A2(n_263),
.B(n_282),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_24),
.B(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_24),
.A2(n_30),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_24),
.A2(n_84),
.B(n_283),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_25),
.B(n_32),
.Y(n_143)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_27),
.B(n_129),
.CON(n_128),
.SN(n_128)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_29),
.A2(n_31),
.B1(n_128),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_30),
.B(n_283),
.Y(n_282)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_31),
.A2(n_44),
.A3(n_47),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_33),
.A2(n_37),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_37),
.B(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_67),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_57),
.C(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_42),
.A2(n_75),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_43),
.A2(n_55),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_43),
.A2(n_55),
.B1(n_123),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_43),
.A2(n_55),
.B1(n_156),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_43),
.A2(n_55),
.B1(n_77),
.B2(n_301),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_45),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_45),
.B(n_48),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_45),
.A2(n_61),
.B(n_129),
.C(n_200),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_52),
.A2(n_87),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_57),
.A2(n_67),
.B1(n_74),
.B2(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_65),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_65),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_58),
.A2(n_62),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_58),
.A2(n_180),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_58),
.A2(n_62),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_58),
.A2(n_62),
.B1(n_179),
.B2(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_58),
.A2(n_62),
.B1(n_103),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_58),
.A2(n_119),
.B(n_256),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_62),
.B(n_129),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_64),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_66),
.B(n_120),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.C(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_69),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_73),
.B(n_322),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_74),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_78),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_75),
.A2(n_78),
.B(n_88),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_311),
.A3(n_323),
.B1(n_329),
.B2(n_330),
.C(n_332),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_293),
.B(n_310),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_269),
.B(n_292),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_161),
.B(n_246),
.C(n_268),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_148),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_99),
.B(n_148),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_132),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_101),
.B(n_116),
.C(n_132),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_102),
.B(n_107),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_104),
.B(n_190),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_110),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_108),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_108),
.A2(n_147),
.B1(n_215),
.B2(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_108),
.A2(n_147),
.B(n_288),
.Y(n_287)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_109),
.B(n_129),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_112),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_127),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_134),
.B(n_139),
.C(n_141),
.Y(n_266)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_144),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_149),
.A2(n_150),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_245),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_238),
.B(n_244),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_191),
.B(n_237),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_181),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_165),
.B(n_181),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_174),
.C(n_177),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_166),
.A2(n_167),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_169),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_210),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_188),
.C(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_231),
.B(n_236),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_211),
.B(n_230),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_194),
.B(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_196),
.B1(n_199),
.B2(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_219),
.B(n_229),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_217),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_224),
.B(n_228),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_266),
.B2(n_267),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_258),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_258),
.C(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_261),
.C(n_265),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_271),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_291),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_284),
.B2(n_285),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_285),
.C(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_287),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_289),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_304),
.B(n_307),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_295),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_308),
.B2(n_309),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_303),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_303),
.C(n_309),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_313),
.C(n_319),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_313),
.B1(n_314),
.B2(n_328),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_321),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_321),
.Y(n_330)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);


endmodule