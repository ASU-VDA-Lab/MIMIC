module real_jpeg_32860_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_0),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_1),
.A2(n_295),
.B1(n_296),
.B2(n_299),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_1),
.A2(n_295),
.B1(n_445),
.B2(n_449),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_1),
.A2(n_295),
.B1(n_542),
.B2(n_544),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_2),
.A2(n_162),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_2),
.A2(n_217),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_2),
.A2(n_217),
.B1(n_459),
.B2(n_461),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_2),
.A2(n_217),
.B1(n_581),
.B2(n_583),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_3),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_3),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_4),
.A2(n_387),
.B1(n_389),
.B2(n_390),
.Y(n_386)
);

INVx2_ASAP7_75t_R g389 ( 
.A(n_4),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_4),
.A2(n_389),
.B1(n_481),
.B2(n_484),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_4),
.A2(n_389),
.B1(n_563),
.B2(n_566),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_51),
.B1(n_54),
.B2(n_58),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_58),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_5),
.A2(n_58),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_5),
.A2(n_58),
.B1(n_411),
.B2(n_414),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_44),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_6),
.A2(n_44),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_6),
.A2(n_44),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_7),
.A2(n_161),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_7),
.A2(n_161),
.B1(n_421),
.B2(n_423),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_7),
.A2(n_161),
.B1(n_532),
.B2(n_535),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_8),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_8),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_8),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_13),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_36),
.B1(n_45),
.B2(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_14),
.B(n_167),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_14),
.A2(n_196),
.A3(n_203),
.B1(n_204),
.B2(n_209),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_71),
.B1(n_232),
.B2(n_236),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_14),
.A2(n_339),
.B(n_342),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_14),
.B(n_343),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_15),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_87)
);

INVx2_ASAP7_75t_R g93 ( 
.A(n_15),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_15),
.A2(n_93),
.B1(n_252),
.B2(n_255),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_15),
.A2(n_93),
.B1(n_356),
.B2(n_361),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_15),
.A2(n_93),
.B1(n_467),
.B2(n_471),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_16),
.A2(n_433),
.B1(n_434),
.B2(n_488),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_16),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_16),
.A2(n_352),
.B1(n_488),
.B2(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_17),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_17),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_17),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_18),
.A2(n_433),
.B1(n_435),
.B2(n_436),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_18),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_18),
.A2(n_435),
.B1(n_518),
.B2(n_522),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_19),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_19),
.Y(n_206)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_19),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_548),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_498),
.B(n_546),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_399),
.B(n_495),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_311),
.B(n_398),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_263),
.B(n_310),
.Y(n_29)
);

AOI21x1_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_191),
.B(n_262),
.Y(n_30)
);

OAI21x1_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_153),
.B(n_190),
.Y(n_31)
);

AOI22x1_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_82),
.B1(n_151),
.B2(n_152),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_72),
.B(n_81),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_61),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_35),
.B(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_45),
.B1(n_50),
.B2(n_59),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_40),
.Y(n_160)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_40),
.Y(n_164)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_45),
.A2(n_87),
.B1(n_96),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_45),
.A2(n_386),
.B1(n_432),
.B2(n_438),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_45),
.A2(n_74),
.B1(n_432),
.B2(n_487),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_45),
.A2(n_487),
.B(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_46),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_46),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_47),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_53),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_59),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_62),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_62),
.A2(n_135),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_62),
.A2(n_135),
.B1(n_272),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_62),
.A2(n_135),
.B1(n_348),
.B2(n_444),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_63),
.Y(n_258)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AO21x2_ASAP7_75t_L g135 ( 
.A1(n_64),
.A2(n_123),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_115),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_114),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_71),
.B(n_210),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_SL g301 ( 
.A(n_71),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_101),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_95),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_85),
.A2(n_158),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_85),
.A2(n_214),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_85),
.A2(n_294),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_R g293 ( 
.A(n_99),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_100),
.Y(n_384)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_128),
.B2(n_150),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_102),
.B(n_150),
.Y(n_154)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_120),
.B2(n_122),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_108),
.Y(n_299)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_108),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_117),
.Y(n_279)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_134),
.B1(n_141),
.B2(n_149),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_134),
.A2(n_251),
.B1(n_258),
.B2(n_259),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_134),
.A2(n_258),
.B1(n_569),
.B2(n_573),
.Y(n_568)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_135),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_135),
.A2(n_444),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_135),
.A2(n_479),
.B1(n_480),
.B2(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_140),
.Y(n_351)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_143),
.Y(n_483)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_147),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_148),
.Y(n_448)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_148),
.Y(n_521)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_148),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_149),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_155),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_179),
.C(n_188),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_160),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_179),
.B1(n_188),
.B2(n_189),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_167),
.A2(n_539),
.B1(n_540),
.B2(n_541),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_167),
.A2(n_540),
.B1(n_541),
.B2(n_562),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_168),
.A2(n_204),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_174),
.B2(n_176),
.Y(n_168)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_169),
.Y(n_572)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_175),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_175),
.Y(n_450)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g262 ( 
.A(n_192),
.B(n_193),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_220),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_250),
.C(n_261),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_212),
.B1(n_218),
.B2(n_219),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_201),
.Y(n_422)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_201),
.Y(n_545)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g306 ( 
.A(n_206),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_206),
.Y(n_565)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_250),
.B1(n_260),
.B2(n_261),
.Y(n_220)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_231),
.B1(n_239),
.B2(n_240),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_222),
.A2(n_239),
.B1(n_240),
.B2(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_222),
.A2(n_239),
.B1(n_284),
.B2(n_355),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g419 ( 
.A1(n_222),
.A2(n_239),
.B1(n_355),
.B2(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_222),
.A2(n_239),
.B1(n_420),
.B2(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_222),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_227),
.Y(n_543)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_228),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_229),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_230),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_238),
.Y(n_289)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_248),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_248),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_249),
.Y(n_426)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_258),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_265),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_282),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_280),
.B2(n_281),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_268),
.B(n_280),
.C(n_282),
.Y(n_397)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_283),
.B(n_291),
.C(n_301),
.Y(n_364)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_300),
.B2(n_301),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_316),
.B1(n_324),
.B2(n_338),
.Y(n_315)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_302),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_302),
.A2(n_324),
.B1(n_410),
.B2(n_466),
.Y(n_465)
);

OAI22x1_ASAP7_75t_SL g529 ( 
.A1(n_302),
.A2(n_324),
.B1(n_466),
.B2(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_302),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_306),
.Y(n_362)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_397),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g398 ( 
.A(n_312),
.B(n_397),
.Y(n_398)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_363),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_313),
.B(n_364),
.C(n_365),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_346),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_315),
.B(n_347),
.C(n_354),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_316),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_322),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_323),
.Y(n_582)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_325),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_325),
.B(n_531),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_331),
.B1(n_333),
.B2(n_335),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_330),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_334),
.Y(n_585)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx4f_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVx3_ASAP7_75t_SL g472 ( 
.A(n_341),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_383),
.B1(n_394),
.B2(n_396),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_366),
.B(n_396),
.Y(n_427)
);

OAI32xp33_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_370),
.A3(n_374),
.B1(n_376),
.B2(n_382),
.Y(n_366)
);

OAI32xp33_ASAP7_75t_L g395 ( 
.A1(n_367),
.A2(n_370),
.A3(n_374),
.B1(n_376),
.B2(n_382),
.Y(n_395)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx11_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_490),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_451),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_402),
.B(n_451),
.C(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_428),
.C(n_430),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_403),
.B(n_494),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_427),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_418),
.B2(n_419),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_427),
.C(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_417),
.Y(n_470)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_426),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_429),
.B(n_430),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_443),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_443),
.Y(n_476)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_442),
.Y(n_515)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_502),
.C(n_503),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_474),
.B1(n_475),
.B2(n_489),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_456),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_456),
.A2(n_476),
.B1(n_489),
.B2(n_504),
.Y(n_503)
);

AO22x1_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_464),
.B1(n_465),
.B2(n_473),
.Y(n_456)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_464),
.B(n_473),
.C(n_504),
.Y(n_506)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_476),
.Y(n_504)
);

INVxp33_ASAP7_75t_SL g502 ( 
.A(n_477),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_486),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_478),
.B(n_486),
.Y(n_527)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_493),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_505),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_501),
.B(n_505),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_506),
.B(n_509),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g554 ( 
.A(n_506),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_526),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_508),
.B(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_516),
.B2(n_525),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_510),
.A2(n_511),
.B1(n_577),
.B2(n_578),
.Y(n_576)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_511),
.B(n_516),
.Y(n_588)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_516),
.Y(n_525)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_517),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_528),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_527),
.B(n_557),
.C(n_558),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_538),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_529),
.Y(n_558)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVxp33_ASAP7_75t_SL g546 ( 
.A(n_547),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_R g548 ( 
.A(n_549),
.B(n_589),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_555),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_550),
.B(n_555),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_551),
.A2(n_552),
.B(n_553),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_559),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_575),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_561),
.A2(n_568),
.B(n_574),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_568),
.Y(n_574)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx8_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_588),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_587),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_586),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_582),
.Y(n_581)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);


endmodule