module fake_netlist_6_2305_n_2420 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2420);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2420;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_822;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_907;
wire n_1446;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_2101;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_1165;
wire n_2008;
wire n_2192;
wire n_2345;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_890;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_1270;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_1222;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2322;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_875;
wire n_1678;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_740;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g705 ( 
.A(n_569),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_186),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_175),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_462),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_239),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_234),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_456),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_633),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_628),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_135),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_404),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_550),
.Y(n_716)
);

CKINVDCx14_ASAP7_75t_R g717 ( 
.A(n_607),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_7),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_585),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_593),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_702),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_508),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_499),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_559),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_201),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_554),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_638),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_590),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_586),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_653),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_664),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_207),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_619),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_572),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_435),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_563),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_207),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_173),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_283),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_377),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_576),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_183),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_420),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_663),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_596),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_613),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_630),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_38),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_551),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_98),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_650),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_654),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_623),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_684),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_624),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_448),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_655),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_357),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_286),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_243),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_553),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_172),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_608),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_579),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_21),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_657),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_682),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_697),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_651),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_399),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_587),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_365),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_615),
.Y(n_773)
);

CKINVDCx16_ASAP7_75t_R g774 ( 
.A(n_284),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_662),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_162),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_652),
.Y(n_777)
);

CKINVDCx14_ASAP7_75t_R g778 ( 
.A(n_406),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_629),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_47),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_605),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_601),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_374),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_375),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_575),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_552),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_610),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_614),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_469),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_485),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_627),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_20),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_671),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_414),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_39),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_255),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_363),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_10),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_670),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_561),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_82),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_302),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_681),
.Y(n_804)
);

CKINVDCx16_ASAP7_75t_R g805 ( 
.A(n_187),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_389),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_645),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_458),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_606),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_667),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_646),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_196),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_135),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_142),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_617),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_349),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_127),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_102),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_441),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_656),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_163),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_64),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_666),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_142),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_685),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_620),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_157),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_410),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_288),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_291),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_228),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_163),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_636),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_266),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_339),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_597),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_603),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_665),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_600),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_282),
.Y(n_840)
);

BUFx2_ASAP7_75t_SL g841 ( 
.A(n_641),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_173),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_224),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_595),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_251),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_195),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_634),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_165),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_350),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_403),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_126),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_612),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_604),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_345),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_189),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_253),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_599),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_543),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_58),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_98),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_431),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_532),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_618),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_616),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_589),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_696),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_378),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_132),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_317),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_254),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_416),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_584),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_162),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_609),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_274),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_299),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_197),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_141),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_555),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_464),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_480),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_647),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_611),
.Y(n_883)
);

BUFx5_ASAP7_75t_L g884 ( 
.A(n_643),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_233),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_227),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_96),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_683),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_117),
.Y(n_889)
);

BUFx10_ASAP7_75t_L g890 ( 
.A(n_677),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_693),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_548),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_231),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_351),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_75),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_621),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_10),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_591),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_251),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_592),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_461),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_602),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_335),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_632),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_9),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_15),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_659),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_279),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_302),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_275),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_219),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_688),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_194),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_55),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_261),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_62),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_49),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_265),
.Y(n_918)
);

CKINVDCx14_ASAP7_75t_R g919 ( 
.A(n_230),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_564),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_676),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_542),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_504),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_367),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_512),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_495),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_644),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_193),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_509),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_658),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_141),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_639),
.Y(n_932)
);

BUFx10_ASAP7_75t_L g933 ( 
.A(n_224),
.Y(n_933)
);

CKINVDCx14_ASAP7_75t_R g934 ( 
.A(n_257),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_625),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_156),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_649),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_326),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_384),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_476),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_364),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_661),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_16),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_669),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_594),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_336),
.Y(n_946)
);

CKINVDCx16_ASAP7_75t_R g947 ( 
.A(n_626),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_687),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_549),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_521),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_642),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_186),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_673),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_58),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_635),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_330),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_203),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_598),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_519),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_254),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_303),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_686),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_71),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_379),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_631),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_263),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_237),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_249),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_219),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_622),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_108),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_560),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_84),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_660),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_73),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_402),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_668),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_230),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_478),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_648),
.Y(n_980)
);

BUFx10_ASAP7_75t_L g981 ( 
.A(n_474),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_588),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_291),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_146),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_352),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_640),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_18),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_263),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_562),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_280),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_884),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_708),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_712),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_725),
.Y(n_994)
);

NOR2xp67_ASAP7_75t_L g995 ( 
.A(n_765),
.B(n_0),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_713),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_748),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_715),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_884),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_711),
.B(n_1),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_884),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_719),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_759),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_868),
.B(n_0),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_760),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_919),
.B(n_1),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_793),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_729),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_802),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_747),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_803),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_818),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_723),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_934),
.B(n_2),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_737),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_821),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_726),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_727),
.Y(n_1018)
);

CKINVDCx16_ASAP7_75t_R g1019 ( 
.A(n_774),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_834),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_805),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_992),
.B(n_717),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_1019),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_994),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_997),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_993),
.B(n_778),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_1005),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1007),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_1006),
.B(n_879),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1011),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_1012),
.Y(n_1031)
);

CKINVDCx8_ASAP7_75t_R g1032 ( 
.A(n_998),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1016),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1002),
.B(n_858),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_1020),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1003),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1013),
.B(n_757),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1003),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_991),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1017),
.B(n_836),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1018),
.B(n_850),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1009),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1009),
.B(n_989),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_999),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1001),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1014),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1000),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1004),
.B(n_937),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_995),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_996),
.B(n_764),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1008),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1036),
.B(n_786),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_1032),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1022),
.B(n_724),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1045),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_1046),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1028),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1039),
.Y(n_1058)
);

OAI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_1047),
.A2(n_870),
.B1(n_875),
.B2(n_846),
.C(n_845),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_1039),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1037),
.B(n_780),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_1023),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1044),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1050),
.A2(n_838),
.B1(n_849),
.B2(n_828),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_1039),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1040),
.B(n_740),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1024),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_1033),
.Y(n_1068)
);

INVx8_ASAP7_75t_L g1069 ( 
.A(n_1026),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1038),
.B(n_951),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1021),
.Y(n_1071)
);

OR2x2_ASAP7_75t_SL g1072 ( 
.A(n_1049),
.B(n_947),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_1029),
.B(n_722),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1030),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1042),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1025),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1048),
.B(n_706),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1025),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1027),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1027),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1031),
.Y(n_1081)
);

AO21x2_ASAP7_75t_L g1082 ( 
.A1(n_1034),
.A2(n_716),
.B(n_705),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_1031),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_1035),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1043),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_1041),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1051),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1039),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1028),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1022),
.B(n_758),
.Y(n_1090)
);

AND2x2_ASAP7_75t_SL g1091 ( 
.A(n_1023),
.B(n_940),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1037),
.B(n_1010),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1039),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1036),
.B(n_974),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_1023),
.B(n_876),
.Y(n_1095)
);

AO22x2_ASAP7_75t_L g1096 ( 
.A1(n_1073),
.A2(n_796),
.B1(n_812),
.B2(n_707),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1057),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1061),
.B(n_720),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1089),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1055),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1055),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1086),
.A2(n_985),
.B1(n_728),
.B2(n_790),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_1077),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1053),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1074),
.Y(n_1105)
);

AO22x2_ASAP7_75t_L g1106 ( 
.A1(n_1071),
.A2(n_984),
.B1(n_813),
.B2(n_916),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1067),
.Y(n_1107)
);

OR2x6_ASAP7_75t_L g1108 ( 
.A(n_1062),
.B(n_841),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1085),
.B(n_754),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1076),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1079),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1083),
.B(n_877),
.Y(n_1112)
);

NAND2x1p5_ASAP7_75t_L g1113 ( 
.A(n_1075),
.B(n_809),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1063),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1063),
.Y(n_1115)
);

NAND2x1p5_ASAP7_75t_L g1116 ( 
.A(n_1056),
.B(n_721),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1078),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_SL g1118 ( 
.A1(n_1092),
.A2(n_718),
.B1(n_750),
.B2(n_709),
.Y(n_1118)
);

AO22x2_ASAP7_75t_L g1119 ( 
.A1(n_1077),
.A2(n_990),
.B1(n_885),
.B2(n_895),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1080),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1064),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1087),
.B(n_878),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_1084),
.B(n_785),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1066),
.B(n_1054),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1081),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1090),
.A2(n_804),
.B1(n_735),
.B2(n_741),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1052),
.B(n_840),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1068),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1058),
.B(n_730),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1068),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1088),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1093),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1060),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1070),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1094),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1082),
.Y(n_1136)
);

AO22x2_ASAP7_75t_L g1137 ( 
.A1(n_1091),
.A2(n_913),
.B1(n_936),
.B2(n_905),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1095),
.B(n_1069),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_1069),
.B(n_938),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1095),
.Y(n_1140)
);

AO22x2_ASAP7_75t_L g1141 ( 
.A1(n_1072),
.A2(n_966),
.B1(n_957),
.B2(n_952),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1072),
.B(n_710),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1065),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1059),
.Y(n_1144)
);

AO22x2_ASAP7_75t_L g1145 ( 
.A1(n_1073),
.A2(n_969),
.B1(n_776),
.B2(n_824),
.Y(n_1145)
);

AO22x2_ASAP7_75t_L g1146 ( 
.A1(n_1073),
.A2(n_910),
.B1(n_928),
.B2(n_742),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1057),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1057),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1085),
.B(n_840),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1057),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1077),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1061),
.B(n_733),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1095),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1057),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1057),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1061),
.B(n_734),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1067),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1053),
.Y(n_1158)
);

OAI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_1059),
.A2(n_983),
.B1(n_791),
.B2(n_756),
.C(n_761),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1057),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1061),
.B(n_745),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1057),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1083),
.B(n_755),
.Y(n_1163)
);

AO22x2_ASAP7_75t_L g1164 ( 
.A1(n_1085),
.A2(n_767),
.B1(n_769),
.B2(n_766),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1085),
.B(n_775),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1086),
.A2(n_743),
.B1(n_744),
.B2(n_731),
.Y(n_1167)
);

AO22x2_ASAP7_75t_L g1168 ( 
.A1(n_1085),
.A2(n_794),
.B1(n_795),
.B2(n_789),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1061),
.B(n_798),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1061),
.B(n_806),
.Y(n_1170)
);

AO22x2_ASAP7_75t_L g1171 ( 
.A1(n_1085),
.A2(n_808),
.B1(n_835),
.B2(n_807),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1067),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1067),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1057),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_1077),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1085),
.B(n_839),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1067),
.Y(n_1177)
);

OAI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_1059),
.A2(n_925),
.B1(n_865),
.B2(n_854),
.C(n_857),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1085),
.B(n_972),
.Y(n_1179)
);

AO22x2_ASAP7_75t_L g1180 ( 
.A1(n_1085),
.A2(n_852),
.B1(n_862),
.B2(n_853),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_L g1181 ( 
.A(n_1086),
.B(n_884),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1085),
.B(n_977),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1057),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1067),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1057),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_SL g1186 ( 
.A(n_1064),
.B(n_856),
.C(n_831),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1057),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1053),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_L g1189 ( 
.A(n_1086),
.B(n_884),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1085),
.B(n_911),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1061),
.B(n_714),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1057),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_1095),
.Y(n_1193)
);

OAI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1059),
.A2(n_949),
.B1(n_866),
.B2(n_871),
.C(n_874),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1057),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1067),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1124),
.B(n_746),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1098),
.B(n_749),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1191),
.B(n_864),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1121),
.B(n_860),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1152),
.B(n_751),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1156),
.B(n_752),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1161),
.B(n_753),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1169),
.B(n_763),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1170),
.B(n_1103),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1128),
.B(n_882),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1151),
.B(n_768),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1175),
.B(n_770),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1149),
.B(n_911),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1123),
.B(n_771),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1100),
.B(n_891),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1190),
.B(n_933),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1101),
.B(n_1097),
.Y(n_1213)
);

AND2x2_ASAP7_75t_SL g1214 ( 
.A(n_1138),
.B(n_883),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1134),
.B(n_869),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1109),
.B(n_772),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1102),
.B(n_773),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1135),
.B(n_897),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1165),
.B(n_777),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1099),
.B(n_896),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1176),
.B(n_779),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1147),
.B(n_781),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1148),
.B(n_902),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1150),
.B(n_782),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1154),
.B(n_783),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1155),
.B(n_784),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1160),
.B(n_921),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1162),
.B(n_1166),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1127),
.B(n_933),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1104),
.B(n_968),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1174),
.B(n_787),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1183),
.B(n_788),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1185),
.B(n_792),
.Y(n_1233)
);

NAND2xp33_ASAP7_75t_SL g1234 ( 
.A(n_1158),
.B(n_800),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1108),
.B(n_732),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1187),
.B(n_801),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_SL g1237 ( 
.A(n_1188),
.B(n_810),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1192),
.B(n_811),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1195),
.B(n_815),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1193),
.B(n_816),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1144),
.B(n_819),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1193),
.B(n_820),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1167),
.B(n_1113),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1130),
.B(n_922),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_SL g1245 ( 
.A(n_1140),
.B(n_823),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1126),
.B(n_825),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1142),
.B(n_1114),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1153),
.B(n_826),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1115),
.B(n_833),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1105),
.B(n_837),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_SL g1251 ( 
.A(n_1179),
.B(n_844),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1110),
.B(n_939),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1163),
.B(n_847),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1111),
.B(n_861),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1157),
.B(n_948),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1172),
.B(n_863),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1173),
.B(n_867),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1177),
.B(n_872),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_SL g1259 ( 
.A(n_1182),
.B(n_880),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1184),
.B(n_956),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1196),
.B(n_881),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1117),
.B(n_888),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1120),
.B(n_892),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1125),
.B(n_894),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_SL g1265 ( 
.A(n_1112),
.B(n_898),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_SL g1266 ( 
.A(n_1143),
.B(n_900),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1107),
.B(n_901),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1116),
.B(n_907),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1122),
.B(n_923),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1108),
.B(n_738),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1136),
.B(n_924),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1133),
.B(n_926),
.Y(n_1272)
);

NAND2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1131),
.B(n_927),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1118),
.B(n_929),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1129),
.B(n_930),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1132),
.B(n_935),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1186),
.B(n_941),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1146),
.B(n_942),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1145),
.B(n_944),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_SL g1280 ( 
.A(n_1141),
.B(n_945),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1181),
.B(n_959),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1137),
.B(n_946),
.Y(n_1282)
);

NAND2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1096),
.B(n_950),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1189),
.B(n_965),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1164),
.B(n_953),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1164),
.B(n_955),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1168),
.B(n_958),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1168),
.B(n_962),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_SL g1289 ( 
.A(n_1171),
.B(n_970),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1171),
.B(n_976),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1180),
.B(n_980),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1180),
.B(n_986),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1119),
.B(n_722),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1139),
.B(n_739),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1139),
.B(n_979),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1106),
.B(n_736),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1159),
.B(n_903),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1178),
.B(n_736),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1194),
.B(n_890),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1124),
.B(n_890),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1121),
.B(n_762),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1124),
.B(n_920),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1124),
.B(n_920),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1124),
.B(n_912),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1124),
.B(n_981),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1124),
.B(n_932),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1124),
.B(n_981),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1124),
.B(n_964),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1124),
.B(n_884),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1124),
.B(n_904),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1124),
.B(n_904),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_SL g1312 ( 
.A(n_1121),
.B(n_797),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1124),
.B(n_904),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1128),
.B(n_329),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1124),
.B(n_982),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1124),
.B(n_982),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1124),
.B(n_982),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1124),
.B(n_799),
.Y(n_1318)
);

NAND2xp33_ASAP7_75t_SL g1319 ( 
.A(n_1121),
.B(n_814),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1124),
.B(n_817),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1124),
.B(n_822),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1124),
.B(n_827),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1124),
.B(n_829),
.Y(n_1323)
);

NAND2xp33_ASAP7_75t_SL g1324 ( 
.A(n_1121),
.B(n_830),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1124),
.B(n_832),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1124),
.B(n_842),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1124),
.B(n_843),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1124),
.B(n_848),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1103),
.B(n_851),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1124),
.B(n_855),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1124),
.B(n_859),
.Y(n_1331)
);

NAND2xp33_ASAP7_75t_SL g1332 ( 
.A(n_1121),
.B(n_873),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1124),
.B(n_886),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1124),
.B(n_887),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1124),
.B(n_889),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1124),
.B(n_893),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1124),
.B(n_899),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1124),
.B(n_906),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1124),
.B(n_908),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1124),
.B(n_909),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1124),
.B(n_914),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1128),
.B(n_331),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1124),
.B(n_915),
.Y(n_1343)
);

NAND2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1121),
.B(n_917),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1124),
.B(n_918),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1124),
.B(n_931),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1124),
.B(n_943),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1124),
.B(n_954),
.Y(n_1348)
);

INVx5_ASAP7_75t_L g1349 ( 
.A(n_1235),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1320),
.B(n_960),
.Y(n_1350)
);

AOI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1199),
.A2(n_963),
.B(n_961),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1209),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1212),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_R g1354 ( 
.A(n_1234),
.B(n_967),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1329),
.B(n_971),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1327),
.B(n_973),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1335),
.B(n_975),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1304),
.B(n_1306),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1308),
.A2(n_987),
.B(n_988),
.C(n_978),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1214),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1213),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1247),
.A2(n_1243),
.B(n_1313),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1228),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1206),
.B(n_332),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1206),
.B(n_333),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1314),
.B(n_334),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1244),
.B(n_337),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_1216),
.B(n_338),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1211),
.A2(n_341),
.B(n_340),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1252),
.A2(n_343),
.B(n_342),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1255),
.A2(n_346),
.B(n_344),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1246),
.A2(n_348),
.B(n_353),
.C(n_347),
.Y(n_1372)
);

AOI221x1_ASAP7_75t_L g1373 ( 
.A1(n_1283),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1309),
.A2(n_355),
.B(n_354),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1281),
.A2(n_358),
.B(n_356),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1260),
.Y(n_1376)
);

NAND2x1_ASAP7_75t_L g1377 ( 
.A(n_1314),
.B(n_1342),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1244),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1284),
.A2(n_360),
.B(n_359),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1342),
.B(n_5),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1318),
.A2(n_362),
.B(n_361),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1220),
.A2(n_368),
.B(n_366),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1223),
.A2(n_1227),
.B(n_1310),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1295),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1276),
.A2(n_370),
.B(n_369),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1200),
.B(n_6),
.Y(n_1386)
);

CKINVDCx8_ASAP7_75t_R g1387 ( 
.A(n_1297),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1311),
.A2(n_372),
.B(n_371),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1230),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1297),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1229),
.B(n_7),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1205),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1315),
.A2(n_376),
.B(n_373),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1316),
.A2(n_381),
.B(n_380),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1317),
.A2(n_383),
.B(n_382),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1256),
.A2(n_386),
.B(n_385),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1272),
.A2(n_388),
.B(n_387),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1197),
.A2(n_1254),
.B(n_1224),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1257),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1321),
.A2(n_391),
.B1(n_392),
.B2(n_390),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1270),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1271),
.A2(n_698),
.A3(n_699),
.B(n_695),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1258),
.A2(n_394),
.B(n_393),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1322),
.B(n_8),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1237),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1301),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1261),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1241),
.A2(n_11),
.B(n_8),
.C(n_9),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1323),
.A2(n_396),
.B(n_395),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1240),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1198),
.A2(n_398),
.B(n_397),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1325),
.B(n_11),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1326),
.A2(n_401),
.B(n_400),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1328),
.A2(n_407),
.B(n_405),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1222),
.A2(n_409),
.B(n_408),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1330),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_1416)
);

O2A1O1Ixp5_ASAP7_75t_L g1417 ( 
.A1(n_1300),
.A2(n_700),
.B(n_701),
.C(n_694),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1225),
.A2(n_1231),
.B(n_1226),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1232),
.A2(n_412),
.B(n_411),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1331),
.B(n_12),
.Y(n_1420)
);

O2A1O1Ixp5_ASAP7_75t_SL g1421 ( 
.A1(n_1296),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1249),
.A2(n_415),
.B(n_413),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1333),
.B(n_16),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1262),
.A2(n_418),
.B(n_417),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1275),
.A2(n_421),
.B(n_419),
.Y(n_1425)
);

AO32x2_ASAP7_75t_L g1426 ( 
.A1(n_1285),
.A2(n_19),
.A3(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1334),
.A2(n_1337),
.B(n_1338),
.C(n_1336),
.Y(n_1427)
);

AO31x2_ASAP7_75t_L g1428 ( 
.A1(n_1289),
.A2(n_703),
.A3(n_704),
.B(n_692),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1339),
.A2(n_21),
.B(n_17),
.C(n_19),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1263),
.A2(n_423),
.B(n_422),
.Y(n_1430)
);

AOI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1264),
.A2(n_425),
.B(n_424),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1340),
.A2(n_427),
.B(n_426),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1341),
.B(n_22),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1343),
.B(n_22),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1233),
.A2(n_429),
.B(n_428),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1293),
.A2(n_23),
.B(n_24),
.Y(n_1436)
);

AOI211x1_ASAP7_75t_L g1437 ( 
.A1(n_1286),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1236),
.A2(n_432),
.B(n_430),
.Y(n_1438)
);

INVx5_ASAP7_75t_L g1439 ( 
.A(n_1248),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1267),
.A2(n_1278),
.B(n_1250),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1347),
.B(n_25),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1312),
.Y(n_1443)
);

NOR2xp67_ASAP7_75t_L g1444 ( 
.A(n_1302),
.B(n_433),
.Y(n_1444)
);

AO31x2_ASAP7_75t_L g1445 ( 
.A1(n_1291),
.A2(n_679),
.A3(n_680),
.B(n_678),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1348),
.B(n_434),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1201),
.B(n_26),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1202),
.A2(n_437),
.B1(n_438),
.B2(n_436),
.Y(n_1448)
);

AOI21xp33_ASAP7_75t_L g1449 ( 
.A1(n_1277),
.A2(n_27),
.B(n_28),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1238),
.A2(n_440),
.B(n_439),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1280),
.A2(n_691),
.A3(n_690),
.B(n_443),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1239),
.A2(n_1279),
.B(n_1268),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1319),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1203),
.B(n_27),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1273),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_L g1456 ( 
.A(n_1251),
.B(n_442),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1242),
.B(n_1253),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1204),
.B(n_28),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1324),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1303),
.B(n_29),
.Y(n_1460)
);

AO31x2_ASAP7_75t_L g1461 ( 
.A1(n_1287),
.A2(n_674),
.A3(n_675),
.B(n_672),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1210),
.A2(n_445),
.B(n_444),
.Y(n_1462)
);

AO21x1_ASAP7_75t_L g1463 ( 
.A1(n_1288),
.A2(n_29),
.B(n_30),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1290),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1362),
.A2(n_1292),
.B(n_1221),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1423),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1383),
.A2(n_1422),
.B(n_1403),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1361),
.B(n_1305),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1363),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1443),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1384),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1352),
.B(n_1332),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1350),
.B(n_1344),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1355),
.B(n_1274),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1373),
.A2(n_1307),
.A3(n_1282),
.B(n_1259),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1358),
.A2(n_1219),
.B(n_1208),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1377),
.B(n_1207),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1398),
.A2(n_1427),
.B(n_1418),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1405),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1353),
.B(n_1215),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1356),
.B(n_1217),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1452),
.A2(n_1299),
.B(n_1298),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1369),
.A2(n_1266),
.B(n_1269),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1384),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1459),
.Y(n_1485)
);

NOR2x1_ASAP7_75t_R g1486 ( 
.A(n_1349),
.B(n_1218),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1349),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_R g1488 ( 
.A(n_1439),
.B(n_1294),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1378),
.B(n_1245),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1401),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1392),
.Y(n_1491)
);

NAND2x1p5_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1265),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1387),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1456),
.A2(n_447),
.B(n_446),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1391),
.B(n_30),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1406),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1434),
.B(n_31),
.C(n_32),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1463),
.A2(n_450),
.B(n_449),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1412),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1380),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1441),
.A2(n_452),
.B(n_451),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1381),
.A2(n_454),
.B(n_453),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1390),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1376),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1366),
.B(n_455),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1396),
.A2(n_459),
.B(n_457),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1407),
.Y(n_1507)
);

AOI22x1_ASAP7_75t_L g1508 ( 
.A1(n_1455),
.A2(n_463),
.B1(n_465),
.B2(n_460),
.Y(n_1508)
);

AND2x6_ASAP7_75t_L g1509 ( 
.A(n_1364),
.B(n_466),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1388),
.A2(n_468),
.B(n_467),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1365),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1404),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1357),
.A2(n_471),
.B(n_470),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1351),
.B(n_31),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1446),
.A2(n_473),
.B(n_472),
.Y(n_1515)
);

AO31x2_ASAP7_75t_L g1516 ( 
.A1(n_1464),
.A2(n_477),
.A3(n_479),
.B(n_475),
.Y(n_1516)
);

BUFx8_ASAP7_75t_L g1517 ( 
.A(n_1426),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1453),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1399),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1410),
.Y(n_1520)
);

NOR2xp67_ASAP7_75t_SL g1521 ( 
.A(n_1386),
.B(n_33),
.Y(n_1521)
);

BUFx4_ASAP7_75t_R g1522 ( 
.A(n_1360),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1394),
.A2(n_482),
.B(n_481),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1409),
.A2(n_1414),
.B(n_1413),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1424),
.A2(n_1430),
.B(n_1371),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1431),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1370),
.A2(n_484),
.B(n_483),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1389),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1457),
.B(n_486),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1359),
.A2(n_488),
.B(n_487),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1382),
.A2(n_490),
.B(n_489),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1425),
.A2(n_492),
.B(n_491),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1395),
.A2(n_1374),
.B(n_1417),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1420),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1440),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1433),
.B(n_36),
.Y(n_1536)
);

AOI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1444),
.A2(n_494),
.B(n_493),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1385),
.A2(n_497),
.B(n_496),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1449),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.C(n_40),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1411),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1432),
.A2(n_500),
.B(n_498),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1442),
.A2(n_502),
.B(n_501),
.Y(n_1542)
);

AOI22x1_ASAP7_75t_L g1543 ( 
.A1(n_1415),
.A2(n_1419),
.B1(n_1438),
.B2(n_1435),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1367),
.B(n_37),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1460),
.B(n_40),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1397),
.A2(n_505),
.B(n_503),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1462),
.A2(n_507),
.B(n_506),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1450),
.A2(n_511),
.B(n_510),
.Y(n_1548)
);

INVx8_ASAP7_75t_L g1549 ( 
.A(n_1368),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1447),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1408),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1454),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1458),
.A2(n_1416),
.B(n_1429),
.C(n_1436),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1400),
.B(n_513),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1448),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.C(n_47),
.Y(n_1555)
);

INVx4_ASAP7_75t_SL g1556 ( 
.A(n_1461),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1437),
.B(n_1354),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1375),
.A2(n_515),
.B(n_514),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1426),
.B(n_44),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1461),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1379),
.A2(n_1372),
.B(n_1393),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1421),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1451),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1428),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1451),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1428),
.B(n_45),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1445),
.B(n_1402),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1445),
.B(n_516),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1402),
.B(n_46),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1384),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1361),
.B(n_48),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1361),
.Y(n_1572)
);

AOI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1362),
.A2(n_518),
.B(n_517),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1423),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1355),
.B(n_50),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1384),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1362),
.A2(n_522),
.B(n_520),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1361),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1380),
.B(n_523),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1362),
.A2(n_525),
.B(n_524),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1361),
.B(n_51),
.Y(n_1581)
);

AO31x2_ASAP7_75t_L g1582 ( 
.A1(n_1362),
.A2(n_527),
.A3(n_528),
.B(n_526),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1361),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1362),
.A2(n_530),
.B(n_529),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1401),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1578),
.Y(n_1586)
);

AO21x1_ASAP7_75t_L g1587 ( 
.A1(n_1551),
.A2(n_52),
.B(n_53),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1572),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1470),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1535),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1491),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1536),
.B(n_54),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1583),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1575),
.B(n_54),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1504),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1519),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1469),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1555),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1484),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1507),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1503),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1512),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1534),
.Y(n_1603)
);

INVx5_ASAP7_75t_SL g1604 ( 
.A(n_1579),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1499),
.B(n_56),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1581),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1479),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1484),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1576),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1468),
.B(n_57),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1566),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1576),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1569),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1471),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1487),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1550),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1559),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1511),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1563),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1465),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1545),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1467),
.A2(n_533),
.B(n_531),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1526),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1517),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1525),
.A2(n_535),
.B(n_534),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1477),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1520),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1557),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1565),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1482),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1567),
.A2(n_537),
.B(n_536),
.Y(n_1632)
);

O2A1O1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1553),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1490),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1481),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1585),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1473),
.B(n_63),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1496),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1495),
.B(n_65),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1496),
.Y(n_1640)
);

OAI221xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1574),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1516),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1570),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1532),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1474),
.B(n_67),
.Y(n_1645)
);

INVxp33_ASAP7_75t_L g1646 ( 
.A(n_1472),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1493),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1516),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1489),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1568),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1478),
.A2(n_539),
.B(n_538),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1480),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1529),
.B(n_540),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1544),
.B(n_69),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1580),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1514),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1564),
.A2(n_544),
.B(n_541),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1485),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1466),
.B(n_70),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1582),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1475),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1533),
.A2(n_546),
.B(n_545),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_R g1664 ( 
.A(n_1589),
.B(n_1608),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1607),
.B(n_1606),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1615),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1599),
.B(n_1505),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_R g1668 ( 
.A(n_1638),
.B(n_1549),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_R g1669 ( 
.A(n_1640),
.B(n_1579),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1620),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1634),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1609),
.B(n_1505),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1630),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_R g1675 ( 
.A(n_1636),
.B(n_1500),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1618),
.B(n_1475),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1592),
.B(n_1521),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1658),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1549),
.Y(n_1679)
);

XNOR2xp5_ASAP7_75t_L g1680 ( 
.A(n_1646),
.B(n_1492),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1647),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1628),
.B(n_1610),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1602),
.B(n_1497),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1617),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_R g1685 ( 
.A(n_1619),
.B(n_1509),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_R g1686 ( 
.A(n_1653),
.B(n_1524),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1637),
.B(n_1522),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_R g1688 ( 
.A(n_1653),
.B(n_1502),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1515),
.Y(n_1689)
);

INVx8_ASAP7_75t_L g1690 ( 
.A(n_1647),
.Y(n_1690)
);

CKINVDCx12_ASAP7_75t_R g1691 ( 
.A(n_1654),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_R g1692 ( 
.A(n_1659),
.B(n_1483),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1647),
.Y(n_1693)
);

BUFx10_ASAP7_75t_L g1694 ( 
.A(n_1613),
.Y(n_1694)
);

OR2x4_ASAP7_75t_L g1695 ( 
.A(n_1625),
.B(n_1488),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1603),
.B(n_1476),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1494),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1633),
.B(n_1501),
.Y(n_1698)
);

NAND2xp33_ASAP7_75t_R g1699 ( 
.A(n_1645),
.B(n_1577),
.Y(n_1699)
);

XOR2x2_ASAP7_75t_SL g1700 ( 
.A(n_1635),
.B(n_1518),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_R g1701 ( 
.A(n_1611),
.B(n_1542),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1643),
.B(n_1486),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1614),
.B(n_1612),
.Y(n_1703)
);

XNOR2xp5_ASAP7_75t_L g1704 ( 
.A(n_1594),
.B(n_1528),
.Y(n_1704)
);

BUFx10_ASAP7_75t_L g1705 ( 
.A(n_1616),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_R g1706 ( 
.A(n_1596),
.B(n_1509),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1591),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1605),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1666),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1676),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1703),
.B(n_1696),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1663),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1677),
.B(n_1639),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1678),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1708),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1671),
.B(n_1661),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1661),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1670),
.B(n_1630),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1681),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1690),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1679),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1674),
.B(n_1590),
.Y(n_1724)
);

OAI222xp33_ASAP7_75t_L g1725 ( 
.A1(n_1698),
.A2(n_1641),
.B1(n_1622),
.B2(n_1652),
.C1(n_1508),
.C2(n_1627),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1665),
.B(n_1590),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1682),
.B(n_1595),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1673),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1683),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1689),
.B(n_1624),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1709),
.B(n_1588),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1697),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1680),
.B(n_1593),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1707),
.B(n_1642),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1667),
.B(n_1601),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1672),
.B(n_1648),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1693),
.B(n_1600),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1697),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1690),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1693),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1692),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1687),
.B(n_1604),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_1597),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1705),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1698),
.A2(n_1587),
.B1(n_1539),
.B2(n_1554),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1694),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1691),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1686),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1704),
.A2(n_1598),
.B1(n_1530),
.B2(n_1513),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1702),
.B(n_1621),
.Y(n_1752)
);

NOR2xp67_ASAP7_75t_L g1753 ( 
.A(n_1675),
.B(n_1644),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1685),
.B(n_1604),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1695),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1701),
.B(n_1631),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1699),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1711),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1720),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1757),
.B(n_1660),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1733),
.B(n_1664),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1747),
.B(n_1560),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1713),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1719),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1756),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1562),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1741),
.B(n_1632),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1755),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1744),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1713),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

AOI222xp33_ASAP7_75t_L g1772 ( 
.A1(n_1750),
.A2(n_1509),
.B1(n_1498),
.B2(n_1556),
.C1(n_1541),
.C2(n_95),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1734),
.B(n_1632),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1718),
.B(n_1668),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1710),
.B(n_1657),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1748),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1729),
.B(n_1657),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1714),
.B(n_1655),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1724),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1716),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1728),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1726),
.Y(n_1782)
);

OAI31xp33_ASAP7_75t_L g1783 ( 
.A1(n_1725),
.A2(n_1750),
.A3(n_1751),
.B(n_1745),
.Y(n_1783)
);

OAI31xp33_ASAP7_75t_L g1784 ( 
.A1(n_1738),
.A2(n_1688),
.A3(n_1669),
.B(n_1540),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1715),
.B(n_1749),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1736),
.B(n_1651),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1740),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1717),
.B(n_1651),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1723),
.B(n_1662),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1731),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1738),
.B(n_1626),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1752),
.A2(n_1543),
.B1(n_1561),
.B2(n_1558),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1753),
.A2(n_1538),
.B(n_1548),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1735),
.B(n_1623),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1727),
.B(n_1527),
.Y(n_1796)
);

INVx5_ASAP7_75t_L g1797 ( 
.A(n_1746),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1730),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1730),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1752),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1737),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1721),
.B(n_1531),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1740),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1746),
.Y(n_1804)
);

AO21x2_ASAP7_75t_L g1805 ( 
.A1(n_1755),
.A2(n_1584),
.B(n_1573),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1754),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1722),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1739),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1742),
.B(n_1547),
.Y(n_1809)
);

AOI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1750),
.A2(n_1546),
.B(n_1506),
.C(n_1523),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1712),
.B(n_71),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1740),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1751),
.A2(n_1510),
.B1(n_1537),
.B2(n_74),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1711),
.B(n_72),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1720),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1732),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1757),
.B(n_72),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1746),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1732),
.B(n_74),
.Y(n_1819)
);

NOR2xp67_ASAP7_75t_L g1820 ( 
.A(n_1741),
.B(n_75),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1757),
.B(n_76),
.Y(n_1821)
);

NAND2x1_ASAP7_75t_L g1822 ( 
.A(n_1753),
.B(n_76),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1757),
.B(n_77),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1711),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1720),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1763),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1770),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1780),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1798),
.B(n_77),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1800),
.B(n_78),
.Y(n_1830)
);

AND3x2_ASAP7_75t_L g1831 ( 
.A(n_1783),
.B(n_1804),
.C(n_1817),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1765),
.B(n_78),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1764),
.B(n_79),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1776),
.B(n_79),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1782),
.B(n_80),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1816),
.B(n_80),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1781),
.B(n_81),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1793),
.B(n_82),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1771),
.B(n_83),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1758),
.B(n_1824),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1775),
.B(n_83),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1799),
.B(n_84),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1759),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1779),
.B(n_85),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1815),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1825),
.B(n_1773),
.Y(n_1846)
);

INVxp67_ASAP7_75t_SL g1847 ( 
.A(n_1777),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1790),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1801),
.B(n_85),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1806),
.B(n_1774),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1767),
.B(n_1760),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1768),
.B(n_86),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1803),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1769),
.B(n_87),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1778),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1791),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1786),
.B(n_87),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1761),
.B(n_88),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1812),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1762),
.B(n_88),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1788),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1766),
.B(n_89),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1811),
.B(n_89),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1814),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1789),
.B(n_90),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1796),
.B(n_90),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1797),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1802),
.B(n_1821),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1823),
.B(n_91),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1795),
.B(n_1818),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1807),
.Y(n_1871)
);

NOR2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1822),
.B(n_91),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1808),
.B(n_92),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1787),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1784),
.B(n_92),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1797),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1818),
.B(n_1797),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1819),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1819),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1822),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1809),
.B(n_93),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1785),
.B(n_1820),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1805),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1792),
.B(n_1794),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1813),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1772),
.B(n_93),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1810),
.B(n_94),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1765),
.B(n_94),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1763),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1765),
.B(n_95),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1765),
.B(n_96),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1763),
.Y(n_1892)
);

NAND2x1p5_ASAP7_75t_L g1893 ( 
.A(n_1797),
.B(n_547),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1765),
.B(n_97),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1763),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1798),
.B(n_97),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1818),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1765),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1765),
.B(n_99),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1765),
.B(n_99),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1765),
.B(n_100),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1763),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1763),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1818),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1765),
.B(n_100),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1765),
.B(n_101),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1765),
.B(n_101),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1765),
.B(n_102),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1763),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1898),
.B(n_103),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1847),
.B(n_103),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1840),
.B(n_104),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1862),
.B(n_105),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1826),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1868),
.B(n_106),
.Y(n_1915)
);

OAI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1886),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.C(n_110),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1885),
.A2(n_112),
.B1(n_109),
.B2(n_111),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1875),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.C(n_114),
.Y(n_1918)
);

NAND2xp33_ASAP7_75t_SL g1919 ( 
.A(n_1872),
.B(n_113),
.Y(n_1919)
);

AO221x2_ASAP7_75t_L g1920 ( 
.A1(n_1834),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.C(n_117),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1882),
.B(n_115),
.Y(n_1921)
);

OAI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1880),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1841),
.Y(n_1923)
);

NOR2x1_ASAP7_75t_L g1924 ( 
.A(n_1877),
.B(n_118),
.Y(n_1924)
);

AO221x2_ASAP7_75t_L g1925 ( 
.A1(n_1878),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.C(n_122),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1861),
.B(n_120),
.Y(n_1926)
);

OAI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1863),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_124),
.Y(n_1927)
);

NOR4xp25_ASAP7_75t_SL g1928 ( 
.A(n_1876),
.B(n_125),
.C(n_123),
.D(n_124),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1884),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1831),
.B(n_128),
.Y(n_1930)
);

OAI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1866),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1893),
.B(n_129),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_SL g1933 ( 
.A1(n_1888),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1933)
);

NAND2xp33_ASAP7_75t_SL g1934 ( 
.A(n_1852),
.B(n_133),
.Y(n_1934)
);

NAND2xp33_ASAP7_75t_R g1935 ( 
.A(n_1897),
.B(n_133),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1871),
.B(n_134),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1851),
.B(n_134),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1859),
.Y(n_1938)
);

INVxp33_ASAP7_75t_L g1939 ( 
.A(n_1870),
.Y(n_1939)
);

NAND2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1905),
.B(n_136),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1856),
.B(n_137),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1828),
.B(n_138),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1832),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1864),
.B(n_139),
.Y(n_1944)
);

OAI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1867),
.A2(n_143),
.B1(n_139),
.B2(n_140),
.Y(n_1945)
);

CKINVDCx14_ASAP7_75t_R g1946 ( 
.A(n_1858),
.Y(n_1946)
);

OAI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1900),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.C(n_146),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1879),
.B(n_144),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1881),
.A2(n_1865),
.B1(n_1857),
.B2(n_1850),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1881),
.A2(n_148),
.B1(n_145),
.B2(n_147),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1869),
.B(n_147),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1843),
.B(n_1845),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1904),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1874),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1855),
.B(n_149),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1859),
.B(n_150),
.Y(n_1956)
);

INVxp33_ASAP7_75t_SL g1957 ( 
.A(n_1836),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1827),
.Y(n_1958)
);

OAI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1908),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_1959)
);

OAI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1849),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1848),
.B(n_154),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1835),
.B(n_155),
.Y(n_1962)
);

NOR2x1_ASAP7_75t_L g1963 ( 
.A(n_1890),
.B(n_1891),
.Y(n_1963)
);

OAI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1873),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1853),
.B(n_158),
.Y(n_1965)
);

NOR4xp25_ASAP7_75t_SL g1966 ( 
.A(n_1889),
.B(n_161),
.C(n_159),
.D(n_160),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1892),
.B(n_159),
.Y(n_1967)
);

NAND2xp33_ASAP7_75t_SL g1968 ( 
.A(n_1894),
.B(n_160),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1895),
.B(n_161),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1902),
.B(n_164),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1903),
.B(n_164),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1909),
.B(n_165),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1846),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1899),
.B(n_166),
.Y(n_1974)
);

AO221x2_ASAP7_75t_L g1975 ( 
.A1(n_1837),
.A2(n_1883),
.B1(n_1906),
.B2(n_1907),
.C(n_1901),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_SL g1976 ( 
.A1(n_1830),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1833),
.B(n_167),
.Y(n_1977)
);

A2O1A1Ixp33_ASAP7_75t_L g1978 ( 
.A1(n_1844),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1838),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1860),
.B(n_169),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1842),
.B(n_170),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1854),
.B(n_171),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1844),
.B(n_171),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_SL g1984 ( 
.A(n_1839),
.B(n_172),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1829),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_1985)
);

CKINVDCx8_ASAP7_75t_R g1986 ( 
.A(n_1896),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1897),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1887),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1887),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1897),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_SL g1991 ( 
.A(n_1872),
.B(n_180),
.Y(n_1991)
);

OAI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1887),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1887),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_1993)
);

OAI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1887),
.A2(n_188),
.B1(n_185),
.B2(n_187),
.C(n_189),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1898),
.B(n_188),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_SL g1996 ( 
.A(n_1872),
.B(n_190),
.Y(n_1996)
);

NOR4xp25_ASAP7_75t_SL g1997 ( 
.A(n_1876),
.B(n_192),
.C(n_190),
.D(n_191),
.Y(n_1997)
);

OAI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1886),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_R g1999 ( 
.A(n_1831),
.B(n_194),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1851),
.B(n_195),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1826),
.Y(n_2001)
);

OAI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1886),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_2002)
);

OAI22xp5_ASAP7_75t_SL g2003 ( 
.A1(n_1886),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1882),
.B(n_199),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1887),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1872),
.B(n_202),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1898),
.B(n_203),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1898),
.B(n_204),
.Y(n_2008)
);

OAI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1886),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1914),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1999),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_SL g2012 ( 
.A(n_1935),
.B(n_205),
.C(n_206),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1923),
.B(n_208),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1958),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2001),
.Y(n_2015)
);

AOI222xp33_ASAP7_75t_L g2016 ( 
.A1(n_2003),
.A2(n_210),
.B1(n_212),
.B2(n_208),
.C1(n_209),
.C2(n_211),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1937),
.B(n_209),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1953),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1930),
.B(n_210),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1943),
.B(n_212),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1952),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1957),
.B(n_213),
.Y(n_2022)
);

INVx1_ASAP7_75t_SL g2023 ( 
.A(n_1987),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1938),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1975),
.B(n_214),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2000),
.B(n_214),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1973),
.B(n_215),
.Y(n_2027)
);

INVx4_ASAP7_75t_L g2028 ( 
.A(n_1990),
.Y(n_2028)
);

INVxp67_ASAP7_75t_L g2029 ( 
.A(n_1921),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1975),
.B(n_215),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1986),
.Y(n_2031)
);

AND2x4_ASAP7_75t_SL g2032 ( 
.A(n_1949),
.B(n_216),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1979),
.B(n_216),
.Y(n_2033)
);

INVx1_ASAP7_75t_SL g2034 ( 
.A(n_1963),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_1924),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1946),
.B(n_217),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1911),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2004),
.B(n_217),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1965),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1915),
.B(n_218),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_1956),
.B(n_218),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1936),
.B(n_220),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1942),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1941),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_1918),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1926),
.B(n_221),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1912),
.B(n_222),
.Y(n_2047)
);

NAND2xp33_ASAP7_75t_L g2048 ( 
.A(n_1919),
.B(n_223),
.Y(n_2048)
);

HB1xp67_ASAP7_75t_L g2049 ( 
.A(n_1967),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1969),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1961),
.B(n_223),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1944),
.B(n_225),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1970),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1971),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1916),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1972),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1955),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1983),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1910),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1995),
.B(n_228),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2007),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1962),
.B(n_2008),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1913),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1981),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1948),
.B(n_229),
.Y(n_2065)
);

NAND2x1p5_ASAP7_75t_L g2066 ( 
.A(n_1933),
.B(n_229),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1982),
.B(n_232),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1920),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1977),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1974),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1920),
.B(n_1940),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1934),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1925),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1980),
.B(n_232),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_1968),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1925),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1950),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1991),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1951),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1932),
.B(n_233),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1931),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1959),
.B(n_234),
.Y(n_2082)
);

INVx1_ASAP7_75t_SL g2083 ( 
.A(n_1996),
.Y(n_2083)
);

INVx1_ASAP7_75t_SL g2084 ( 
.A(n_2006),
.Y(n_2084)
);

AO21x2_ASAP7_75t_L g2085 ( 
.A1(n_1922),
.A2(n_235),
.B(n_236),
.Y(n_2085)
);

INVxp67_ASAP7_75t_SL g2086 ( 
.A(n_1964),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1984),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1985),
.B(n_1988),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1989),
.B(n_235),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1960),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1947),
.Y(n_2091)
);

BUFx2_ASAP7_75t_SL g2092 ( 
.A(n_1954),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_R g2093 ( 
.A(n_1928),
.B(n_236),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1993),
.B(n_237),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2005),
.B(n_238),
.Y(n_2095)
);

OR2x6_ASAP7_75t_L g2096 ( 
.A(n_1976),
.B(n_238),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1998),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_1917),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2002),
.B(n_239),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1927),
.B(n_240),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2009),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1929),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1978),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1992),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_1994),
.B(n_240),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_1945),
.Y(n_2106)
);

OAI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_1966),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_1997),
.Y(n_2108)
);

AND3x1_ASAP7_75t_L g2109 ( 
.A(n_1930),
.B(n_241),
.C(n_242),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1914),
.Y(n_2110)
);

INVx1_ASAP7_75t_SL g2111 ( 
.A(n_1999),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_1930),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1923),
.B(n_244),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1938),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1938),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_1921),
.Y(n_2116)
);

INVx3_ASAP7_75t_L g2117 ( 
.A(n_1986),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1921),
.Y(n_2118)
);

INVxp67_ASAP7_75t_SL g2119 ( 
.A(n_1956),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1923),
.B(n_245),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_1938),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_1999),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_1938),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1923),
.B(n_247),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1914),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1939),
.B(n_248),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1923),
.B(n_249),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1923),
.B(n_250),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_1986),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1923),
.B(n_250),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1914),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1986),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1914),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1939),
.B(n_252),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1939),
.B(n_252),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1914),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1938),
.Y(n_2137)
);

INVxp67_ASAP7_75t_L g2138 ( 
.A(n_1921),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_1999),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1914),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1914),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_1986),
.Y(n_2142)
);

AO21x2_ASAP7_75t_L g2143 ( 
.A1(n_1999),
.A2(n_255),
.B(n_256),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1914),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_1999),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1938),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_1999),
.Y(n_2147)
);

NOR2x1_ASAP7_75t_L g2148 ( 
.A(n_1956),
.B(n_256),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1914),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_1937),
.B(n_257),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1939),
.B(n_258),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1914),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1939),
.B(n_258),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1914),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_1938),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_1937),
.B(n_259),
.Y(n_2156)
);

AOI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_1930),
.A2(n_259),
.B(n_260),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1986),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1939),
.B(n_260),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1938),
.B(n_261),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_1937),
.B(n_262),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1930),
.A2(n_265),
.B1(n_262),
.B2(n_264),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_1939),
.B(n_264),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2092),
.A2(n_2068),
.B1(n_2086),
.B2(n_2091),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2034),
.B(n_266),
.Y(n_2165)
);

NAND2x1_ASAP7_75t_L g2166 ( 
.A(n_2024),
.B(n_267),
.Y(n_2166)
);

OAI33xp33_ASAP7_75t_L g2167 ( 
.A1(n_2025),
.A2(n_2030),
.A3(n_2073),
.B1(n_2071),
.B2(n_2090),
.B3(n_2097),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2119),
.B(n_267),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2117),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2029),
.B(n_268),
.Y(n_2170)
);

OAI31xp33_ASAP7_75t_L g2171 ( 
.A1(n_2035),
.A2(n_270),
.A3(n_268),
.B(n_269),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2116),
.B(n_269),
.Y(n_2172)
);

OAI21xp33_ASAP7_75t_SL g2173 ( 
.A1(n_2118),
.A2(n_270),
.B(n_271),
.Y(n_2173)
);

INVx2_ASAP7_75t_SL g2174 ( 
.A(n_2031),
.Y(n_2174)
);

AOI21xp33_ASAP7_75t_L g2175 ( 
.A1(n_2100),
.A2(n_271),
.B(n_272),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2010),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2132),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2048),
.A2(n_272),
.B(n_273),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2138),
.B(n_273),
.Y(n_2179)
);

AOI21xp33_ASAP7_75t_L g2180 ( 
.A1(n_2016),
.A2(n_2104),
.B(n_2108),
.Y(n_2180)
);

AOI211xp5_ASAP7_75t_L g2181 ( 
.A1(n_2019),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2014),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2015),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2012),
.A2(n_276),
.B(n_277),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2110),
.Y(n_2185)
);

OAI221xp5_ASAP7_75t_L g2186 ( 
.A1(n_2122),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.C(n_280),
.Y(n_2186)
);

OAI21xp33_ASAP7_75t_L g2187 ( 
.A1(n_2045),
.A2(n_278),
.B(n_281),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2063),
.B(n_281),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2125),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2098),
.B(n_282),
.Y(n_2190)
);

INVxp67_ASAP7_75t_SL g2191 ( 
.A(n_2087),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2131),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_2158),
.B(n_283),
.Y(n_2193)
);

AOI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_2103),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2133),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2136),
.Y(n_2196)
);

AOI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2082),
.A2(n_285),
.B(n_287),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_2011),
.B(n_287),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2058),
.B(n_288),
.Y(n_2199)
);

AOI21xp33_ASAP7_75t_L g2200 ( 
.A1(n_2102),
.A2(n_289),
.B(n_290),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2140),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2059),
.B(n_289),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2076),
.B(n_290),
.Y(n_2203)
);

INVx1_ASAP7_75t_SL g2204 ( 
.A(n_2111),
.Y(n_2204)
);

OAI32xp33_ASAP7_75t_L g2205 ( 
.A1(n_2066),
.A2(n_294),
.A3(n_292),
.B1(n_293),
.B2(n_295),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2064),
.B(n_292),
.Y(n_2206)
);

AOI322xp5_ASAP7_75t_L g2207 ( 
.A1(n_2088),
.A2(n_293),
.A3(n_294),
.B1(n_295),
.B2(n_296),
.C1(n_297),
.C2(n_298),
.Y(n_2207)
);

INVxp67_ASAP7_75t_L g2208 ( 
.A(n_2143),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2103),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2209)
);

OAI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_2157),
.A2(n_299),
.B(n_300),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2069),
.B(n_300),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2129),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2077),
.B(n_301),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2079),
.B(n_301),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2044),
.B(n_303),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2141),
.Y(n_2216)
);

AOI222xp33_ASAP7_75t_L g2217 ( 
.A1(n_2094),
.A2(n_306),
.B1(n_308),
.B2(n_304),
.C1(n_305),
.C2(n_307),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2109),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_2218)
);

INVx1_ASAP7_75t_SL g2219 ( 
.A(n_2139),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2096),
.A2(n_307),
.B(n_308),
.Y(n_2220)
);

INVx1_ASAP7_75t_SL g2221 ( 
.A(n_2145),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2096),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2049),
.B(n_309),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2070),
.B(n_310),
.Y(n_2224)
);

OAI32xp33_ASAP7_75t_L g2225 ( 
.A1(n_2075),
.A2(n_313),
.A3(n_311),
.B1(n_312),
.B2(n_314),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2114),
.B(n_312),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_SL g2227 ( 
.A(n_2036),
.B(n_313),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2043),
.B(n_314),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2115),
.B(n_315),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2101),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2144),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2147),
.B(n_316),
.Y(n_2232)
);

BUFx2_ASAP7_75t_SL g2233 ( 
.A(n_2142),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2041),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2149),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2137),
.B(n_318),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2152),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2148),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2154),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_2121),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2021),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2056),
.B(n_318),
.Y(n_2242)
);

INVx1_ASAP7_75t_SL g2243 ( 
.A(n_2078),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2146),
.B(n_319),
.Y(n_2244)
);

OAI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2072),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2083),
.B(n_320),
.Y(n_2246)
);

AOI21xp33_ASAP7_75t_L g2247 ( 
.A1(n_2093),
.A2(n_2105),
.B(n_2084),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_L g2248 ( 
.A(n_2028),
.B(n_2106),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2123),
.Y(n_2249)
);

NAND4xp25_ASAP7_75t_L g2250 ( 
.A(n_2055),
.B(n_323),
.C(n_321),
.D(n_322),
.Y(n_2250)
);

AOI22xp33_ASAP7_75t_L g2251 ( 
.A1(n_2081),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2155),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2061),
.B(n_324),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2037),
.B(n_325),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2018),
.B(n_325),
.Y(n_2255)
);

XNOR2xp5_ASAP7_75t_L g2256 ( 
.A(n_2023),
.B(n_326),
.Y(n_2256)
);

NAND3xp33_ASAP7_75t_SL g2257 ( 
.A(n_2112),
.B(n_327),
.C(n_328),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2039),
.Y(n_2258)
);

INVxp67_ASAP7_75t_L g2259 ( 
.A(n_2160),
.Y(n_2259)
);

XOR2xp5_ASAP7_75t_L g2260 ( 
.A(n_2162),
.B(n_2099),
.Y(n_2260)
);

AOI221xp5_ASAP7_75t_L g2261 ( 
.A1(n_2089),
.A2(n_2095),
.B1(n_2107),
.B2(n_2020),
.C(n_2113),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2050),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2053),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2054),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2057),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2062),
.B(n_2160),
.Y(n_2266)
);

INVxp67_ASAP7_75t_L g2267 ( 
.A(n_2022),
.Y(n_2267)
);

INVx1_ASAP7_75t_SL g2268 ( 
.A(n_2032),
.Y(n_2268)
);

INVx1_ASAP7_75t_SL g2269 ( 
.A(n_2080),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2033),
.Y(n_2270)
);

AOI21xp33_ASAP7_75t_SL g2271 ( 
.A1(n_2085),
.A2(n_556),
.B(n_557),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2046),
.B(n_2126),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_2013),
.B(n_558),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2046),
.B(n_689),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2240),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2243),
.B(n_2249),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2176),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2269),
.B(n_2120),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2182),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2252),
.B(n_2124),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2183),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2234),
.B(n_2027),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2238),
.B(n_2038),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2208),
.B(n_2052),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2185),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2169),
.B(n_2134),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_2180),
.A2(n_2067),
.B1(n_2074),
.B2(n_2135),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2204),
.B(n_2047),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2233),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2189),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2174),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2212),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2219),
.B(n_2040),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2221),
.B(n_2151),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_2167),
.A2(n_2159),
.B1(n_2163),
.B2(n_2153),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2177),
.B(n_2065),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2192),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2191),
.B(n_2017),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2164),
.B(n_2127),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2195),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2259),
.B(n_2026),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2247),
.B(n_2128),
.Y(n_2302)
);

NOR2x1_ASAP7_75t_L g2303 ( 
.A(n_2165),
.B(n_2166),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2267),
.B(n_2130),
.Y(n_2304)
);

INVx1_ASAP7_75t_SL g2305 ( 
.A(n_2227),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2248),
.B(n_2150),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_2266),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2271),
.B(n_2156),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2268),
.B(n_2161),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2270),
.B(n_2042),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2272),
.B(n_2051),
.Y(n_2311)
);

INVx1_ASAP7_75t_SL g2312 ( 
.A(n_2202),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2196),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2260),
.B(n_2060),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2213),
.B(n_2214),
.Y(n_2315)
);

AOI222xp33_ASAP7_75t_L g2316 ( 
.A1(n_2257),
.A2(n_565),
.B1(n_566),
.B2(n_567),
.C1(n_568),
.C2(n_570),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2226),
.B(n_571),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2261),
.B(n_573),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2201),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2224),
.B(n_574),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2197),
.B(n_577),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2216),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2231),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2235),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2173),
.B(n_2223),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2229),
.B(n_578),
.Y(n_2326)
);

NAND2x1_ASAP7_75t_L g2327 ( 
.A(n_2237),
.B(n_580),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2239),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2173),
.B(n_2168),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2236),
.B(n_581),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2206),
.B(n_582),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2244),
.B(n_583),
.Y(n_2332)
);

INVx1_ASAP7_75t_SL g2333 ( 
.A(n_2255),
.Y(n_2333)
);

OAI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2218),
.A2(n_2230),
.B1(n_2181),
.B2(n_2184),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2275),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2301),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2276),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2277),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2279),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2289),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2303),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2281),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2285),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2290),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2305),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2297),
.Y(n_2346)
);

INVx5_ASAP7_75t_L g2347 ( 
.A(n_2291),
.Y(n_2347)
);

NAND2xp33_ASAP7_75t_L g2348 ( 
.A(n_2333),
.B(n_2245),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2300),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2296),
.Y(n_2350)
);

INVx3_ASAP7_75t_SL g2351 ( 
.A(n_2317),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2313),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2312),
.Y(n_2353)
);

INVx8_ASAP7_75t_L g2354 ( 
.A(n_2326),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2325),
.B(n_2203),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2319),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2322),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2323),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2324),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2328),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2286),
.Y(n_2361)
);

BUFx2_ASAP7_75t_L g2362 ( 
.A(n_2298),
.Y(n_2362)
);

HB1xp67_ASAP7_75t_L g2363 ( 
.A(n_2309),
.Y(n_2363)
);

INVx1_ASAP7_75t_SL g2364 ( 
.A(n_2306),
.Y(n_2364)
);

HB1xp67_ASAP7_75t_L g2365 ( 
.A(n_2288),
.Y(n_2365)
);

INVxp67_ASAP7_75t_L g2366 ( 
.A(n_2283),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2341),
.A2(n_2287),
.B1(n_2334),
.B2(n_2295),
.Y(n_2367)
);

NAND3xp33_ASAP7_75t_L g2368 ( 
.A(n_2348),
.B(n_2171),
.C(n_2207),
.Y(n_2368)
);

NOR2x1_ASAP7_75t_L g2369 ( 
.A(n_2340),
.B(n_2318),
.Y(n_2369)
);

NOR3xp33_ASAP7_75t_L g2370 ( 
.A(n_2355),
.B(n_2302),
.C(n_2284),
.Y(n_2370)
);

AOI211xp5_ASAP7_75t_L g2371 ( 
.A1(n_2345),
.A2(n_2222),
.B(n_2205),
.C(n_2175),
.Y(n_2371)
);

NAND5xp2_ASAP7_75t_L g2372 ( 
.A(n_2337),
.B(n_2336),
.C(n_2366),
.D(n_2362),
.E(n_2335),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2363),
.A2(n_2314),
.B(n_2329),
.Y(n_2373)
);

NOR3xp33_ASAP7_75t_L g2374 ( 
.A(n_2353),
.B(n_2365),
.C(n_2364),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2361),
.Y(n_2375)
);

AOI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2354),
.A2(n_2299),
.B(n_2308),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2347),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2347),
.B(n_2286),
.Y(n_2378)
);

NAND3xp33_ASAP7_75t_L g2379 ( 
.A(n_2350),
.B(n_2217),
.C(n_2220),
.Y(n_2379)
);

OAI21xp5_ASAP7_75t_SL g2380 ( 
.A1(n_2340),
.A2(n_2210),
.B(n_2178),
.Y(n_2380)
);

AND4x1_ASAP7_75t_L g2381 ( 
.A(n_2360),
.B(n_2246),
.C(n_2304),
.D(n_2316),
.Y(n_2381)
);

NOR3x1_ASAP7_75t_L g2382 ( 
.A(n_2338),
.B(n_2294),
.C(n_2282),
.Y(n_2382)
);

NOR3xp33_ASAP7_75t_L g2383 ( 
.A(n_2339),
.B(n_2307),
.C(n_2292),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2351),
.B(n_2293),
.Y(n_2384)
);

O2A1O1Ixp5_ASAP7_75t_L g2385 ( 
.A1(n_2378),
.A2(n_2343),
.B(n_2344),
.C(n_2342),
.Y(n_2385)
);

OA22x2_ASAP7_75t_L g2386 ( 
.A1(n_2380),
.A2(n_2262),
.B1(n_2263),
.B2(n_2258),
.Y(n_2386)
);

NAND4xp25_ASAP7_75t_L g2387 ( 
.A(n_2372),
.B(n_2315),
.C(n_2280),
.D(n_2278),
.Y(n_2387)
);

OAI211xp5_ASAP7_75t_SL g2388 ( 
.A1(n_2367),
.A2(n_2349),
.B(n_2352),
.C(n_2346),
.Y(n_2388)
);

AOI221xp5_ASAP7_75t_L g2389 ( 
.A1(n_2368),
.A2(n_2358),
.B1(n_2359),
.B2(n_2357),
.C(n_2356),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2371),
.A2(n_2251),
.B1(n_2311),
.B2(n_2209),
.Y(n_2390)
);

AOI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2370),
.A2(n_2225),
.B1(n_2200),
.B2(n_2250),
.C(n_2187),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2373),
.A2(n_2179),
.B1(n_2172),
.B2(n_2170),
.C(n_2310),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2377),
.B(n_2374),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2385),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2393),
.Y(n_2395)
);

NOR2x1_ASAP7_75t_L g2396 ( 
.A(n_2387),
.B(n_2384),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2386),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2391),
.B(n_2376),
.Y(n_2398)
);

NOR2x1_ASAP7_75t_L g2399 ( 
.A(n_2388),
.B(n_2379),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2392),
.B(n_2375),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2389),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2394),
.B(n_2383),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_R g2403 ( 
.A(n_2395),
.B(n_2198),
.Y(n_2403)
);

NAND2xp33_ASAP7_75t_SL g2404 ( 
.A(n_2397),
.B(n_2327),
.Y(n_2404)
);

NAND2xp33_ASAP7_75t_SL g2405 ( 
.A(n_2400),
.B(n_2390),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2396),
.B(n_2382),
.Y(n_2406)
);

AOI211x1_ASAP7_75t_L g2407 ( 
.A1(n_2406),
.A2(n_2381),
.B(n_2398),
.C(n_2401),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2405),
.A2(n_2399),
.B1(n_2369),
.B2(n_2354),
.Y(n_2408)
);

NAND4xp25_ASAP7_75t_L g2409 ( 
.A(n_2407),
.B(n_2402),
.C(n_2404),
.D(n_2232),
.Y(n_2409)
);

XNOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2409),
.B(n_2408),
.Y(n_2410)
);

AOI31xp33_ASAP7_75t_L g2411 ( 
.A1(n_2410),
.A2(n_2403),
.A3(n_2256),
.B(n_2190),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2410),
.A2(n_2264),
.B1(n_2265),
.B2(n_2321),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2412),
.A2(n_2215),
.B1(n_2254),
.B2(n_2253),
.Y(n_2413)
);

OAI322xp33_ASAP7_75t_L g2414 ( 
.A1(n_2411),
.A2(n_2193),
.A3(n_2320),
.B1(n_2242),
.B2(n_2228),
.C1(n_2211),
.C2(n_2331),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2414),
.A2(n_2199),
.B(n_2188),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2413),
.Y(n_2416)
);

BUFx2_ASAP7_75t_L g2417 ( 
.A(n_2416),
.Y(n_2417)
);

XOR2xp5_ASAP7_75t_L g2418 ( 
.A(n_2415),
.B(n_2194),
.Y(n_2418)
);

AOI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2418),
.A2(n_2273),
.B1(n_2332),
.B2(n_2330),
.C(n_2241),
.Y(n_2419)
);

AOI211xp5_ASAP7_75t_L g2420 ( 
.A1(n_2419),
.A2(n_2417),
.B(n_2274),
.C(n_2186),
.Y(n_2420)
);


endmodule