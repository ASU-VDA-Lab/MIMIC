module real_jpeg_17994_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_0),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_148),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_0),
.B(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_2),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_3),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_3),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_3),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_3),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_3),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_3),
.B(n_333),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_4),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_74),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_4),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_5),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_9),
.B1(n_113),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_5),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_6),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_6),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_6),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_6),
.B(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_9),
.B(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_11),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_12),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_13),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_13),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_13),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_13),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_13),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_13),
.B(n_246),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_13),
.B(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_14),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_14),
.Y(n_318)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_15),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_206),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_205),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_156),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_20),
.B(n_156),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.C(n_121),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_21),
.B(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_23),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_26),
.B(n_35),
.C(n_36),
.Y(n_194)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_54),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_43),
.A2(n_49),
.B(n_54),
.C(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_48),
.B(n_53),
.Y(n_176)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_52),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_63),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_63),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_55),
.Y(n_124)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_63),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_65),
.B(n_158),
.C(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_80),
.C(n_87),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_66),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_71),
.C(n_77),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_69),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_80),
.A2(n_81),
.B1(n_87),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_86),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_87),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.C(n_94),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_88),
.A2(n_94),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_90),
.B(n_219),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_92),
.Y(n_302)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_94),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_96),
.B(n_121),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_111),
.C(n_120),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_102),
.C(n_105),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_108),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_103),
.Y(n_252)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_105),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_107),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_108),
.B(n_140),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_120),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_127),
.B(n_134),
.Y(n_126)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_119),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_138),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_122),
.B(n_126),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_128),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_128),
.B(n_228),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_137),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_138),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.C(n_150),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_139),
.B(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_144),
.A2(n_145),
.B1(n_150),
.B2(n_151),
.Y(n_241)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_179),
.B2(n_180),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_174),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_203),
.B2(n_204),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_201),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_201),
.B(n_250),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_232),
.B(n_348),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_208),
.B(n_210),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_217),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_223),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_230),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_230),
.Y(n_291)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_256),
.B(n_347),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_253),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_236),
.B(n_253),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_237),
.A2(n_238),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_240),
.B(n_242),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.C(n_249),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_249),
.B(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_341),
.B(n_346),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_295),
.B(n_340),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_287),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_259),
.B(n_287),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_276),
.C(n_285),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_260),
.A2(n_261),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_269),
.C(n_271),
.Y(n_289)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_285),
.B1(n_286),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_290),
.C(n_292),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_309),
.B(n_339),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_305),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_297),
.B(n_305),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.C(n_303),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_303),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_306),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_324),
.B(n_338),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_321),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_311),
.B(n_321),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_319),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_328),
.B(n_337),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_326),
.B(n_327),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_342),
.B(n_343),
.Y(n_346)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);


endmodule