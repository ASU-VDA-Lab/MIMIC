module fake_jpeg_10627_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_20),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_5),
.B1(n_6),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_21),
.B1(n_13),
.B2(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_6),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_12),
.B1(n_9),
.B2(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_29),
.B1(n_10),
.B2(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_1),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_7),
.B(n_10),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_12),
.B1(n_20),
.B2(n_10),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_7),
.C(n_10),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_16),
.C(n_15),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_26),
.C(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_35),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_42),
.B(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_41),
.Y(n_48)
);

XNOR2x1_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_26),
.Y(n_47)
);

OAI221xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.C(n_28),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_49),
.B(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_4),
.B1(n_38),
.B2(n_45),
.Y(n_52)
);


endmodule