module fake_jpeg_3405_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_8),
.B1(n_11),
.B2(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_9),
.B(n_3),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_20),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_22),
.B(n_16),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_18),
.B1(n_17),
.B2(n_12),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp67_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_27),
.C(n_24),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_22),
.B(n_10),
.C(n_12),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_41),
.C(n_33),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_34),
.B1(n_27),
.B2(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_41),
.C(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_42),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_26),
.Y(n_48)
);

AOI211xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_38),
.B(n_14),
.C(n_4),
.Y(n_49)
);

NOR4xp25_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_4),
.C(n_14),
.D(n_32),
.Y(n_50)
);


endmodule