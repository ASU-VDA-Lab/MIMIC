module fake_jpeg_27733_n_275 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_51),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_27),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_23),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_38),
.B1(n_20),
.B2(n_22),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_64),
.B1(n_2),
.B2(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_38),
.B1(n_56),
.B2(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_36),
.B1(n_24),
.B2(n_33),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_76),
.B1(n_79),
.B2(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_73),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_89),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_22),
.B1(n_24),
.B2(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_29),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_73),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_31),
.B1(n_25),
.B2(n_23),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_30),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_99),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_101),
.Y(n_129)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_35),
.C(n_30),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_18),
.B1(n_30),
.B2(n_3),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_116),
.B1(n_88),
.B2(n_89),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_59),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_1),
.C(n_2),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_59),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_118),
.B1(n_103),
.B2(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_74),
.B1(n_85),
.B2(n_83),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_82),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_60),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_9),
.Y(n_138)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_121),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_14),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_138),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_97),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_91),
.B(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_146),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_105),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_138),
.B(n_133),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_145),
.B1(n_150),
.B2(n_119),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_99),
.B1(n_95),
.B2(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_93),
.B(n_81),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_92),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_156),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_123),
.B1(n_95),
.B2(n_101),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_159),
.B1(n_161),
.B2(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_132),
.B1(n_148),
.B2(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_116),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_165),
.B(n_177),
.Y(n_183)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_173),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_83),
.B1(n_85),
.B2(n_74),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_168),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_175),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_81),
.B(n_124),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_174),
.B(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_109),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_108),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_135),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_143),
.B1(n_142),
.B2(n_128),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_172),
.B1(n_98),
.B2(n_175),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_94),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_136),
.B1(n_135),
.B2(n_134),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_136),
.B(n_144),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_154),
.B(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_199),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_9),
.B(n_10),
.Y(n_198)
);

OAI322xp33_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_160),
.A3(n_174),
.B1(n_191),
.B2(n_197),
.C1(n_199),
.C2(n_186),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_134),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_167),
.B(n_11),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_177),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_161),
.C(n_157),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_159),
.C(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_215),
.C(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_163),
.B1(n_155),
.B2(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_183),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_170),
.C(n_165),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_153),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_219),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_201),
.B(n_190),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_220),
.B1(n_194),
.B2(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_172),
.C(n_166),
.Y(n_222)
);

OAI321xp33_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_186),
.A3(n_190),
.B1(n_192),
.B2(n_200),
.C(n_182),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_211),
.B1(n_222),
.B2(n_215),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_219),
.B(n_104),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_201),
.B1(n_184),
.B2(n_188),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_227),
.B1(n_212),
.B2(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_187),
.B1(n_181),
.B2(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_15),
.Y(n_246)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

NAND4xp25_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_204),
.C(n_181),
.D(n_183),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_246),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_217),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_245),
.B(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_237),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_234),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_11),
.B(n_13),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_11),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_228),
.B(n_226),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_255),
.B(n_245),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_256),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_68),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_229),
.B(n_236),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_238),
.C(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_252),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_239),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_262),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_236),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_265),
.B(n_257),
.C(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_235),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_235),
.B(n_248),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_263),
.B(n_233),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.C(n_233),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_256),
.C(n_267),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_272),
.C(n_68),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_68),
.Y(n_275)
);


endmodule