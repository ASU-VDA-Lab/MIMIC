module fake_netlist_6_2610_n_1023 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1023);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1023;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_880;
wire n_981;
wire n_476;
wire n_792;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_267;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_63),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_138),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_56),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_13),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_76),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_132),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_79),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_75),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_36),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_41),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_46),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_176),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_86),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_101),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_127),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_77),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_83),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_93),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_16),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_182),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_196),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_34),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_22),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_116),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_44),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_130),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_12),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_59),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_43),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_58),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_51),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_62),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_38),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_137),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_109),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_142),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_119),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_164),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_87),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_158),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_193),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_162),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_139),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_186),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_61),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_60),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_194),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_104),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_39),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_103),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_180),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_17),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_50),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_73),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_128),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_135),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_110),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_24),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_224),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_225),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_238),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_239),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_223),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_250),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_228),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_230),
.B(n_0),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_203),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_228),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_252),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_254),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_230),
.B(n_0),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_216),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_256),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_220),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_258),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_254),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_212),
.B(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_264),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_212),
.B(n_1),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_262),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_281),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_202),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_282),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_242),
.B(n_2),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_208),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_273),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_273),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_204),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_206),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_209),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_214),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_210),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_265),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_338),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_338),
.B(n_265),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_205),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_285),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_340),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_265),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_339),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_285),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_293),
.A2(n_248),
.B(n_222),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_305),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_331),
.B(n_207),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_337),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_292),
.B(n_222),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_337),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_R g378 ( 
.A(n_298),
.B(n_217),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_309),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_298),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_299),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_290),
.B(n_248),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_287),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_287),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_299),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_311),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_300),
.B(n_213),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_R g393 ( 
.A(n_300),
.B(n_218),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_SL g395 ( 
.A(n_301),
.B(n_247),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_324),
.B(n_215),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_304),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_R g398 ( 
.A(n_310),
.B(n_219),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_344),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_378),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_314),
.Y(n_408)
);

NAND2x1p5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_221),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_314),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_255),
.B1(n_277),
.B2(n_205),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_316),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_393),
.B(n_316),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_229),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_327),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_327),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_328),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_379),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_398),
.B(n_328),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_375),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_364),
.B(n_330),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_351),
.B(n_330),
.Y(n_436)
);

CKINVDCx8_ASAP7_75t_R g437 ( 
.A(n_370),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_351),
.B(n_231),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_359),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_375),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_383),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_382),
.B(n_308),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_364),
.B(n_323),
.Y(n_447)
);

BUFx4_ASAP7_75t_L g448 ( 
.A(n_345),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_227),
.C(n_226),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_377),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_388),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_317),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

BUFx8_ASAP7_75t_SL g457 ( 
.A(n_377),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_346),
.Y(n_458)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

CKINVDCx8_ASAP7_75t_R g462 ( 
.A(n_390),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_355),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_364),
.B(n_232),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_233),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_360),
.B(n_371),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_385),
.A2(n_205),
.B1(n_255),
.B2(n_277),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_353),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_235),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_385),
.A2(n_396),
.B1(n_344),
.B2(n_355),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_360),
.B(n_237),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_371),
.B(n_240),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_402),
.B(n_401),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_366),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_385),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_357),
.B(n_335),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_380),
.B(n_241),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_410),
.A2(n_381),
.B1(n_386),
.B2(n_380),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_476),
.B(n_396),
.Y(n_481)
);

CKINVDCx11_ASAP7_75t_R g482 ( 
.A(n_437),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_408),
.B(n_394),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_460),
.A2(n_459),
.B1(n_467),
.B2(n_409),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_475),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_396),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_SL g490 ( 
.A(n_432),
.B(n_321),
.C(n_320),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_425),
.B(n_400),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_403),
.B(n_400),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_459),
.A2(n_349),
.B(n_347),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_445),
.B(n_352),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_444),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_381),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_403),
.B(n_347),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_405),
.B(n_357),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_415),
.B(n_386),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_470),
.B(n_404),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_415),
.B(n_423),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_446),
.B(n_354),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_404),
.B(n_397),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_354),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_428),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_454),
.B(n_356),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_407),
.B(n_356),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_458),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_423),
.B(n_426),
.Y(n_513)
);

NAND2x1_ASAP7_75t_L g514 ( 
.A(n_420),
.B(n_350),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_455),
.A2(n_399),
.B1(n_397),
.B2(n_348),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_234),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_440),
.B(n_399),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_426),
.A2(n_336),
.B1(n_243),
.B2(n_271),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_236),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_406),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_246),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_436),
.B(n_249),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_434),
.B(n_255),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_459),
.A2(n_260),
.B1(n_261),
.B2(n_269),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_436),
.A2(n_268),
.B1(n_253),
.B2(n_257),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_447),
.B(n_259),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_L g530 ( 
.A(n_449),
.B(n_266),
.C(n_263),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_465),
.B(n_276),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_469),
.B(n_283),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_409),
.B(n_255),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_438),
.B(n_284),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_438),
.B(n_358),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_444),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_438),
.B(n_358),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_409),
.B(n_277),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_442),
.B(n_270),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_432),
.A2(n_289),
.B1(n_247),
.B2(n_267),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_433),
.B(n_471),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_442),
.B(n_272),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_434),
.A2(n_286),
.B1(n_278),
.B2(n_251),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_452),
.B(n_277),
.Y(n_547)
);

BUFx6f_ASAP7_75t_SL g548 ( 
.A(n_443),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_422),
.B(n_418),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_413),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_411),
.B(n_440),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_422),
.B(n_251),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_452),
.B(n_350),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_451),
.B(n_350),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_464),
.A2(n_251),
.B1(n_289),
.B2(n_267),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_451),
.B(n_350),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_422),
.A2(n_245),
.B1(n_350),
.B2(n_4),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_451),
.B(n_350),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_444),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_472),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_488),
.B(n_456),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_479),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_519),
.B(n_485),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_SL g567 ( 
.A(n_543),
.B(n_450),
.C(n_441),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_527),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_484),
.B(n_474),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_461),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_524),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_491),
.B(n_461),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_482),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_483),
.B(n_461),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_524),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_517),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_525),
.B(n_418),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_SL g580 ( 
.A(n_490),
.B(n_450),
.C(n_441),
.Y(n_580)
);

AO22x1_ASAP7_75t_L g581 ( 
.A1(n_495),
.A2(n_448),
.B1(n_466),
.B2(n_443),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_519),
.B(n_416),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_485),
.B(n_507),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_495),
.B(n_443),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_548),
.B(n_437),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_507),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_500),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_509),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_539),
.Y(n_590)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_500),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_429),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_483),
.B(n_444),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_513),
.A2(n_478),
.B1(n_473),
.B2(n_420),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_548),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

AOI221xp5_ASAP7_75t_L g597 ( 
.A1(n_503),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.C(n_6),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_487),
.B(n_462),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_513),
.B(n_444),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_503),
.A2(n_473),
.B1(n_420),
.B2(n_430),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_493),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_512),
.B(n_473),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_SL g603 ( 
.A(n_502),
.B(n_448),
.C(n_457),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_521),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_534),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_501),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_525),
.B(n_544),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_SL g609 ( 
.A(n_498),
.B(n_457),
.C(n_462),
.Y(n_609)
);

OR2x2_ASAP7_75t_SL g610 ( 
.A(n_504),
.B(n_3),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_547),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_498),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_558),
.B(n_412),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_558),
.B(n_412),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_562),
.B(n_412),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_538),
.B(n_540),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_480),
.B(n_412),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_492),
.B(n_412),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_418),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_544),
.A2(n_439),
.B1(n_431),
.B2(n_430),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_515),
.B(n_427),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_506),
.B(n_5),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_537),
.Y(n_628)
);

BUFx12f_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_608),
.A2(n_529),
.B(n_546),
.C(n_555),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_596),
.A2(n_552),
.B(n_541),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_608),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_601),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_596),
.A2(n_552),
.B(n_541),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_563),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_618),
.B(n_551),
.Y(n_637)
);

AO21x1_ASAP7_75t_L g638 ( 
.A1(n_593),
.A2(n_526),
.B(n_535),
.Y(n_638)
);

AO31x2_ASAP7_75t_L g639 ( 
.A1(n_571),
.A2(n_532),
.A3(n_531),
.B(n_516),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_571),
.A2(n_535),
.B(n_494),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_592),
.B(n_481),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_569),
.A2(n_604),
.B(n_578),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_613),
.A2(n_553),
.B(n_508),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_615),
.A2(n_616),
.B1(n_570),
.B2(n_597),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_599),
.B(n_520),
.Y(n_645)
);

OAI21x1_ASAP7_75t_SL g646 ( 
.A1(n_615),
.A2(n_536),
.B(n_489),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_599),
.B(n_550),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_573),
.B(n_550),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_573),
.B(n_499),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_612),
.B(n_518),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_575),
.B(n_511),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_530),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

NOR2x1_ASAP7_75t_L g654 ( 
.A(n_584),
.B(n_523),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_628),
.A2(n_510),
.B(n_505),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_587),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_566),
.B(n_497),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_624),
.A2(n_557),
.B(n_554),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_623),
.A2(n_560),
.B(n_549),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_606),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_623),
.A2(n_549),
.B(n_514),
.Y(n_661)
);

OAI21x1_ASAP7_75t_SL g662 ( 
.A1(n_616),
.A2(n_545),
.B(n_542),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_570),
.A2(n_561),
.B(n_528),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_593),
.A2(n_547),
.B(n_430),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_605),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_597),
.A2(n_439),
.B1(n_431),
.B2(n_430),
.Y(n_666)
);

AOI211x1_ASAP7_75t_L g667 ( 
.A1(n_568),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_575),
.A2(n_579),
.B(n_621),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_625),
.A2(n_439),
.B(n_431),
.C(n_430),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_598),
.B(n_7),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_625),
.A2(n_439),
.B(n_431),
.C(n_427),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_619),
.A2(n_620),
.B(n_600),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_589),
.A2(n_431),
.B(n_427),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_621),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_611),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_583),
.B(n_427),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_611),
.Y(n_677)
);

AOI221x1_ASAP7_75t_L g678 ( 
.A1(n_622),
.A2(n_439),
.B1(n_427),
.B2(n_14),
.C(n_15),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_594),
.A2(n_579),
.B(n_627),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_622),
.A2(n_583),
.B(n_602),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_586),
.Y(n_681)
);

AOI211x1_ASAP7_75t_L g682 ( 
.A1(n_581),
.A2(n_10),
.B(n_13),
.C(n_14),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_564),
.A2(n_565),
.B(n_586),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_587),
.Y(n_684)
);

NAND2x1_ASAP7_75t_L g685 ( 
.A(n_590),
.B(n_418),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_626),
.B(n_418),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_566),
.B(n_52),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_665),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_650),
.A2(n_629),
.B1(n_588),
.B2(n_582),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_634),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_673),
.A2(n_564),
.B(n_565),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_645),
.B(n_614),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_637),
.A2(n_585),
.B1(n_650),
.B2(n_636),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_642),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_658),
.A2(n_564),
.B(n_565),
.Y(n_696)
);

BUFx12f_ASAP7_75t_L g697 ( 
.A(n_660),
.Y(n_697)
);

NOR2x1_ASAP7_75t_SL g698 ( 
.A(n_647),
.B(n_564),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_643),
.A2(n_590),
.B(n_614),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_647),
.Y(n_700)
);

A2O1A1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_630),
.A2(n_582),
.B(n_580),
.C(n_617),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_637),
.A2(n_591),
.B1(n_587),
.B2(n_617),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_653),
.Y(n_703)
);

BUFx4f_ASAP7_75t_L g704 ( 
.A(n_656),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_648),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_632),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_632),
.B(n_611),
.Y(n_707)
);

BUFx12f_ASAP7_75t_L g708 ( 
.A(n_656),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_655),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_645),
.B(n_591),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_648),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_656),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_631),
.A2(n_602),
.B(n_580),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_672),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_663),
.A2(n_668),
.B(n_641),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_635),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_644),
.A2(n_591),
.B1(n_610),
.B2(n_567),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_664),
.A2(n_640),
.B(n_659),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_644),
.A2(n_567),
.B(n_603),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_683),
.B(n_572),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_SL g721 ( 
.A1(n_682),
.A2(n_595),
.B1(n_574),
.B2(n_576),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_649),
.A2(n_54),
.B(n_53),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_SL g723 ( 
.A1(n_669),
.A2(n_603),
.B(n_609),
.C(n_108),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_675),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_670),
.A2(n_609),
.B1(n_17),
.B2(n_18),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_684),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_680),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_654),
.B(n_19),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

BUFx12f_ASAP7_75t_L g731 ( 
.A(n_633),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_649),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_679),
.A2(n_111),
.B(n_199),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_677),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_657),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_664),
.A2(n_106),
.B(n_195),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_688),
.B(n_55),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_676),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_688),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_657),
.B(n_20),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_681),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_738),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_693),
.B(n_676),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_719),
.A2(n_646),
.B1(n_652),
.B2(n_638),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_717),
.A2(n_662),
.B1(n_651),
.B2(n_686),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_694),
.A2(n_686),
.B1(n_687),
.B2(n_651),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_706),
.B(n_633),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_704),
.B(n_681),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_690),
.A2(n_721),
.B1(n_728),
.B2(n_739),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_708),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_727),
.A2(n_666),
.B1(n_678),
.B2(n_667),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_730),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_689),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_SL g754 ( 
.A1(n_701),
.A2(n_671),
.B(n_733),
.C(n_732),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_715),
.A2(n_687),
.B(n_666),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_689),
.Y(n_756)
);

CKINVDCx16_ASAP7_75t_R g757 ( 
.A(n_697),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_740),
.B(n_674),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_699),
.B(n_661),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_691),
.B(n_639),
.Y(n_760)
);

AO21x2_ASAP7_75t_L g761 ( 
.A1(n_718),
.A2(n_639),
.B(n_674),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_697),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_708),
.Y(n_763)
);

AOI221xp5_ASAP7_75t_L g764 ( 
.A1(n_725),
.A2(n_674),
.B1(n_639),
.B2(n_685),
.C(n_25),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_737),
.A2(n_639),
.B1(n_674),
.B2(n_24),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_734),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_704),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_732),
.B(n_21),
.Y(n_768)
);

NAND2x1_ASAP7_75t_L g769 ( 
.A(n_741),
.B(n_57),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_737),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_734),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_703),
.B(n_64),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_731),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_710),
.A2(n_26),
.B(n_27),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_738),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_703),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_741),
.B(n_65),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_702),
.B(n_27),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_731),
.Y(n_779)
);

CKINVDCx6p67_ASAP7_75t_R g780 ( 
.A(n_712),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_705),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_707),
.A2(n_118),
.B(n_192),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_724),
.B(n_28),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_714),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_700),
.B(n_705),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_711),
.A2(n_700),
.B1(n_720),
.B2(n_704),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_720),
.Y(n_787)
);

CKINVDCx6p67_ASAP7_75t_R g788 ( 
.A(n_712),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_711),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_720),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_735),
.B(n_31),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_729),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_729),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_714),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_707),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_737),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_713),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_718),
.A2(n_121),
.B(n_191),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_696),
.A2(n_120),
.B(n_189),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_726),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_713),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_695),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_776),
.B(n_742),
.Y(n_803)
);

AOI221xp5_ASAP7_75t_L g804 ( 
.A1(n_796),
.A2(n_723),
.B1(n_722),
.B2(n_709),
.C(n_716),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_776),
.B(n_696),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_789),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_774),
.A2(n_737),
.B1(n_736),
.B2(n_709),
.Y(n_807)
);

AOI33xp33_ASAP7_75t_L g808 ( 
.A1(n_770),
.A2(n_32),
.A3(n_33),
.B1(n_35),
.B2(n_36),
.B3(n_37),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_778),
.A2(n_698),
.B1(n_736),
.B2(n_699),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_758),
.B(n_716),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_785),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_SL g812 ( 
.A1(n_749),
.A2(n_695),
.B(n_37),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_744),
.A2(n_692),
.B(n_698),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_766),
.A2(n_692),
.B1(n_38),
.B2(n_39),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_743),
.B(n_35),
.Y(n_815)
);

AOI221xp5_ASAP7_75t_L g816 ( 
.A1(n_764),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.C(n_44),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_743),
.B(n_40),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_745),
.A2(n_42),
.B(n_45),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_L g819 ( 
.A1(n_790),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_778),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_780),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_787),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_742),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_791),
.A2(n_49),
.B1(n_50),
.B2(n_66),
.Y(n_824)
);

OAI221xp5_ASAP7_75t_L g825 ( 
.A1(n_751),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.C(n_70),
.Y(n_825)
);

AND2x2_ASAP7_75t_SL g826 ( 
.A(n_765),
.B(n_71),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_772),
.A2(n_72),
.B1(n_74),
.B2(n_78),
.Y(n_827)
);

OAI211xp5_ASAP7_75t_L g828 ( 
.A1(n_781),
.A2(n_80),
.B(n_81),
.C(n_84),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_802),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_772),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_756),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_831)
);

AO221x2_ASAP7_75t_L g832 ( 
.A1(n_786),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_787),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_760),
.B(n_98),
.Y(n_834)
);

OAI211xp5_ASAP7_75t_L g835 ( 
.A1(n_768),
.A2(n_99),
.B(n_100),
.C(n_102),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_785),
.B(n_105),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_772),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_777),
.A2(n_753),
.B1(n_795),
.B2(n_747),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_775),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_784),
.Y(n_840)
);

OAI221xp5_ASAP7_75t_L g841 ( 
.A1(n_746),
.A2(n_115),
.B1(n_117),
.B2(n_122),
.C(n_124),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_777),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_756),
.B(n_141),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_759),
.B(n_143),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_775),
.B(n_200),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_757),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_761),
.B(n_188),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_777),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_848)
);

AOI221xp5_ASAP7_75t_L g849 ( 
.A1(n_754),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.C(n_154),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_799),
.A2(n_155),
.B(n_157),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_747),
.B(n_159),
.Y(n_851)
);

OAI211xp5_ASAP7_75t_L g852 ( 
.A1(n_783),
.A2(n_160),
.B(n_163),
.C(n_166),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_810),
.B(n_761),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_810),
.B(n_811),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_805),
.B(n_797),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_829),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_805),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_805),
.B(n_801),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_829),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_806),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_840),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_840),
.Y(n_862)
);

INVx8_ASAP7_75t_L g863 ( 
.A(n_844),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_803),
.B(n_794),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_826),
.A2(n_771),
.B1(n_755),
.B2(n_762),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_803),
.B(n_794),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_784),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_839),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_844),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_839),
.B(n_759),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_822),
.Y(n_871)
);

AOI221xp5_ASAP7_75t_L g872 ( 
.A1(n_816),
.A2(n_754),
.B1(n_782),
.B2(n_752),
.C(n_800),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_823),
.B(n_759),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_847),
.Y(n_874)
);

AO221x2_ASAP7_75t_L g875 ( 
.A1(n_812),
.A2(n_818),
.B1(n_814),
.B2(n_832),
.C(n_817),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_847),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_813),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_844),
.Y(n_878)
);

NOR2x1_ASAP7_75t_SL g879 ( 
.A(n_844),
.B(n_798),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_822),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_822),
.B(n_759),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_833),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_850),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_833),
.B(n_798),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_850),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_834),
.B(n_799),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_845),
.Y(n_887)
);

NOR2x1_ASAP7_75t_L g888 ( 
.A(n_871),
.B(n_821),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_857),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_854),
.B(n_853),
.Y(n_890)
);

AOI221xp5_ASAP7_75t_L g891 ( 
.A1(n_865),
.A2(n_820),
.B1(n_815),
.B2(n_819),
.C(n_824),
.Y(n_891)
);

AOI221xp5_ASAP7_75t_L g892 ( 
.A1(n_865),
.A2(n_825),
.B1(n_849),
.B2(n_841),
.C(n_852),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_856),
.Y(n_893)
);

OR2x6_ASAP7_75t_L g894 ( 
.A(n_863),
.B(n_833),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_860),
.Y(n_895)
);

OAI31xp33_ASAP7_75t_L g896 ( 
.A1(n_877),
.A2(n_835),
.A3(n_828),
.B(n_843),
.Y(n_896)
);

OAI33xp33_ASAP7_75t_L g897 ( 
.A1(n_860),
.A2(n_793),
.A3(n_808),
.B1(n_762),
.B2(n_773),
.B3(n_832),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_866),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_875),
.A2(n_826),
.B1(n_832),
.B2(n_807),
.Y(n_899)
);

BUFx8_ASAP7_75t_L g900 ( 
.A(n_871),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_868),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_856),
.Y(n_902)
);

NAND4xp25_ASAP7_75t_SL g903 ( 
.A(n_872),
.B(n_808),
.C(n_831),
.D(n_846),
.Y(n_903)
);

AOI221xp5_ASAP7_75t_L g904 ( 
.A1(n_877),
.A2(n_834),
.B1(n_836),
.B2(n_804),
.C(n_838),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_859),
.Y(n_905)
);

OAI321xp33_ASAP7_75t_L g906 ( 
.A1(n_872),
.A2(n_848),
.A3(n_842),
.B1(n_827),
.B2(n_837),
.C(n_830),
.Y(n_906)
);

AOI211xp5_ASAP7_75t_L g907 ( 
.A1(n_878),
.A2(n_851),
.B(n_836),
.C(n_821),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_868),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_SL g909 ( 
.A1(n_869),
.A2(n_845),
.B(n_767),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_875),
.A2(n_851),
.B1(n_771),
.B2(n_809),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_854),
.B(n_874),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_911),
.B(n_857),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_890),
.B(n_874),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_898),
.B(n_876),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_894),
.B(n_876),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_901),
.B(n_853),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_901),
.B(n_853),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_893),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_903),
.A2(n_875),
.B1(n_869),
.B2(n_863),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_893),
.B(n_859),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_895),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_908),
.B(n_857),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_908),
.B(n_857),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_889),
.B(n_855),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_888),
.B(n_869),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_SL g926 ( 
.A(n_899),
.B(n_869),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_921),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_914),
.B(n_902),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_920),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_924),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_918),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_916),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_913),
.B(n_905),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_920),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_915),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_918),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_912),
.B(n_889),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_932),
.B(n_912),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_931),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_SL g940 ( 
.A(n_928),
.B(n_899),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_927),
.Y(n_941)
);

NOR2x1_ASAP7_75t_L g942 ( 
.A(n_936),
.B(n_925),
.Y(n_942)
);

NAND4xp75_ASAP7_75t_L g943 ( 
.A(n_929),
.B(n_919),
.C(n_892),
.D(n_896),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_933),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_930),
.B(n_917),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_936),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_935),
.B(n_925),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_929),
.Y(n_948)
);

AOI222xp33_ASAP7_75t_L g949 ( 
.A1(n_940),
.A2(n_926),
.B1(n_891),
.B2(n_897),
.C1(n_904),
.C2(n_906),
.Y(n_949)
);

OAI222xp33_ASAP7_75t_L g950 ( 
.A1(n_947),
.A2(n_910),
.B1(n_925),
.B2(n_894),
.C1(n_878),
.C2(n_926),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_941),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_943),
.A2(n_907),
.B1(n_894),
.B2(n_863),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_946),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_951),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_951),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_952),
.Y(n_956)
);

NOR4xp25_ASAP7_75t_SL g957 ( 
.A(n_955),
.B(n_940),
.C(n_953),
.D(n_950),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_949),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_954),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_955),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_944),
.Y(n_961)
);

NOR2xp67_ASAP7_75t_L g962 ( 
.A(n_959),
.B(n_939),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_957),
.A2(n_942),
.B(n_939),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_958),
.B(n_938),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_SL g965 ( 
.A(n_959),
.B(n_773),
.C(n_945),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_959),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_SL g967 ( 
.A(n_957),
.B(n_948),
.C(n_938),
.Y(n_967)
);

NAND4xp25_ASAP7_75t_L g968 ( 
.A(n_958),
.B(n_750),
.C(n_763),
.D(n_851),
.Y(n_968)
);

AOI222xp33_ASAP7_75t_L g969 ( 
.A1(n_967),
.A2(n_965),
.B1(n_964),
.B2(n_962),
.C1(n_966),
.C2(n_961),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_863),
.B(n_934),
.C(n_763),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_968),
.A2(n_875),
.B(n_934),
.Y(n_971)
);

NOR4xp25_ASAP7_75t_SL g972 ( 
.A(n_966),
.B(n_779),
.C(n_875),
.D(n_750),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_966),
.B(n_937),
.Y(n_973)
);

NAND4xp25_ASAP7_75t_L g974 ( 
.A(n_967),
.B(n_871),
.C(n_886),
.D(n_937),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_963),
.A2(n_931),
.B1(n_923),
.B2(n_922),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_973),
.B(n_779),
.Y(n_976)
);

AOI322xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_863),
.A3(n_909),
.B1(n_886),
.B2(n_880),
.C1(n_882),
.C2(n_883),
.Y(n_977)
);

NOR4xp25_ASAP7_75t_L g978 ( 
.A(n_974),
.B(n_767),
.C(n_883),
.D(n_885),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_969),
.A2(n_900),
.B1(n_863),
.B2(n_881),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_972),
.B(n_780),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_975),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_971),
.A2(n_900),
.B1(n_881),
.B2(n_884),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_973),
.B(n_889),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_981),
.B(n_167),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_979),
.Y(n_985)
);

NAND5xp2_ASAP7_75t_L g986 ( 
.A(n_982),
.B(n_748),
.C(n_886),
.D(n_885),
.E(n_887),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_976),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_983),
.B(n_880),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_978),
.A2(n_882),
.B1(n_792),
.B2(n_884),
.C(n_747),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_977),
.B(n_788),
.Y(n_991)
);

XNOR2xp5_ASAP7_75t_L g992 ( 
.A(n_979),
.B(n_748),
.Y(n_992)
);

NOR2x1_ASAP7_75t_L g993 ( 
.A(n_983),
.B(n_769),
.Y(n_993)
);

OAI221xp5_ASAP7_75t_R g994 ( 
.A1(n_979),
.A2(n_900),
.B1(n_879),
.B2(n_788),
.C(n_884),
.Y(n_994)
);

AOI222xp33_ASAP7_75t_L g995 ( 
.A1(n_989),
.A2(n_879),
.B1(n_884),
.B2(n_887),
.C1(n_881),
.C2(n_873),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_SL g996 ( 
.A(n_987),
.B(n_873),
.C(n_862),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_984),
.Y(n_997)
);

AOI211x1_ASAP7_75t_L g998 ( 
.A1(n_985),
.A2(n_862),
.B(n_873),
.C(n_870),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_988),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_991),
.B(n_992),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_986),
.C(n_990),
.Y(n_1001)
);

AOI211x1_ASAP7_75t_SL g1002 ( 
.A1(n_994),
.A2(n_861),
.B(n_170),
.C(n_171),
.Y(n_1002)
);

NAND5xp2_ASAP7_75t_L g1003 ( 
.A(n_989),
.B(n_870),
.C(n_858),
.D(n_855),
.E(n_867),
.Y(n_1003)
);

NOR2x1p5_ASAP7_75t_L g1004 ( 
.A(n_989),
.B(n_881),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_1004),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_997),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_1000),
.Y(n_1007)
);

OAI21xp33_ASAP7_75t_SL g1008 ( 
.A1(n_995),
.A2(n_858),
.B(n_855),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_999),
.B(n_858),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_L g1010 ( 
.A(n_996),
.B(n_168),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1005),
.B(n_1001),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_1010),
.Y(n_1012)
);

XOR2xp5_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_1002),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_1012),
.A2(n_1006),
.B(n_1009),
.C(n_1008),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_1013),
.A2(n_998),
.B1(n_1003),
.B2(n_866),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1015),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1014),
.Y(n_1017)
);

AO221x1_ASAP7_75t_L g1018 ( 
.A1(n_1017),
.A2(n_1016),
.B1(n_1011),
.B2(n_868),
.C(n_177),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1017),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1018),
.A2(n_868),
.B1(n_861),
.B2(n_864),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1020),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_1021),
.A2(n_1019),
.B1(n_173),
.B2(n_175),
.C(n_178),
.Y(n_1022)
);

AOI211xp5_ASAP7_75t_L g1023 ( 
.A1(n_1022),
.A2(n_172),
.B(n_179),
.C(n_184),
.Y(n_1023)
);


endmodule