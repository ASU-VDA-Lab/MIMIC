module fake_jpeg_22522_n_305 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_25),
.B1(n_27),
.B2(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_25),
.B2(n_29),
.Y(n_44)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_47),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_50),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_30),
.C(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_29),
.B1(n_21),
.B2(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_29),
.B1(n_18),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_29),
.B1(n_21),
.B2(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_82),
.B1(n_85),
.B2(n_17),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_40),
.B1(n_43),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_64),
.B1(n_65),
.B2(n_63),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_40),
.C(n_18),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_0),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_78),
.B1(n_84),
.B2(n_50),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_40),
.B1(n_31),
.B2(n_23),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_32),
.B1(n_22),
.B2(n_19),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_17),
.B1(n_46),
.B2(n_9),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_22),
.B1(n_19),
.B2(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_31),
.B1(n_26),
.B2(n_20),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_92),
.Y(n_116)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_78),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_96),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_58),
.B(n_45),
.C(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_110),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_60),
.B1(n_55),
.B2(n_62),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_114),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_62),
.B1(n_26),
.B2(n_20),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_46),
.B1(n_61),
.B2(n_26),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_92),
.B1(n_77),
.B2(n_103),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_120),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_20),
.B(n_17),
.C(n_46),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_113),
.B(n_71),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_109),
.B1(n_70),
.B2(n_113),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_93),
.Y(n_118)
);

NAND2x1_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_67),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_122),
.A2(n_129),
.B(n_132),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_138),
.B1(n_100),
.B2(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_145),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_75),
.B(n_73),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_121),
.C(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_74),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_86),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_86),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_79),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_67),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_150),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_109),
.B(n_69),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_151),
.B(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_123),
.B1(n_149),
.B2(n_124),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_118),
.B(n_119),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_165),
.B(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_162),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_109),
.B1(n_108),
.B2(n_95),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_177),
.B1(n_123),
.B2(n_127),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_95),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_171),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_130),
.C(n_147),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_97),
.A3(n_88),
.B1(n_105),
.B2(n_10),
.C1(n_12),
.C2(n_16),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_1),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_88),
.B1(n_105),
.B2(n_3),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_175),
.B1(n_143),
.B2(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_179),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_126),
.B1(n_145),
.B2(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_1),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_128),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_2),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_130),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_157),
.Y(n_210)
);

OA21x2_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_129),
.B(n_132),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_197),
.B(n_153),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_200),
.B1(n_166),
.B2(n_177),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_205),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_131),
.B(n_125),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_205),
.B(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_172),
.B1(n_165),
.B2(n_158),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_198),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_199),
.C(n_201),
.Y(n_208)
);

OA21x2_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_149),
.B(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_136),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_134),
.C(n_135),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_2),
.C(n_4),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_204),
.C(n_176),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_4),
.C(n_5),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_5),
.C(n_6),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_171),
.C(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_197),
.B(n_183),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_224),
.Y(n_232)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_192),
.B(n_169),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_178),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_217),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_155),
.B(n_173),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_228),
.B(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_186),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_160),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_229),
.B(n_10),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_187),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_158),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_227),
.B1(n_192),
.B2(n_195),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_170),
.C(n_163),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_199),
.C(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_159),
.B(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_231),
.A2(n_235),
.B(n_216),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_189),
.B(n_184),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_185),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_191),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_214),
.B1(n_223),
.B2(n_222),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_184),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_181),
.C(n_163),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_181),
.C(n_203),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_204),
.C(n_206),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_174),
.C(n_154),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_246),
.B1(n_212),
.B2(n_211),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_215),
.B1(n_229),
.B2(n_217),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_213),
.B(n_218),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_260),
.B(n_235),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_237),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_238),
.C(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_254),
.B(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_11),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_210),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_7),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_266),
.C(n_255),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_243),
.C(n_218),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_268),
.B(n_15),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_230),
.B(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_221),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_5),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_263),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_9),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_258),
.B(n_250),
.C(n_249),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_284),
.B(n_286),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_271),
.C(n_273),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_250),
.B(n_253),
.C(n_249),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_275),
.B(n_6),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_283),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_11),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_282),
.Y(n_296)
);

NAND4xp25_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_266),
.C(n_265),
.D(n_269),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_290),
.B(n_292),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_16),
.B1(n_15),
.B2(n_6),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_281),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_291),
.C(n_300),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_6),
.B(n_280),
.C(n_292),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_299),
.B(n_297),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_303),
.Y(n_305)
);


endmodule