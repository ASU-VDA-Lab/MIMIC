module fake_jpeg_4608_n_197 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_197);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_36),
.A2(n_44),
.B(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_37),
.B(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_21),
.B(n_2),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_27),
.B1(n_15),
.B2(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_26),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_35),
.B1(n_26),
.B2(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_52),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_6),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_8),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_35),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_61),
.Y(n_102)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_68),
.B(n_79),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_34),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_23),
.B1(n_18),
.B2(n_15),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_22),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_88),
.Y(n_104)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_78),
.B1(n_84),
.B2(n_8),
.Y(n_99)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_36),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_8),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_56),
.C(n_77),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_110),
.C(n_101),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_29),
.B1(n_32),
.B2(n_12),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_108),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_9),
.B(n_67),
.C(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_60),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_66),
.B1(n_76),
.B2(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_76),
.B1(n_61),
.B2(n_58),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_58),
.A3(n_65),
.B1(n_82),
.B2(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_65),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_118),
.B(n_125),
.Y(n_156)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_124),
.Y(n_149)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_137),
.Y(n_143)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_98),
.B(n_114),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_97),
.C(n_101),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_139),
.C(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_91),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_110),
.C(n_105),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_92),
.B1(n_95),
.B2(n_116),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_142),
.B(n_156),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_147),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_117),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_105),
.C(n_104),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_104),
.C(n_114),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_155),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_153),
.B(n_154),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_95),
.B(n_114),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_107),
.B(n_112),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_121),
.B1(n_135),
.B2(n_119),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_127),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_120),
.B1(n_130),
.B2(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_164),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_119),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_168),
.B(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_153),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_140),
.B(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_158),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_144),
.A3(n_152),
.B1(n_165),
.B2(n_166),
.C1(n_170),
.C2(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_148),
.C(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_163),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_185),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_188),
.B1(n_181),
.B2(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_173),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_162),
.B1(n_172),
.B2(n_175),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.C(n_176),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_175),
.B1(n_181),
.B2(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_191),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_174),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_192),
.Y(n_197)
);


endmodule