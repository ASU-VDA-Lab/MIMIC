module real_jpeg_30016_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_327, n_326, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_327;
input n_326;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_1),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_33),
.B1(n_35),
.B2(n_134),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_1),
.A2(n_99),
.B1(n_100),
.B2(n_134),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_1),
.A2(n_134),
.B1(n_155),
.B2(n_161),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_34),
.B(n_35),
.C(n_39),
.D(n_42),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_2),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_61),
.B(n_65),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_99),
.B(n_101),
.C(n_102),
.D(n_104),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_2),
.B(n_99),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_2),
.A2(n_100),
.B(n_131),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_2),
.A2(n_83),
.B1(n_155),
.B2(n_161),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_57),
.B1(n_99),
.B2(n_100),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_57),
.B1(n_155),
.B2(n_161),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_5),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_5),
.A2(n_33),
.B1(n_35),
.B2(n_151),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_5),
.A2(n_99),
.B1(n_100),
.B2(n_151),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_5),
.A2(n_151),
.B1(n_155),
.B2(n_161),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_7),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_114),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_7),
.A2(n_99),
.B1(n_100),
.B2(n_114),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_7),
.A2(n_114),
.B1(n_155),
.B2(n_161),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_8),
.A2(n_44),
.B1(n_99),
.B2(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_44),
.B1(n_155),
.B2(n_161),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_10),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_214),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_10),
.A2(n_99),
.B1(n_100),
.B2(n_214),
.Y(n_301)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_11),
.A2(n_35),
.B(n_40),
.C(n_41),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_195),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_12),
.A2(n_99),
.B1(n_100),
.B2(n_195),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_12),
.A2(n_155),
.B1(n_161),
.B2(n_195),
.Y(n_319)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_15),
.A2(n_33),
.B1(n_35),
.B2(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_15),
.A2(n_64),
.B1(n_99),
.B2(n_100),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_15),
.A2(n_64),
.B1(n_155),
.B2(n_161),
.Y(n_206)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_310),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_274),
.A3(n_303),
.B1(n_308),
.B2(n_309),
.C(n_326),
.Y(n_18)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_224),
.A3(n_263),
.B1(n_268),
.B2(n_273),
.C(n_327),
.Y(n_19)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_175),
.C(n_220),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_142),
.B(n_174),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_119),
.B(n_141),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_94),
.B(n_118),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_70),
.B(n_93),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_26),
.B(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_38),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.A3(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_28),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_37),
.Y(n_36)
);

NAND2x1_ASAP7_75t_SL g61 ( 
.A(n_29),
.B(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_33),
.B(n_52),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_35),
.A2(n_100),
.A3(n_101),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_39),
.A2(n_41),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_39),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_39),
.A2(n_41),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_39),
.A2(n_41),
.B1(n_240),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_42),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_56),
.B(n_58),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_45),
.A2(n_58),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_45),
.A2(n_138),
.B1(n_173),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_45),
.A2(n_138),
.B1(n_197),
.B2(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_45),
.A2(n_138),
.B(n_249),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_60),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_55),
.C(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_50),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_50),
.A2(n_102),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_50),
.A2(n_102),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_50),
.A2(n_102),
.B1(n_252),
.B2(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_50),
.A2(n_102),
.B(n_316),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_53),
.B1(n_99),
.B2(n_100),
.Y(n_103)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_56),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_61),
.A2(n_78),
.B1(n_113),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_61),
.A2(n_69),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_61),
.A2(n_194),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_61),
.A2(n_78),
.B(n_213),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_86),
.B(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_SL g212 ( 
.A(n_68),
.Y(n_212)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_83),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_80),
.B(n_92),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_79),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_78),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_75),
.A2(n_77),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_91),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_83),
.B(n_128),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_83),
.A2(n_130),
.B(n_154),
.C(n_155),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_96),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_97),
.B(n_120),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_107),
.CI(n_110),
.CON(n_97),
.SN(n_97)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_100),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_124),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_106),
.A2(n_183),
.B1(n_209),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_106),
.A2(n_183),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_135),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_136),
.C(n_137),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_127),
.C(n_132),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_187),
.B(n_189),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_128),
.A2(n_189),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_128),
.A2(n_231),
.B1(n_259),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_128),
.A2(n_231),
.B1(n_286),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_159),
.B1(n_188),
.B2(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_129),
.A2(n_159),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_131),
.B1(n_155),
.B2(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_144),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_157),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_146),
.B(n_147),
.C(n_157),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_156),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_168),
.C(n_171),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B(n_163),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_164),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_176),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_199),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_177),
.B(n_199),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_191),
.C(n_198),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_181),
.C(n_190),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_186),
.B2(n_190),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B(n_185),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_198),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_196),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_210),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_201),
.B(n_210),
.C(n_219),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_215),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_221),
.B(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_244),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.C(n_243),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_236),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_235),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_233),
.C(n_235),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_242),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_242),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_242),
.A2(n_257),
.B(n_260),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_262),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_254),
.B1(n_255),
.B2(n_261),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_250),
.B(n_253),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_250),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_253),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_253),
.A2(n_276),
.B1(n_277),
.B2(n_288),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_261),
.C(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_269),
.B(n_272),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_291),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_291),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_288),
.C(n_289),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_285),
.B2(n_287),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_280),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_284),
.C(n_285),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_281),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_282),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_284),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_295),
.C(n_299),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_287),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_294),
.C(n_302),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_290),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_302),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_296),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_324),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_323),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_323),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_322),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_315),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_317),
.Y(n_320)
);


endmodule