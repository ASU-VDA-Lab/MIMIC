module fake_jpeg_16632_n_386 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_7),
.B1(n_12),
.B2(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_17),
.B1(n_36),
.B2(n_32),
.Y(n_72)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_21),
.A2(n_13),
.B(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_6),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_8),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_16),
.B1(n_15),
.B2(n_25),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_35),
.Y(n_75)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_8),
.C(n_12),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_29),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_73),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_72),
.A2(n_93),
.B1(n_4),
.B2(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_29),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_75),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_77),
.B(n_82),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g157 ( 
.A(n_81),
.B(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_42),
.B(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_110),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_26),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_87),
.A2(n_104),
.B(n_106),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_38),
.A2(n_18),
.B1(n_31),
.B2(n_28),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_117),
.B1(n_9),
.B2(n_11),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_103),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_19),
.B1(n_18),
.B2(n_32),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_39),
.A2(n_19),
.B1(n_36),
.B2(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_102),
.B1(n_116),
.B2(n_5),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_18),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_111),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_16),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_43),
.B(n_15),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_26),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_44),
.A2(n_37),
.B1(n_32),
.B2(n_17),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_86),
.B1(n_92),
.B2(n_114),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_40),
.B(n_17),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_58),
.B(n_16),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_45),
.A2(n_25),
.B1(n_35),
.B2(n_2),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_63),
.A2(n_25),
.B1(n_8),
.B2(n_3),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_127),
.Y(n_175)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_120),
.Y(n_179)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_122),
.A2(n_140),
.B1(n_144),
.B2(n_146),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_123),
.A2(n_152),
.B1(n_118),
.B2(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_5),
.B1(n_11),
.B2(n_3),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_128),
.A2(n_134),
.B1(n_160),
.B2(n_113),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_135),
.Y(n_176)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_131),
.B(n_139),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_150),
.B1(n_130),
.B2(n_142),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_86),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_4),
.B1(n_10),
.B2(n_13),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_153),
.Y(n_181)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_13),
.B1(n_0),
.B2(n_1),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_68),
.B(n_0),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_145),
.B(n_148),
.Y(n_209)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_13),
.C(n_1),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_73),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_162),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_106),
.B1(n_100),
.B2(n_116),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_99),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_88),
.A2(n_106),
.B1(n_111),
.B2(n_84),
.Y(n_154)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_79),
.A2(n_114),
.B1(n_112),
.B2(n_107),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_163),
.B1(n_122),
.B2(n_119),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_69),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_161),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_79),
.A2(n_109),
.B1(n_112),
.B2(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_74),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_84),
.B(n_71),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_109),
.A2(n_107),
.B1(n_76),
.B2(n_74),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_129),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_67),
.A2(n_81),
.B1(n_97),
.B2(n_76),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_120),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_211),
.B1(n_161),
.B2(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_129),
.B(n_95),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_191),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_95),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_207),
.B(n_181),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_189),
.B(n_188),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_195),
.B1(n_196),
.B2(n_178),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_124),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_194),
.B1(n_213),
.B2(n_178),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_124),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_204),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_137),
.B1(n_123),
.B2(n_138),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_128),
.A2(n_156),
.B1(n_154),
.B2(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

AOI22x1_ASAP7_75t_R g198 ( 
.A1(n_156),
.A2(n_124),
.B1(n_145),
.B2(n_157),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_157),
.B(n_125),
.C(n_127),
.D(n_131),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_133),
.B(n_125),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_199),
.B(n_203),
.Y(n_233)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_141),
.B(n_121),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_159),
.B1(n_164),
.B2(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_215),
.B(n_239),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_217),
.B(n_223),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_218),
.A2(n_228),
.B1(n_229),
.B2(n_240),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_250),
.B(n_243),
.Y(n_257)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_221),
.A2(n_227),
.B1(n_236),
.B2(n_238),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_186),
.B(n_193),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_224),
.A2(n_239),
.B(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_174),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_231),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_206),
.B1(n_210),
.B2(n_212),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_173),
.A2(n_194),
.B1(n_192),
.B2(n_183),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_189),
.B1(n_169),
.B2(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_177),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_191),
.C(n_185),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_222),
.C(n_230),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_176),
.B(n_208),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_175),
.B1(n_182),
.B2(n_188),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_253),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_176),
.B(n_181),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_244),
.B(n_219),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_175),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_180),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_187),
.A2(n_213),
.B(n_172),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_174),
.B(n_197),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_246),
.B(n_233),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_207),
.B1(n_199),
.B2(n_202),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_277),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_205),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_255),
.B(n_256),
.C(n_265),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_244),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_257),
.A2(n_258),
.B(n_259),
.Y(n_309)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_275),
.B1(n_261),
.B2(n_263),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_222),
.A2(n_230),
.B(n_241),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_267),
.A2(n_279),
.B(n_283),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_275),
.B(n_280),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_228),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_276),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_237),
.B(n_225),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_273),
.B(n_281),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_241),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_223),
.B(n_225),
.C(n_221),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_234),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_236),
.A2(n_238),
.B(n_250),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_232),
.Y(n_284)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_216),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_262),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_250),
.B1(n_229),
.B2(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_250),
.B1(n_232),
.B2(n_247),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_294),
.B1(n_295),
.B2(n_306),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_287),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_296),
.B(n_302),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_249),
.B1(n_231),
.B2(n_215),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_220),
.B1(n_272),
.B2(n_274),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_260),
.A2(n_267),
.B1(n_270),
.B2(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_260),
.A2(n_258),
.B1(n_280),
.B2(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_301),
.B(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_268),
.A2(n_256),
.B(n_269),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_277),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_286),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_265),
.A2(n_283),
.B1(n_279),
.B2(n_259),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_307),
.B(n_315),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_268),
.A3(n_266),
.B1(n_278),
.B2(n_255),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_308),
.B(n_310),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_271),
.A2(n_286),
.B(n_285),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_312),
.A2(n_307),
.B1(n_292),
.B2(n_305),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_313),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_271),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_302),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_306),
.C(n_288),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_308),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_324),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_326),
.A2(n_335),
.B1(n_300),
.B2(n_297),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_296),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_327),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_304),
.B(n_294),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_328),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_305),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_329),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_303),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_291),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_303),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_300),
.B(n_288),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_351),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_298),
.C(n_310),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_343),
.C(n_349),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_290),
.C(n_309),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_293),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_348),
.B(n_329),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_299),
.C(n_297),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_320),
.A2(n_293),
.B1(n_313),
.B2(n_289),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_351),
.A2(n_353),
.B1(n_317),
.B2(n_332),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_332),
.A2(n_320),
.B1(n_323),
.B2(n_326),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_354),
.A2(n_365),
.B1(n_340),
.B2(n_328),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_355),
.A2(n_344),
.B(n_346),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_333),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_356),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_325),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_358),
.C(n_362),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_325),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_363),
.C(n_364),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_336),
.C(n_330),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_334),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_336),
.C(n_335),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_324),
.Y(n_365)
);

XOR2x1_ASAP7_75t_SL g366 ( 
.A(n_361),
.B(n_348),
.Y(n_366)
);

AO21x1_ASAP7_75t_L g375 ( 
.A1(n_366),
.A2(n_372),
.B(n_352),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_371),
.Y(n_376)
);

AO221x1_ASAP7_75t_L g372 ( 
.A1(n_362),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.C(n_318),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_373),
.B(n_374),
.Y(n_377)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_369),
.Y(n_374)
);

AOI322xp5_ASAP7_75t_L g379 ( 
.A1(n_375),
.A2(n_366),
.A3(n_360),
.B1(n_370),
.B2(n_323),
.C1(n_346),
.C2(n_350),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_359),
.C(n_363),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_359),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_345),
.Y(n_380)
);

AOI21x1_ASAP7_75t_L g382 ( 
.A1(n_380),
.A2(n_381),
.B(n_370),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_382),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_380),
.B(n_377),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_353),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_338),
.Y(n_386)
);


endmodule