module fake_aes_10113_n_665 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_665);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_665;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_50), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_88), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_8), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_45), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_23), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_86), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_9), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_38), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_81), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_68), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_5), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_20), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_27), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_3), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_31), .Y(n_108) );
BUFx2_ASAP7_75t_SL g109 ( .A(n_32), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_47), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_5), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_28), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_48), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_63), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_43), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_0), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_12), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_52), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_46), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_35), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_25), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_17), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_4), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_51), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_103), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_127), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_105), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_99), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_99), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_92), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_90), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_101), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_127), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
NOR2xp67_ASAP7_75t_L g146 ( .A(n_98), .B(n_3), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_100), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_97), .B(n_4), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_97), .B(n_6), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_101), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_126), .B(n_7), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_100), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_126), .B(n_8), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_104), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_104), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_132), .A2(n_120), .B1(n_102), .B2(n_110), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_141), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_132), .B(n_102), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_131), .B(n_120), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_149), .B(n_93), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_149), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_133), .B(n_94), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_131), .B(n_95), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_149), .B(n_128), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_147), .B(n_106), .Y(n_172) );
AOI22x1_ASAP7_75t_L g173 ( .A1(n_156), .A2(n_109), .B1(n_108), .B2(n_124), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_136), .B(n_90), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_157), .B(n_128), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_157), .B(n_119), .Y(n_178) );
CKINVDCx8_ASAP7_75t_R g179 ( .A(n_130), .Y(n_179) );
BUFx10_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_134), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_139), .B(n_114), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_139), .B(n_111), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_145), .B(n_115), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_178), .A2(n_153), .B1(n_151), .B2(n_146), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_174), .B(n_145), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_167), .B(n_146), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_180), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_166), .A2(n_155), .B1(n_154), .B2(n_138), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_180), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_166), .A2(n_140), .B1(n_155), .B2(n_154), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_178), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_180), .B(n_152), .Y(n_200) );
NOR2x2_ASAP7_75t_L g201 ( .A(n_169), .B(n_140), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_187), .B(n_151), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_175), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_162), .B(n_153), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_159), .B(n_152), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_175), .B(n_111), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_165), .B(n_135), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_181), .B(n_116), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_171), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_171), .B(n_112), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_181), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_176), .B(n_116), .Y(n_214) );
BUFx6f_ASAP7_75t_SL g215 ( .A(n_166), .Y(n_215) );
BUFx8_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_159), .B(n_176), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_158), .B(n_135), .Y(n_219) );
INVxp67_ASAP7_75t_SL g220 ( .A(n_161), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_159), .B(n_152), .Y(n_221) );
AND2x6_ASAP7_75t_L g222 ( .A(n_163), .B(n_118), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_166), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_164), .A2(n_107), .B1(n_113), .B2(n_117), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_166), .B(n_135), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_177), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_168), .B(n_135), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_188), .B(n_123), .Y(n_230) );
INVx5_ASAP7_75t_L g231 ( .A(n_191), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_160), .A2(n_137), .B1(n_143), .B2(n_138), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_179), .B(n_109), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_189), .B(n_123), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_170), .B(n_137), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_204), .B(n_186), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_224), .B(n_160), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_202), .A2(n_185), .B(n_190), .C(n_172), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_199), .B(n_190), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_210), .B(n_179), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_226), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_206), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_227), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_224), .B(n_173), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_226), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_208), .A2(n_172), .B(n_138), .C(n_143), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_192), .A2(n_143), .B(n_137), .C(n_129), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_217), .B(n_137), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_203), .Y(n_253) );
AND3x2_ASAP7_75t_L g254 ( .A(n_201), .B(n_121), .C(n_122), .Y(n_254) );
AND3x2_ASAP7_75t_L g255 ( .A(n_216), .B(n_9), .C(n_10), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_212), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_198), .A2(n_192), .B1(n_220), .B2(n_223), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_208), .A2(n_152), .B(n_150), .C(n_134), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_225), .A2(n_182), .B(n_184), .C(n_173), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
BUFx4f_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_233), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_218), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_218), .B(n_152), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_220), .B(n_152), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_214), .B(n_191), .Y(n_270) );
INVx6_ASAP7_75t_SL g271 ( .A(n_234), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_196), .A2(n_150), .B1(n_134), .B2(n_184), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_196), .B(n_134), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_233), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_233), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_219), .B(n_134), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_211), .B(n_10), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_195), .B(n_150), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_193), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_274), .A2(n_182), .B(n_200), .Y(n_281) );
OR2x6_ASAP7_75t_L g282 ( .A(n_280), .B(n_234), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_246), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_275), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_280), .A2(n_211), .B1(n_215), .B2(n_234), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_275), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_260), .A2(n_236), .B(n_229), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_246), .Y(n_288) );
OR3x4_ASAP7_75t_SL g289 ( .A(n_255), .B(n_216), .C(n_12), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_240), .A2(n_205), .B(n_221), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_275), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_251), .B(n_229), .C(n_194), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_242), .B(n_194), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_278), .A2(n_215), .B1(n_232), .B2(n_222), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_248), .A2(n_200), .B(n_205), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_238), .B(n_197), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_239), .B(n_231), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_250), .A2(n_221), .B(n_230), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_267), .B(n_235), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_275), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_261), .A2(n_209), .B(n_207), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_267), .Y(n_304) );
NOR2x1_ASAP7_75t_R g305 ( .A(n_239), .B(n_231), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_247), .B(n_231), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_253), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_239), .B(n_231), .Y(n_308) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_259), .A2(n_232), .B(n_225), .Y(n_309) );
AOI21x1_ASAP7_75t_L g310 ( .A1(n_273), .A2(n_150), .B(n_134), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_277), .A2(n_222), .B(n_150), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_253), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_277), .A2(n_222), .B(n_150), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_259), .A2(n_222), .B(n_150), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_258), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_290), .A2(n_279), .B(n_269), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_296), .B(n_252), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_282), .A2(n_271), .B1(n_263), .B2(n_243), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_290), .A2(n_269), .B(n_276), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_303), .A2(n_276), .B(n_268), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_285), .A2(n_241), .B1(n_249), .B2(n_263), .C(n_270), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_296), .A2(n_257), .B1(n_262), .B2(n_272), .C(n_263), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_309), .A2(n_271), .B1(n_254), .B2(n_222), .Y(n_326) );
OAI22xp33_ASAP7_75t_SL g327 ( .A1(n_282), .A2(n_271), .B1(n_262), .B2(n_257), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_296), .B(n_256), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_299), .B(n_256), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_299), .B(n_272), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_309), .A2(n_266), .B1(n_265), .B2(n_247), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_305), .A2(n_266), .B(n_237), .C(n_244), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_266), .B1(n_265), .B2(n_247), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_288), .B(n_245), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_292), .A2(n_245), .B(n_244), .C(n_237), .Y(n_336) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_315), .A2(n_268), .B(n_264), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_299), .B(n_264), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_309), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_282), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_282), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_282), .A2(n_16), .B1(n_18), .B2(n_19), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_297), .B(n_18), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_344), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_337), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_318), .B(n_304), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_340), .B(n_316), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_318), .B(n_328), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_340), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_323), .B(n_307), .Y(n_354) );
AO31x2_ASAP7_75t_L g355 ( .A1(n_320), .A2(n_284), .A3(n_286), .B(n_291), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_323), .B(n_312), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_340), .B(n_312), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_324), .B(n_287), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_313), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_329), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_329), .B(n_313), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_330), .B(n_282), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_332), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_343), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_335), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_321), .A2(n_315), .B(n_303), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_330), .B(n_315), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_333), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_338), .B(n_314), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_349), .A2(n_341), .B1(n_326), .B2(n_293), .C(n_339), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_369), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_373), .B(n_331), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_373), .B(n_334), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_350), .A2(n_325), .B1(n_333), .B2(n_319), .Y(n_381) );
NAND3xp33_ASAP7_75t_SL g382 ( .A(n_350), .B(n_345), .C(n_342), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_375), .B(n_338), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
AO21x2_ASAP7_75t_L g385 ( .A1(n_371), .A2(n_336), .B(n_317), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_374), .A2(n_322), .B1(n_325), .B2(n_319), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_371), .A2(n_327), .B(n_314), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_375), .B(n_351), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_374), .A2(n_322), .B1(n_294), .B2(n_292), .C(n_346), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_369), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_351), .B(n_287), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_352), .B(n_287), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_327), .B1(n_297), .B2(n_308), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_352), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_355), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g401 ( .A1(n_364), .A2(n_297), .B(n_308), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_366), .Y(n_402) );
AO21x2_ASAP7_75t_L g403 ( .A1(n_371), .A2(n_310), .B(n_303), .Y(n_403) );
INVx4_ASAP7_75t_L g404 ( .A(n_352), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_367), .B(n_368), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_349), .A2(n_302), .B1(n_289), .B2(n_297), .C(n_308), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_352), .B(n_287), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_360), .A2(n_302), .B1(n_305), .B2(n_284), .C(n_286), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_409), .B(n_348), .Y(n_411) );
AO21x1_ASAP7_75t_L g412 ( .A1(n_381), .A2(n_368), .B(n_357), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_409), .B(n_348), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_400), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_396), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_400), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_409), .B(n_353), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_389), .B(n_361), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_389), .B(n_392), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_404), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_392), .B(n_353), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_377), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_377), .B(n_358), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_379), .B(n_359), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_402), .B(n_358), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_383), .B(n_361), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_379), .B(n_359), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_383), .B(n_365), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_406), .B(n_360), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_402), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_409), .B(n_365), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_380), .B(n_361), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_398), .B(n_361), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_398), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_387), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_380), .B(n_371), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_404), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_405), .B(n_370), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_387), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_406), .B(n_357), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_380), .B(n_370), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_391), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_405), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_401), .B(n_370), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_380), .B(n_372), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_401), .B(n_372), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_386), .B(n_372), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_393), .B(n_355), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_400), .Y(n_460) );
INVxp33_ASAP7_75t_L g461 ( .A(n_381), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_421), .B(n_393), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_412), .B(n_404), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_421), .B(n_407), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_444), .B(n_407), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_444), .B(n_408), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_448), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_415), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_412), .B(n_422), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_461), .B(n_408), .Y(n_471) );
AOI211xp5_ASAP7_75t_L g472 ( .A1(n_434), .A2(n_410), .B(n_390), .C(n_376), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
NAND4xp75_ASAP7_75t_L g474 ( .A(n_449), .B(n_376), .C(n_388), .D(n_356), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_425), .B(n_410), .C(n_395), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_459), .B(n_408), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_459), .B(n_385), .Y(n_478) );
OAI31xp33_ASAP7_75t_L g479 ( .A1(n_422), .A2(n_390), .A3(n_297), .B(n_308), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_436), .Y(n_480) );
NOR2xp67_ASAP7_75t_SL g481 ( .A(n_445), .B(n_388), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_429), .B(n_354), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_414), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g484 ( .A1(n_445), .A2(n_455), .B(n_458), .C(n_457), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_417), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_450), .B(n_385), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_420), .B(n_19), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_450), .B(n_385), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_433), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_423), .B(n_438), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_424), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_416), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_416), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_423), .B(n_385), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_440), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_429), .B(n_356), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_432), .B(n_354), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_438), .B(n_403), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_411), .B(n_403), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_428), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_441), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_456), .B(n_403), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_428), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_424), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_426), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_443), .B(n_403), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_433), .B(n_355), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_456), .B(n_355), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_432), .B(n_453), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_418), .B(n_287), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_419), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_431), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_418), .B(n_363), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_460), .B(n_363), .C(n_298), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_430), .B(n_382), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_452), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_453), .B(n_382), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_418), .B(n_437), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_491), .B(n_430), .Y(n_522) );
OAI32xp33_ASAP7_75t_SL g523 ( .A1(n_475), .A2(n_454), .A3(n_439), .B1(n_442), .B2(n_446), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_505), .Y(n_524) );
XOR2x2_ASAP7_75t_L g525 ( .A(n_472), .B(n_442), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_519), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_497), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_491), .A2(n_451), .B1(n_447), .B2(n_443), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_502), .Y(n_529) );
OAI22xp33_ASAP7_75t_SL g530 ( .A1(n_470), .A2(n_451), .B1(n_447), .B2(n_460), .Y(n_530) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_484), .B(n_435), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_520), .B(n_437), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_469), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_492), .B(n_411), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_468), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_471), .B(n_437), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_512), .B(n_437), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_474), .A2(n_418), .B(n_419), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_479), .A2(n_411), .A3(n_413), .B(n_435), .Y(n_539) );
AND2x4_ASAP7_75t_SL g540 ( .A(n_480), .B(n_413), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_469), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_478), .B(n_416), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_489), .A2(n_413), .B1(n_411), .B2(n_308), .C(n_306), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_473), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_485), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_518), .B(n_413), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_492), .B(n_300), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_463), .A2(n_306), .B(n_301), .C(n_284), .Y(n_550) );
OAI32xp33_ASAP7_75t_L g551 ( .A1(n_518), .A2(n_306), .A3(n_300), .B1(n_291), .B2(n_286), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_516), .A2(n_314), .B1(n_311), .B2(n_300), .Y(n_552) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_508), .A2(n_310), .B(n_311), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_477), .A2(n_306), .B1(n_291), .B2(n_301), .C(n_26), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_514), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_478), .B(n_298), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_474), .A2(n_298), .B1(n_301), .B2(n_311), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_517), .B(n_298), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_462), .B(n_281), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_476), .B(n_281), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
OAI221xp5_ASAP7_75t_SL g564 ( .A1(n_515), .A2(n_496), .B1(n_510), .B2(n_504), .C(n_516), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_476), .B(n_298), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_467), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_482), .A2(n_281), .B1(n_22), .B2(n_24), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_496), .A2(n_295), .B1(n_29), .B2(n_30), .Y(n_568) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_508), .B(n_21), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_487), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_464), .B(n_33), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_501), .B(n_295), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_509), .A2(n_295), .B1(n_36), .B2(n_39), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_498), .B(n_34), .Y(n_574) );
NAND2x1_ASAP7_75t_SL g575 ( .A(n_531), .B(n_521), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_524), .B(n_500), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_530), .B(n_501), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_539), .A2(n_481), .B1(n_504), .B2(n_510), .C(n_499), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_566), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_533), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_535), .B(n_500), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_540), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_526), .B(n_521), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_541), .Y(n_584) );
XNOR2xp5_ASAP7_75t_L g585 ( .A(n_525), .B(n_466), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_539), .B(n_501), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_523), .A2(n_564), .B1(n_528), .B2(n_563), .C(n_527), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_529), .B(n_466), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_529), .B(n_542), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_550), .A2(n_481), .B(n_509), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_538), .B(n_493), .C(n_511), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_544), .B(n_467), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_534), .B(n_465), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_543), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_542), .B(n_465), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_538), .B(n_494), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_522), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_559), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_548), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_549), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_560), .Y(n_603) );
OAI322xp33_ASAP7_75t_L g604 ( .A1(n_547), .A2(n_511), .A3(n_507), .B1(n_506), .B2(n_493), .C1(n_486), .C2(n_490), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_SL g605 ( .A1(n_572), .A2(n_506), .B(n_507), .C(n_494), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_537), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_532), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_554), .A2(n_490), .B(n_486), .Y(n_609) );
NAND2xp33_ASAP7_75t_L g610 ( .A(n_569), .B(n_513), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_582), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_587), .B(n_571), .C(n_555), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_604), .A2(n_536), .B1(n_556), .B2(n_567), .C(n_574), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_577), .A2(n_556), .B1(n_567), .B2(n_551), .C(n_565), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_585), .B(n_561), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_579), .Y(n_617) );
XNOR2x1_ASAP7_75t_L g618 ( .A(n_601), .B(n_513), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_586), .B(n_577), .C(n_578), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_580), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_584), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_584), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_599), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_586), .A2(n_558), .B(n_573), .Y(n_625) );
OAI21xp33_ASAP7_75t_SL g626 ( .A1(n_597), .A2(n_557), .B(n_553), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_590), .A2(n_592), .B1(n_609), .B2(n_591), .C(n_597), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_592), .A2(n_552), .B(n_568), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_595), .Y(n_629) );
AO21x1_ASAP7_75t_L g630 ( .A1(n_610), .A2(n_495), .B(n_488), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_608), .B(n_562), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_598), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_619), .A2(n_581), .B1(n_589), .B2(n_607), .C1(n_588), .C2(n_583), .Y(n_633) );
NOR2xp33_ASAP7_75t_R g634 ( .A(n_624), .B(n_583), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_627), .A2(n_605), .B1(n_576), .B2(n_603), .C(n_600), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_626), .A2(n_606), .B1(n_602), .B2(n_579), .C1(n_593), .C2(n_495), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_628), .A2(n_605), .B(n_596), .C(n_488), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_616), .A2(n_483), .B1(n_41), .B2(n_42), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_620), .Y(n_639) );
NAND2xp33_ASAP7_75t_R g640 ( .A(n_612), .B(n_40), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_623), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_625), .A2(n_483), .B(n_49), .C(n_53), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_611), .B(n_44), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_613), .A2(n_54), .B1(n_56), .B2(n_57), .C(n_59), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_616), .A2(n_60), .B1(n_61), .B2(n_62), .C(n_65), .Y(n_645) );
AOI211xp5_ASAP7_75t_SL g646 ( .A1(n_644), .A2(n_615), .B(n_614), .C(n_621), .Y(n_646) );
OR5x1_ASAP7_75t_L g647 ( .A(n_636), .B(n_618), .C(n_630), .D(n_622), .E(n_621), .Y(n_647) );
AND3x4_ASAP7_75t_L g648 ( .A(n_634), .B(n_631), .C(n_622), .Y(n_648) );
NAND4xp25_ASAP7_75t_SL g649 ( .A(n_635), .B(n_632), .C(n_629), .D(n_617), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_633), .B(n_617), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_637), .B(n_66), .C(n_67), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_639), .A2(n_69), .B1(n_70), .B2(n_71), .Y(n_652) );
OAI211xp5_ASAP7_75t_SL g653 ( .A1(n_646), .A2(n_645), .B(n_638), .C(n_642), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_648), .A2(n_640), .B1(n_643), .B2(n_641), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_650), .B(n_72), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_649), .B(n_651), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_655), .Y(n_657) );
NAND2x1_ASAP7_75t_L g658 ( .A(n_654), .B(n_647), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_656), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_658), .A2(n_653), .B1(n_652), .B2(n_76), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_659), .B(n_74), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_661), .Y(n_662) );
AOI32xp33_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_660), .A3(n_657), .B1(n_78), .B2(n_79), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_75), .A3(n_77), .B1(n_80), .B2(n_82), .C1(n_83), .C2(n_84), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_664), .A2(n_85), .B(n_87), .Y(n_665) );
endmodule