module fake_jpeg_23729_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_22),
.Y(n_26)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_18),
.B1(n_10),
.B2(n_12),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.C(n_24),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_9),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_19),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_43),
.B(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_22),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_19),
.B1(n_11),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_33),
.B1(n_20),
.B2(n_18),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_11),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_43),
.B1(n_20),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_17),
.B1(n_10),
.B2(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_21),
.B(n_14),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_53),
.B2(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_0),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_8),
.C(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_74),
.Y(n_80)
);

XOR2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_64),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_68),
.B1(n_76),
.B2(n_57),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_78),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_77),
.B1(n_48),
.B2(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_77),
.C(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_81),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_94),
.B1(n_89),
.B2(n_5),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_82),
.B1(n_80),
.B2(n_3),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_90),
.C(n_86),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_92),
.B(n_5),
.Y(n_103)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_96),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_98),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_99),
.C(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B1(n_101),
.B2(n_99),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_4),
.C(n_6),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_4),
.C(n_7),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_7),
.Y(n_109)
);


endmodule