module fake_jpeg_16596_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_0),
.Y(n_81)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_60),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_63),
.C(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_79),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_59),
.B1(n_62),
.B2(n_45),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_57),
.B1(n_46),
.B2(n_52),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_55),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_44),
.B1(n_56),
.B2(n_3),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_75),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_84),
.B1(n_80),
.B2(n_4),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_106),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_87),
.B1(n_88),
.B2(n_82),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_107),
.A2(n_101),
.B(n_2),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_1),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_10),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_11),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_13),
.C(n_18),
.Y(n_118)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_37),
.B(n_22),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_21),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_32),
.CI(n_30),
.CON(n_122),
.SN(n_122)
);


endmodule