module fake_jpeg_28167_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

OR2x2_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_9),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_28),
.C(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_14),
.B1(n_19),
.B2(n_21),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_24),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_23),
.B1(n_29),
.B2(n_27),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_55),
.B1(n_57),
.B2(n_22),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_24),
.B(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_50),
.Y(n_62)
);

NAND5xp2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_37),
.C(n_36),
.D(n_24),
.E(n_25),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.C(n_59),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_16),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_54),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_13),
.B1(n_21),
.B2(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_13),
.B(n_12),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_41),
.B1(n_44),
.B2(n_59),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_4),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_43),
.C(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_76),
.C(n_77),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_61),
.C(n_71),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_53),
.C(n_48),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_58),
.C(n_47),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_46),
.B1(n_56),
.B2(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_80),
.B(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_62),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.C(n_73),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_62),
.B(n_69),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.C(n_20),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_83),
.B(n_68),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_73),
.C(n_75),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_91),
.B(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_68),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_97),
.B(n_8),
.C(n_10),
.D(n_6),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);


endmodule