module fake_jpeg_23091_n_136 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx5_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_30),
.A2(n_13),
.B1(n_15),
.B2(n_21),
.Y(n_31)
);

BUFx2_ASAP7_75t_SL g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_11),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_21),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_20),
.B1(n_17),
.B2(n_12),
.Y(n_38)
);

AO22x2_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_28),
.B1(n_22),
.B2(n_13),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_53),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_13),
.B1(n_41),
.B2(n_33),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_28),
.C(n_29),
.Y(n_48)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_42),
.B(n_28),
.C(n_36),
.D(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_22),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_63),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_38),
.B(n_36),
.C(n_33),
.D(n_32),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_48),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_20),
.C(n_17),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_40),
.B1(n_45),
.B2(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_55),
.B(n_59),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_82),
.B(n_91),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_60),
.B(n_61),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_33),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_73),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_67),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_6),
.C(n_9),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_74),
.B1(n_78),
.B2(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_95),
.B1(n_99),
.B2(n_88),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_75),
.C(n_77),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_4),
.C(n_9),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_84),
.B1(n_83),
.B2(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_11),
.B1(n_14),
.B2(n_18),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_27),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_25),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_109),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_3),
.Y(n_116)
);

OAI22x1_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_91),
.B1(n_39),
.B2(n_16),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_18),
.B(n_14),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_7),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_12),
.B1(n_16),
.B2(n_39),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_110),
.C(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_25),
.Y(n_109)
);

AOI321xp33_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_92),
.A3(n_96),
.B1(n_94),
.B2(n_100),
.C(n_102),
.Y(n_112)
);

OAI21x1_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_3),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_116),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_102),
.B1(n_4),
.B2(n_3),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_108),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_124),
.B(n_118),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_112),
.B(n_7),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_7),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_118),
.C(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_8),
.B(n_10),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_8),
.C(n_10),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_123),
.B(n_1),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_133),
.B(n_134),
.C(n_132),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_130),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_2),
.Y(n_136)
);


endmodule