module fake_jpeg_6746_n_285 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_39),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_18),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_54),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_17),
.B1(n_19),
.B2(n_39),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_37),
.B1(n_39),
.B2(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_86),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_34),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_107),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_37),
.B1(n_46),
.B2(n_43),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_105),
.B1(n_89),
.B2(n_70),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_97),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_66),
.C(n_57),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_98),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_43),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_58),
.B(n_55),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_67),
.B(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_44),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_109),
.B(n_113),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_45),
.B1(n_65),
.B2(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_76),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_26),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_30),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_30),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_29),
.B(n_27),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_124),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_134),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_77),
.B1(n_71),
.B2(n_72),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_74),
.Y(n_136)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_113),
.B1(n_94),
.B2(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_149),
.Y(n_169)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_93),
.C(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_152),
.C(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_120),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_94),
.B1(n_98),
.B2(n_109),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_137),
.B1(n_131),
.B2(n_125),
.Y(n_174)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_94),
.C(n_92),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_111),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_99),
.B(n_113),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_164),
.B(n_139),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_112),
.C(n_63),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_101),
.C(n_28),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_101),
.B(n_86),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_166),
.Y(n_192)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_172),
.B(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_115),
.B(n_121),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_121),
.B(n_135),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_174),
.A2(n_175),
.B1(n_158),
.B2(n_156),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_133),
.B1(n_125),
.B2(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_181),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_187),
.B(n_188),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_26),
.B(n_23),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_143),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_162),
.C(n_146),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_22),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_156),
.B1(n_149),
.B2(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_206),
.B1(n_23),
.B2(n_21),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_177),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_152),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.C(n_203),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_207),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_157),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_170),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_167),
.B(n_13),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_84),
.B1(n_73),
.B2(n_28),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_219),
.Y(n_228)
);

AO21x2_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_168),
.B(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_221),
.B1(n_191),
.B2(n_206),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_198),
.B(n_167),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_223),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_227),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_176),
.B(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_217),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_187),
.B(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_179),
.B1(n_177),
.B2(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_74),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_190),
.C(n_203),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_24),
.B(n_2),
.C(n_3),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_84),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_25),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_1),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_21),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_197),
.B(n_193),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_235),
.B(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_215),
.C(n_227),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_192),
.B1(n_32),
.B2(n_25),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_32),
.B1(n_24),
.B2(n_15),
.Y(n_236)
);

BUFx12_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_242),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_251),
.B(n_3),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_1),
.B(n_2),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_254),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_24),
.C(n_14),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_240),
.B1(n_239),
.B2(n_237),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_235),
.B1(n_228),
.B2(n_24),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_14),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_237),
.B1(n_234),
.B2(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_255),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_13),
.B(n_3),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_261),
.A2(n_263),
.B(n_251),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_2),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_244),
.C(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_270),
.C(n_4),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_253),
.B1(n_5),
.B2(n_7),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_256),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_272),
.B(n_275),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_259),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_9),
.C(n_10),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_266),
.C(n_10),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_9),
.B(n_11),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_274),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_281),
.B(n_277),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_282),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_11),
.C(n_12),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_12),
.B(n_256),
.Y(n_285)
);


endmodule