module real_jpeg_941_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_28),
.B1(n_31),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_121)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_7),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_7),
.B(n_22),
.C(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_33),
.B1(n_55),
.B2(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_33),
.B1(n_42),
.B2(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_7),
.B(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_7),
.B(n_39),
.C(n_42),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_53),
.C(n_56),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_95),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_54),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_75),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_66),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_15),
.B(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_61),
.B2(n_62),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.C(n_47),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_18),
.A2(n_19),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_18),
.A2(n_19),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

AOI211xp5_ASAP7_75t_SL g108 ( 
.A1(n_18),
.A2(n_104),
.B(n_109),
.C(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_18),
.B(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_18),
.A2(n_19),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_18),
.A2(n_19),
.B1(n_200),
.B2(n_205),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_18),
.A2(n_19),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_18),
.A2(n_205),
.B(n_216),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_18),
.A2(n_19),
.B1(n_67),
.B2(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_67),
.C(n_71),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_48),
.C(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_19),
.B(n_86),
.Y(n_109)
);

AO21x2_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_32),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_20),
.A2(n_27),
.B1(n_32),
.B2(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_90),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_27),
.Y(n_135)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_28),
.B(n_149),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_34),
.A2(n_47),
.B1(n_48),
.B2(n_70),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_45),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_73),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_41),
.B(n_45),
.Y(n_63)
);

AO21x2_ASAP7_75t_SL g86 ( 
.A1(n_37),
.A2(n_41),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);

OA22x2_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_41),
.Y(n_166)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_44),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_42),
.B(n_160),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_47),
.A2(n_48),
.B1(n_72),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_59),
.B(n_60),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_49),
.A2(n_59),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_54),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_50),
.A2(n_54),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_95),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_56),
.B(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_67),
.Y(n_245)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_71),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_72),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_230),
.B(n_247),
.Y(n_75)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_210),
.B(n_229),
.Y(n_76)
);

AOI21x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_190),
.B(n_209),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_137),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_123),
.B(n_136),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_SL g137 ( 
.A(n_80),
.B(n_138),
.C(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_111),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_98),
.C(n_107),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_97),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_84),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_83),
.A2(n_84),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_86),
.B1(n_103),
.B2(n_104),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_86),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_85),
.A2(n_104),
.B(n_110),
.C(n_181),
.Y(n_184)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_103),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_92),
.C(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_86),
.A2(n_222),
.B(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_86),
.B(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_92),
.B1(n_134),
.B2(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_92),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_91),
.B(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_91),
.A2(n_92),
.B1(n_147),
.B2(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_92),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_92),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_92),
.B(n_103),
.C(n_165),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_94),
.B(n_121),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_107),
.B1(n_108),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_104),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_104),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_142),
.C(n_146),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_104),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_103),
.A2(n_104),
.B1(n_158),
.B2(n_159),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_103),
.A2(n_104),
.B1(n_146),
.B2(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_104),
.B(n_120),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_116),
.C(n_119),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_113),
.A2(n_114),
.B(n_117),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_113),
.A2(n_114),
.B(n_197),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_127),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_133),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_129),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_130),
.A2(n_131),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_153),
.B(n_189),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_150),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_183),
.B(n_188),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_177),
.B(n_182),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_167),
.B(n_176),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_179),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_192),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_208),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_199),
.B1(n_206),
.B2(n_207),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_206),
.C(n_208),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_205),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_202),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_212),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_220),
.B2(n_221),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_220),
.C(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_234),
.B1(n_235),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_242),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_241),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_239),
.C(n_240),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_246),
.Y(n_249)
);


endmodule