module fake_ariane_2505_n_995 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_995);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_995;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_222;
wire n_703;
wire n_478;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_727;
wire n_699;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_288;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_52),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_6),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_93),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_187),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_58),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_22),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_97),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_149),
.Y(n_205)
);

BUFx8_ASAP7_75t_SL g206 ( 
.A(n_111),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_36),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_67),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_143),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_165),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_8),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_92),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_13),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_152),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_22),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_155),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_73),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_6),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_39),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_138),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_68),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_186),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_14),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_175),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_188),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_64),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_79),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_118),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_70),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_82),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_43),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

BUFx2_ASAP7_75t_SL g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_145),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_15),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_1),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_125),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_122),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_78),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_121),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_182),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_28),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_61),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_150),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_80),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_46),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_87),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_66),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_21),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_51),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_160),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_13),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_139),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_181),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_72),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_237),
.Y(n_280)
);

BUFx8_ASAP7_75t_SL g281 ( 
.A(n_272),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_202),
.B(n_0),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

BUFx8_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

CKINVDCx11_ASAP7_75t_R g286 ( 
.A(n_234),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_194),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g292 ( 
.A(n_224),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_194),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_38),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_206),
.B(n_40),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_208),
.B(n_0),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_198),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_214),
.B(n_1),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_215),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_226),
.B(n_2),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_210),
.B(n_2),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_3),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_241),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_213),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_191),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_266),
.B(n_4),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

BUFx8_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_223),
.B(n_231),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_218),
.B(n_5),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_238),
.B(n_5),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_7),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_193),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_250),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_251),
.B(n_7),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_260),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_278),
.B1(n_234),
.B2(n_244),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_308),
.A2(n_261),
.B1(n_270),
.B2(n_276),
.Y(n_335)
);

AO22x2_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_247),
.B1(n_278),
.B2(n_244),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_195),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_277),
.B1(n_273),
.B2(n_268),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_196),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_267),
.B1(n_264),
.B2(n_262),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_259),
.B1(n_258),
.B2(n_256),
.Y(n_342)
);

AO22x2_ASAP7_75t_L g343 ( 
.A1(n_280),
.A2(n_206),
.B1(n_9),
.B2(n_10),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

AO22x2_ASAP7_75t_L g345 ( 
.A1(n_280),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_255),
.B1(n_254),
.B2(n_245),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_292),
.A2(n_240),
.B1(n_239),
.B2(n_197),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_R g353 ( 
.A1(n_302),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_283),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_327),
.B1(n_332),
.B2(n_325),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_204),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_291),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_294),
.B(n_205),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_221),
.B1(n_236),
.B2(n_233),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_305),
.A2(n_207),
.B1(n_209),
.B2(n_211),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_324),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g365 ( 
.A1(n_304),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_229),
.B1(n_228),
.B2(n_227),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_R g367 ( 
.A1(n_307),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_R g368 ( 
.A1(n_281),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_316),
.A2(n_225),
.B1(n_222),
.B2(n_219),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_312),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_316),
.A2(n_238),
.B1(n_17),
.B2(n_18),
.Y(n_371)
);

OR2x6_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_16),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_310),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_324),
.A2(n_238),
.B1(n_20),
.B2(n_23),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_322),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_324),
.A2(n_238),
.B1(n_26),
.B2(n_27),
.Y(n_377)
);

BUFx6f_ASAP7_75t_SL g378 ( 
.A(n_301),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_320),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_320),
.B(n_238),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_321),
.B(n_238),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

OA22x2_ASAP7_75t_L g383 ( 
.A1(n_312),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_323),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_323),
.B(n_31),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_303),
.B(n_32),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_330),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_321),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_321),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_339),
.B(n_330),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_334),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_336),
.B(n_286),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

AOI21x1_ASAP7_75t_L g407 ( 
.A1(n_381),
.A2(n_328),
.B(n_326),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_373),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_337),
.B(n_303),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_358),
.A2(n_326),
.B(n_297),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_359),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_339),
.B(n_303),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_340),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_378),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

BUFx6f_ASAP7_75t_SL g419 ( 
.A(n_372),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_336),
.B(n_285),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_338),
.B(n_330),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_330),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_383),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_295),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

OR2x6_ASAP7_75t_L g430 ( 
.A(n_343),
.B(n_295),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_345),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_377),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_371),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_369),
.B(n_306),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_364),
.B(n_311),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_374),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_346),
.B(n_296),
.Y(n_442)
);

XNOR2x2_ASAP7_75t_L g443 ( 
.A(n_355),
.B(n_301),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_352),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_379),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_354),
.B(n_342),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_335),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_353),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_367),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_368),
.B(n_311),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_336),
.B(n_306),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_348),
.Y(n_459)
);

XOR2x2_ASAP7_75t_L g460 ( 
.A(n_334),
.B(n_35),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_336),
.B(n_306),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_300),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_391),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_409),
.B(n_318),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_414),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_408),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_300),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_431),
.B(n_318),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_428),
.B(n_319),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_416),
.B(n_319),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_296),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_441),
.B(n_296),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_433),
.B(n_309),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_400),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_400),
.Y(n_484)
);

AND2x6_ASAP7_75t_SL g485 ( 
.A(n_452),
.B(n_282),
.Y(n_485)
);

BUFx5_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_428),
.B(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_428),
.B(n_309),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_412),
.B(n_296),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_430),
.B(n_309),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_393),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_414),
.B(n_440),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_426),
.B(n_296),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_426),
.B(n_296),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_443),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_309),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_456),
.B(n_309),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_461),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_463),
.B(n_314),
.Y(n_511)
);

AND2x2_ASAP7_75t_SL g512 ( 
.A(n_447),
.B(n_300),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_447),
.B(n_300),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_423),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_446),
.A2(n_297),
.B1(n_314),
.B2(n_300),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_396),
.B(n_314),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_396),
.B(n_314),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_427),
.B(n_314),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_418),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_289),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_423),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_444),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_446),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_425),
.B(n_298),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_436),
.B(n_297),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_444),
.B(n_290),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_454),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_429),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_390),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_395),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_435),
.B(n_282),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_442),
.B(n_293),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_482),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_442),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_495),
.B(n_445),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_495),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_497),
.B(n_445),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_543),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_482),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_495),
.B(n_417),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_548),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_531),
.B(n_453),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_495),
.B(n_401),
.Y(n_560)
);

CKINVDCx6p67_ASAP7_75t_R g561 ( 
.A(n_535),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_531),
.B(n_451),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_462),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_482),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_527),
.Y(n_566)
);

NOR2x1_ASAP7_75t_L g567 ( 
.A(n_535),
.B(n_457),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_545),
.B(n_460),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_487),
.B(n_535),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_540),
.B(n_460),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_401),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_487),
.B(n_403),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_497),
.B(n_293),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_470),
.B(n_455),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_529),
.B(n_455),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_510),
.B(n_420),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_505),
.B(n_297),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_497),
.B(n_297),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_543),
.B(n_298),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_543),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_530),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_505),
.B(n_297),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_543),
.B(n_298),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_539),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_474),
.B(n_297),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_529),
.B(n_290),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_543),
.B(n_298),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_533),
.B(n_493),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_542),
.B(n_298),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_512),
.B(n_514),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_466),
.B(n_290),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_467),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_510),
.B(n_287),
.Y(n_602)
);

BUFx8_ASAP7_75t_SL g603 ( 
.A(n_542),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_506),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_469),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_530),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_473),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_474),
.B(n_42),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_542),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_498),
.B(n_287),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_520),
.B(n_287),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_539),
.B(n_287),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_506),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_506),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_502),
.B(n_44),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_569),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_599),
.B(n_486),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_566),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_586),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_595),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_595),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_591),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_571),
.Y(n_624)
);

BUFx6f_ASAP7_75t_SL g625 ( 
.A(n_560),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_558),
.Y(n_626)
);

INVx8_ASAP7_75t_L g627 ( 
.A(n_595),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_576),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_609),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_553),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_559),
.B(n_468),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_602),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_615),
.B(n_481),
.Y(n_634)
);

BUFx8_ASAP7_75t_L g635 ( 
.A(n_562),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

INVx5_ASAP7_75t_SL g637 ( 
.A(n_561),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_604),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_611),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_582),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_570),
.B(n_502),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_578),
.B(n_468),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_601),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx6_ASAP7_75t_L g645 ( 
.A(n_579),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_570),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_550),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_566),
.Y(n_648)
);

CKINVDCx6p67_ASAP7_75t_R g649 ( 
.A(n_570),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_578),
.B(n_528),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_551),
.A2(n_484),
.B1(n_483),
.B2(n_563),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_552),
.B(n_557),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_603),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_550),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_557),
.Y(n_655)
);

BUFx12f_ASAP7_75t_L g656 ( 
.A(n_560),
.Y(n_656)
);

BUFx2_ASAP7_75t_SL g657 ( 
.A(n_608),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_556),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_604),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_608),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_579),
.B(n_607),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_605),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_568),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_556),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_573),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_605),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_552),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_595),
.A2(n_469),
.B1(n_502),
.B2(n_517),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_580),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_568),
.B(n_528),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_552),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_573),
.B(n_502),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_588),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_556),
.Y(n_674)
);

CKINVDCx9p33_ASAP7_75t_R g675 ( 
.A(n_660),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_627),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_657),
.A2(n_599),
.B1(n_572),
.B2(n_581),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_635),
.A2(n_548),
.B1(n_512),
.B2(n_514),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_648),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_670),
.B(n_534),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_628),
.A2(n_548),
.B1(n_564),
.B2(n_541),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_663),
.A2(n_548),
.B1(n_564),
.B2(n_541),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_665),
.A2(n_541),
.B1(n_537),
.B2(n_574),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_669),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_616),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_619),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_616),
.Y(n_688)
);

BUFx12f_ASAP7_75t_L g689 ( 
.A(n_635),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_669),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_625),
.A2(n_537),
.B1(n_574),
.B2(n_512),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_673),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_640),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_640),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_625),
.A2(n_537),
.B1(n_574),
.B2(n_514),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_643),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_673),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_625),
.A2(n_567),
.B1(n_473),
.B2(n_551),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_643),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_634),
.A2(n_546),
.B1(n_606),
.B2(n_615),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_635),
.A2(n_473),
.B1(n_486),
.B2(n_534),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_656),
.A2(n_473),
.B1(n_486),
.B2(n_521),
.Y(n_702)
);

CKINVDCx14_ASAP7_75t_R g703 ( 
.A(n_653),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_627),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_632),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_627),
.Y(n_706)
);

CKINVDCx11_ASAP7_75t_R g707 ( 
.A(n_653),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_624),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_656),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_655),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_662),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_666),
.Y(n_712)
);

BUFx12f_ASAP7_75t_L g713 ( 
.A(n_623),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_634),
.A2(n_642),
.B1(n_650),
.B2(n_631),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_623),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_672),
.A2(n_473),
.B1(n_486),
.B2(n_521),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_634),
.A2(n_583),
.B1(n_589),
.B2(n_539),
.Y(n_717)
);

BUFx2_ASAP7_75t_R g718 ( 
.A(n_671),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_627),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_634),
.A2(n_546),
.B1(n_600),
.B2(n_575),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_626),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_651),
.A2(n_600),
.B1(n_575),
.B2(n_544),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_633),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_639),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_641),
.A2(n_473),
.B1(n_486),
.B2(n_522),
.Y(n_725)
);

BUFx4_ASAP7_75t_SL g726 ( 
.A(n_626),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_641),
.A2(n_473),
.B1(n_486),
.B2(n_522),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_621),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_687),
.B(n_655),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

AOI222xp33_ASAP7_75t_L g731 ( 
.A1(n_691),
.A2(n_547),
.B1(n_641),
.B2(n_525),
.C1(n_485),
.C2(n_652),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_677),
.A2(n_509),
.B1(n_549),
.B2(n_547),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_678),
.A2(n_509),
.B1(n_549),
.B2(n_501),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_700),
.A2(n_668),
.B1(n_645),
.B2(n_637),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_695),
.A2(n_501),
.B1(n_489),
.B2(n_500),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_724),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_679),
.B(n_493),
.Y(n_737)
);

CKINVDCx14_ASAP7_75t_R g738 ( 
.A(n_703),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_675),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_SL g740 ( 
.A1(n_714),
.A2(n_477),
.B(n_652),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_720),
.A2(n_652),
.B1(n_621),
.B2(n_622),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_684),
.A2(n_479),
.B1(n_486),
.B2(n_621),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_721),
.A2(n_722),
.B1(n_683),
.B2(n_708),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_682),
.A2(n_486),
.B1(n_622),
.B2(n_491),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_689),
.Y(n_745)
);

OAI21xp33_ASAP7_75t_L g746 ( 
.A1(n_681),
.A2(n_476),
.B(n_508),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_689),
.A2(n_649),
.B1(n_555),
.B2(n_607),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_708),
.A2(n_645),
.B1(n_637),
.B2(n_618),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_724),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_698),
.A2(n_486),
.B1(n_492),
.B2(n_491),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_687),
.B(n_485),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_710),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_705),
.A2(n_500),
.B1(n_489),
.B2(n_492),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_717),
.A2(n_491),
.B1(n_492),
.B2(n_525),
.Y(n_755)
);

OAI222xp33_ASAP7_75t_L g756 ( 
.A1(n_705),
.A2(n_671),
.B1(n_555),
.B2(n_519),
.C1(n_667),
.C2(n_496),
.Y(n_756)
);

BUFx4f_ASAP7_75t_SL g757 ( 
.A(n_713),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_709),
.A2(n_508),
.B1(n_511),
.B2(n_488),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_711),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_709),
.A2(n_511),
.B1(n_471),
.B2(n_488),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_701),
.B(n_617),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_711),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_SL g763 ( 
.A1(n_702),
.A2(n_496),
.B(n_618),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_716),
.A2(n_645),
.B1(n_637),
.B2(n_659),
.Y(n_764)
);

AOI21xp33_ASAP7_75t_L g765 ( 
.A1(n_685),
.A2(n_507),
.B(n_524),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_685),
.A2(n_471),
.B1(n_478),
.B2(n_475),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_712),
.B(n_636),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_676),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_710),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_690),
.A2(n_478),
.B1(n_475),
.B2(n_480),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_725),
.A2(n_637),
.B1(n_638),
.B2(n_644),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_690),
.Y(n_772)
);

INVx3_ASAP7_75t_SL g773 ( 
.A(n_715),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_692),
.A2(n_480),
.B1(n_646),
.B2(n_481),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_680),
.A2(n_481),
.B1(n_607),
.B2(n_646),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_712),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_713),
.A2(n_649),
.B1(n_539),
.B2(n_481),
.Y(n_777)
);

BUFx8_ASAP7_75t_SL g778 ( 
.A(n_707),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_727),
.A2(n_644),
.B1(n_630),
.B2(n_607),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_676),
.Y(n_780)
);

INVx5_ASAP7_75t_SL g781 ( 
.A(n_726),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_728),
.A2(n_644),
.B1(n_630),
.B2(n_661),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_680),
.A2(n_524),
.B1(n_636),
.B2(n_610),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_692),
.A2(n_597),
.B1(n_536),
.B2(n_589),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_718),
.B(n_697),
.Y(n_785)
);

OAI21xp33_ASAP7_75t_L g786 ( 
.A1(n_723),
.A2(n_538),
.B(n_494),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_676),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_697),
.A2(n_592),
.B1(n_583),
.B2(n_544),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_706),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_706),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_740),
.B(n_723),
.C(n_593),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_743),
.B(n_593),
.C(n_554),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_739),
.A2(n_728),
.B1(n_719),
.B2(n_706),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_731),
.A2(n_704),
.B1(n_719),
.B2(n_688),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_732),
.A2(n_704),
.B1(n_719),
.B2(n_688),
.Y(n_795)
);

OAI221xp5_ASAP7_75t_L g796 ( 
.A1(n_752),
.A2(n_490),
.B1(n_523),
.B2(n_526),
.C(n_519),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_741),
.A2(n_728),
.B1(n_704),
.B2(n_490),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_732),
.A2(n_693),
.B1(n_699),
.B2(n_696),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_785),
.A2(n_704),
.B1(n_728),
.B2(n_699),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_759),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_729),
.B(n_686),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_763),
.A2(n_704),
.B1(n_490),
.B2(n_612),
.Y(n_802)
);

AOI222xp33_ASAP7_75t_L g803 ( 
.A1(n_756),
.A2(n_523),
.B1(n_533),
.B2(n_592),
.C1(n_597),
.C2(n_696),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_734),
.A2(n_694),
.B1(n_693),
.B2(n_686),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_735),
.A2(n_612),
.B1(n_617),
.B2(n_620),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_735),
.A2(n_612),
.B1(n_617),
.B2(n_620),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_736),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_733),
.A2(n_694),
.B1(n_544),
.B2(n_526),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_748),
.B(n_658),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_762),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_767),
.B(n_620),
.C(n_617),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_733),
.A2(n_758),
.B1(n_777),
.B2(n_760),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_750),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_746),
.A2(n_526),
.B1(n_513),
.B2(n_515),
.Y(n_814)
);

OAI222xp33_ASAP7_75t_L g815 ( 
.A1(n_761),
.A2(n_515),
.B1(n_513),
.B2(n_590),
.C1(n_465),
.C2(n_472),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_776),
.B(n_647),
.Y(n_816)
);

OAI222xp33_ASAP7_75t_L g817 ( 
.A1(n_783),
.A2(n_590),
.B1(n_465),
.B2(n_472),
.C1(n_674),
.C2(n_526),
.Y(n_817)
);

AOI221xp5_ASAP7_75t_L g818 ( 
.A1(n_754),
.A2(n_533),
.B1(n_504),
.B2(n_503),
.C(n_658),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_755),
.A2(n_613),
.B1(n_614),
.B2(n_536),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_SL g820 ( 
.A1(n_738),
.A2(n_661),
.B(n_620),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_754),
.A2(n_614),
.B1(n_613),
.B2(n_533),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_744),
.A2(n_647),
.B1(n_565),
.B2(n_587),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_730),
.A2(n_647),
.B1(n_565),
.B2(n_587),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_753),
.B(n_674),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_737),
.B(n_664),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_769),
.B(n_664),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_742),
.A2(n_516),
.B1(n_532),
.B2(n_584),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_730),
.B(n_633),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_772),
.B(n_633),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_749),
.A2(n_783),
.B1(n_764),
.B2(n_771),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_787),
.B(n_633),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_747),
.A2(n_584),
.B1(n_465),
.B2(n_472),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_SL g833 ( 
.A1(n_779),
.A2(n_598),
.B1(n_596),
.B2(n_654),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_757),
.A2(n_598),
.B1(n_596),
.B2(n_654),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_788),
.A2(n_516),
.B1(n_598),
.B2(n_596),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_751),
.A2(n_516),
.B1(n_518),
.B2(n_585),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_745),
.A2(n_518),
.B1(n_594),
.B2(n_585),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_789),
.B(n_654),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_812),
.A2(n_773),
.B1(n_790),
.B2(n_781),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_810),
.B(n_768),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_810),
.B(n_768),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_SL g842 ( 
.A(n_831),
.B(n_778),
.C(n_781),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_800),
.B(n_780),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_830),
.B(n_780),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_809),
.B(n_773),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_801),
.B(n_745),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_786),
.C(n_765),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_824),
.B(n_781),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_L g849 ( 
.A(n_811),
.B(n_784),
.C(n_775),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_794),
.A2(n_775),
.B1(n_774),
.B2(n_784),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_826),
.B(n_816),
.Y(n_851)
);

NAND4xp25_ASAP7_75t_L g852 ( 
.A(n_828),
.B(n_782),
.C(n_766),
.D(n_770),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_792),
.B(n_654),
.C(n_747),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_825),
.B(n_518),
.Y(n_854)
);

OAI221xp5_ASAP7_75t_L g855 ( 
.A1(n_794),
.A2(n_757),
.B1(n_594),
.B2(n_288),
.C(n_284),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_838),
.B(n_45),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_829),
.B(n_47),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_SL g858 ( 
.A(n_820),
.B(n_284),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_L g859 ( 
.A(n_818),
.B(n_796),
.C(n_799),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_SL g860 ( 
.A1(n_802),
.A2(n_49),
.B(n_50),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_795),
.B(n_288),
.C(n_284),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_807),
.B(n_53),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_793),
.B(n_54),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_833),
.B(n_284),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_804),
.B(n_55),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_795),
.B(n_56),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_797),
.B(n_57),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_798),
.B(n_59),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_834),
.B(n_60),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_823),
.B(n_817),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_837),
.B(n_814),
.C(n_808),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_819),
.B(n_62),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_837),
.B(n_288),
.C(n_284),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_803),
.A2(n_288),
.B1(n_284),
.B2(n_74),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_819),
.B(n_63),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_851),
.B(n_822),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_862),
.A2(n_805),
.B(n_806),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_847),
.B(n_827),
.C(n_835),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_875),
.A2(n_821),
.B1(n_832),
.B2(n_836),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_848),
.B(n_845),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_840),
.B(n_841),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_863),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_843),
.B(n_821),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_846),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_854),
.B(n_844),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_854),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_839),
.B(n_860),
.C(n_844),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_859),
.B(n_815),
.C(n_75),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_868),
.B(n_65),
.C(n_76),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_871),
.B(n_77),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_849),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_853),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_857),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_L g895 ( 
.A(n_871),
.B(n_288),
.C(n_83),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_856),
.B(n_81),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_864),
.B(n_84),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_882),
.B(n_842),
.Y(n_898)
);

XNOR2xp5_ASAP7_75t_L g899 ( 
.A(n_888),
.B(n_892),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_885),
.B(n_870),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_893),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_886),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_883),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_891),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_881),
.B(n_865),
.Y(n_905)
);

NAND4xp75_ASAP7_75t_L g906 ( 
.A(n_897),
.B(n_865),
.C(n_866),
.D(n_867),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_887),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_894),
.Y(n_908)
);

NAND4xp75_ASAP7_75t_L g909 ( 
.A(n_877),
.B(n_876),
.C(n_873),
.D(n_869),
.Y(n_909)
);

XNOR2xp5_ASAP7_75t_L g910 ( 
.A(n_879),
.B(n_875),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_884),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_901),
.B(n_877),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_901),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_911),
.Y(n_914)
);

XNOR2x1_ASAP7_75t_L g915 ( 
.A(n_899),
.B(n_896),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_908),
.B(n_878),
.Y(n_916)
);

XNOR2xp5_ASAP7_75t_L g917 ( 
.A(n_899),
.B(n_895),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_903),
.Y(n_918)
);

XNOR2xp5_ASAP7_75t_L g919 ( 
.A(n_910),
.B(n_880),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_918),
.Y(n_920)
);

XOR2x2_ASAP7_75t_L g921 ( 
.A(n_919),
.B(n_910),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_917),
.A2(n_909),
.B1(n_906),
.B2(n_904),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_915),
.Y(n_923)
);

OA22x2_ASAP7_75t_L g924 ( 
.A1(n_916),
.A2(n_911),
.B1(n_902),
.B2(n_898),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_916),
.A2(n_898),
.B1(n_905),
.B2(n_900),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_912),
.A2(n_909),
.B1(n_906),
.B2(n_889),
.Y(n_926)
);

BUFx2_ASAP7_75t_R g927 ( 
.A(n_923),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_926),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_920),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_925),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_922),
.Y(n_931)
);

OAI222xp33_ASAP7_75t_L g932 ( 
.A1(n_931),
.A2(n_924),
.B1(n_912),
.B2(n_914),
.C1(n_921),
.C2(n_900),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_928),
.A2(n_913),
.B1(n_905),
.B2(n_914),
.Y(n_933)
);

AOI221xp5_ASAP7_75t_L g934 ( 
.A1(n_931),
.A2(n_880),
.B1(n_890),
.B2(n_907),
.C(n_872),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_933),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_SL g936 ( 
.A1(n_932),
.A2(n_929),
.B(n_927),
.C(n_930),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_SL g937 ( 
.A1(n_934),
.A2(n_929),
.B(n_855),
.C(n_861),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_933),
.Y(n_938)
);

NOR2x1_ASAP7_75t_L g939 ( 
.A(n_938),
.B(n_874),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_935),
.A2(n_890),
.B1(n_878),
.B2(n_858),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_937),
.A2(n_852),
.B1(n_850),
.B2(n_288),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_936),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_938),
.B(n_850),
.Y(n_943)
);

NOR4xp25_ASAP7_75t_L g944 ( 
.A(n_938),
.B(n_86),
.C(n_88),
.D(n_90),
.Y(n_944)
);

AOI31xp33_ASAP7_75t_L g945 ( 
.A1(n_938),
.A2(n_91),
.A3(n_94),
.B(n_95),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_939),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_943),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_941),
.Y(n_948)
);

AO22x1_ASAP7_75t_L g949 ( 
.A1(n_942),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_945),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_940),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_944),
.Y(n_952)
);

OAI211xp5_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_105),
.B(n_107),
.C(n_108),
.Y(n_953)
);

NOR2xp67_ASAP7_75t_L g954 ( 
.A(n_950),
.B(n_109),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_946),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_SL g956 ( 
.A1(n_948),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_947),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_949),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_957),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_955),
.A2(n_951),
.B1(n_116),
.B2(n_117),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_958),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_954),
.A2(n_115),
.B1(n_124),
.B2(n_126),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_956),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_953),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_957),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_962),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_965),
.A2(n_961),
.B1(n_963),
.B2(n_964),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_959),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_960),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_970)
);

AO22x2_ASAP7_75t_L g971 ( 
.A1(n_966),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_959),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_962),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_959),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_959),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_975),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_972),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_974),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_968),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_971),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_967),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_980),
.A2(n_973),
.B1(n_970),
.B2(n_969),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_978),
.A2(n_190),
.B1(n_151),
.B2(n_153),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_977),
.A2(n_147),
.B1(n_154),
.B2(n_156),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_977),
.A2(n_189),
.B1(n_158),
.B2(n_159),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_982),
.Y(n_986)
);

XOR2x1_ASAP7_75t_L g987 ( 
.A(n_983),
.B(n_976),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_984),
.Y(n_988)
);

AO22x2_ASAP7_75t_L g989 ( 
.A1(n_986),
.A2(n_981),
.B1(n_979),
.B2(n_985),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_988),
.A2(n_981),
.B1(n_162),
.B2(n_164),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_987),
.A2(n_157),
.B1(n_166),
.B2(n_167),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_989),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_990),
.Y(n_993)
);

AOI221xp5_ASAP7_75t_L g994 ( 
.A1(n_992),
.A2(n_991),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_994)
);

AOI211xp5_ASAP7_75t_L g995 ( 
.A1(n_994),
.A2(n_993),
.B(n_173),
.C(n_176),
.Y(n_995)
);


endmodule