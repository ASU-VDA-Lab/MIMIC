module fake_jpeg_27163_n_40 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_1),
.B(n_0),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_5),
.B(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_19),
.B1(n_12),
.B2(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

OR2x4_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_19)
);

BUFx24_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_16),
.B1(n_22),
.B2(n_26),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

AOI221xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_19),
.B1(n_9),
.B2(n_11),
.C(n_8),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_13),
.C(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_11),
.Y(n_31)
);

AOI21x1_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_13),
.B(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_36),
.C(n_31),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.C(n_33),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_23),
.A3(n_25),
.B1(n_27),
.B2(n_35),
.C1(n_29),
.C2(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_23),
.Y(n_40)
);


endmodule