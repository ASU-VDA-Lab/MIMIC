module real_jpeg_33447_n_19 (n_17, n_8, n_0, n_141, n_2, n_139, n_142, n_143, n_10, n_137, n_9, n_12, n_146, n_6, n_136, n_11, n_14, n_138, n_7, n_18, n_3, n_145, n_144, n_5, n_4, n_1, n_140, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_141;
input n_2;
input n_139;
input n_142;
input n_143;
input n_10;
input n_137;
input n_9;
input n_12;
input n_146;
input n_6;
input n_136;
input n_11;
input n_14;
input n_138;
input n_7;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_1;
input n_140;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_0),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_95),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_2),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_4),
.A2(n_83),
.A3(n_85),
.B1(n_93),
.B2(n_115),
.C1(n_117),
.C2(n_146),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_7),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_14),
.B1(n_49),
.B2(n_53),
.C(n_57),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_9),
.B(n_49),
.C(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_11),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_100),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_12),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_13),
.B(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_16),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_16),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_133),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_123),
.B(n_130),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_32),
.B(n_121),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_24),
.B(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_39),
.B(n_120),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

AOI31xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_75),
.A3(n_105),
.B(n_110),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_69),
.C(n_70),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_61),
.B(n_68),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_138),
.Y(n_53)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_92),
.C(n_99),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_111),
.B(n_114),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_99),
.C(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_142),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OA21x2_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_136),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_137),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_139),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_140),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_141),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_143),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_144),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_145),
.Y(n_108)
);


endmodule