module fake_jpeg_9179_n_31 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_31);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_6),
.B1(n_1),
.B2(n_5),
.Y(n_17)
);

NAND2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_14),
.B1(n_0),
.B2(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_9),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_1),
.C(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_19),
.B2(n_16),
.Y(n_27)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_22),
.B(n_20),
.C(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_28),
.Y(n_30)
);

XNOR2x2_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_27),
.Y(n_31)
);


endmodule