module fake_jpeg_16365_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_5),
.C(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

OAI32xp33_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_28),
.A3(n_13),
.B1(n_17),
.B2(n_7),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_5),
.C(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_16),
.B1(n_19),
.B2(n_11),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_31),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_43),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_41),
.B1(n_30),
.B2(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_7),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_26),
.C(n_17),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_42),
.C(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_50),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_26),
.B(n_11),
.C(n_18),
.D(n_19),
.Y(n_46)
);

NOR2xp67_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_51),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_39),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_18),
.B(n_17),
.C(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_59),
.C(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_46),
.B1(n_52),
.B2(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_32),
.C(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_47),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

XOR2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_53),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_45),
.B1(n_51),
.B2(n_36),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_58),
.B(n_53),
.C(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_65),
.B1(n_66),
.B2(n_64),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_64),
.B1(n_69),
.B2(n_36),
.Y(n_72)
);


endmodule