module real_jpeg_11116_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_15),
.Y(n_25)
);

OA21x2_ASAP7_75t_L g10 ( 
.A1(n_2),
.A2(n_11),
.B(n_12),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_11),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_9),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g9 ( 
.A1(n_4),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_9)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_5),
.A2(n_10),
.B1(n_13),
.B2(n_16),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_15),
.B1(n_17),
.B2(n_21),
.C(n_22),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_24),
.Y(n_23)
);


endmodule