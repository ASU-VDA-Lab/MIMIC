module real_jpeg_6553_n_30 (n_17, n_8, n_0, n_21, n_168, n_2, n_29, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_28, n_171, n_169, n_162, n_167, n_23, n_11, n_14, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_29;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_28;
input n_171;
input n_169;
input n_162;
input n_167;
input n_23;
input n_11;
input n_14;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_0),
.B(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_1),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_2),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_3),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_54),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_5),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_44),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_6),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_6),
.B(n_146),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_7),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_60),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_8),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_9),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_12),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_12),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_33),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_16),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_16),
.B(n_106),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_17),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_18),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_20),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_21),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_50),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_91),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_26),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_26),
.B(n_143),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_28),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_29),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_29),
.B(n_128),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_154),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_153),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_35),
.B(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_141),
.B(n_150),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_121),
.B(n_135),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_64),
.B(n_109),
.C(n_118),
.Y(n_41)
);

NOR4xp25_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.C(n_53),
.D(n_59),
.Y(n_42)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_70),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_120),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_125),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_105),
.B(n_108),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_98),
.B(n_104),
.Y(n_65)
);

AO221x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_75),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B(n_94),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_79),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_93),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_89),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_103),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_144),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B(n_115),
.C(n_116),
.D(n_117),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_131),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_131),
.B(n_136),
.C(n_139),
.D(n_140),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_159),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_162),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_163),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_164),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_165),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_166),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_167),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_168),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_169),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_170),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_171),
.Y(n_107)
);


endmodule