module real_jpeg_23182_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_11),
.Y(n_13)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_5),
.A2(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_5),
.B(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_14),
.B(n_16),
.C(n_26),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_9),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_9),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_8),
.B(n_33),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_15),
.B1(n_32),
.B2(n_34),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_12),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_15),
.A2(n_20),
.B(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_21),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);


endmodule