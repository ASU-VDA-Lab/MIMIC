module fake_jpeg_4004_n_209 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_27),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_31),
.B1(n_20),
.B2(n_15),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_11),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_21),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_39),
.B1(n_41),
.B2(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_15),
.B1(n_13),
.B2(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_15),
.B1(n_20),
.B2(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_43),
.B1(n_19),
.B2(n_16),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_15),
.B1(n_13),
.B2(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_14),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_16),
.B1(n_19),
.B2(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_32),
.Y(n_45)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_21),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_51),
.A3(n_41),
.B1(n_37),
.B2(n_19),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_21),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_25),
.B(n_21),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_27),
.B1(n_31),
.B2(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_31),
.CON(n_89),
.SN(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_37),
.Y(n_72)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_35),
.B1(n_34),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_52),
.B1(n_47),
.B2(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_77),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_52),
.B1(n_35),
.B2(n_46),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_68),
.C(n_67),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_86),
.C(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_52),
.B1(n_35),
.B2(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_38),
.B(n_22),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_72),
.B(n_69),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_58),
.C(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_31),
.B1(n_12),
.B2(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_74),
.B1(n_69),
.B2(n_73),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_61),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.C(n_104),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_71),
.C(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_73),
.C(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_83),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_91),
.B1(n_102),
.B2(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_91),
.B1(n_88),
.B2(n_80),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

BUFx12f_ASAP7_75t_SL g112 ( 
.A(n_105),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_116),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_122),
.B(n_94),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_120),
.B(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_86),
.C(n_90),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_104),
.C(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_61),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_130),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_76),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_86),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_84),
.B1(n_80),
.B2(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_87),
.C(n_63),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_61),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_63),
.C(n_66),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_66),
.C(n_58),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_137),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_77),
.B1(n_33),
.B2(n_48),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_111),
.B(n_120),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_28),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_28),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_145),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_117),
.B(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_133),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_122),
.B1(n_108),
.B2(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_55),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_107),
.B(n_116),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_137),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_17),
.C(n_66),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_12),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_125),
.C(n_132),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_134),
.C(n_138),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_140),
.C(n_123),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_130),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

NAND2x1_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_58),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_75),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_75),
.C(n_17),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_155),
.B1(n_149),
.B2(n_33),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_44),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_151),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_175),
.B(n_33),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_33),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_152),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_7),
.B(n_11),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_155),
.C(n_75),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_0),
.C(n_1),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_55),
.B(n_8),
.C(n_9),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_33),
.B1(n_48),
.B2(n_44),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_0),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_33),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_0),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_187),
.B(n_177),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_172),
.C(n_9),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_188),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_180),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_200),
.C(n_2),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_2),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_181),
.B(n_9),
.C(n_8),
.D(n_7),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_201),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_0),
.B(n_1),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_189),
.C2(n_169),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_191),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_205),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_197),
.B(n_5),
.Y(n_206)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_202),
.B(n_5),
.C(n_6),
.D(n_4),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_207),
.Y(n_209)
);


endmodule