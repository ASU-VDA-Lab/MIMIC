module real_jpeg_11654_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_264, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_264;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_0),
.A2(n_46),
.B1(n_49),
.B2(n_61),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_0),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_127)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_5),
.A2(n_28),
.B1(n_46),
.B2(n_49),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_9),
.A2(n_46),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_38),
.B1(n_46),
.B2(n_49),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_10),
.A2(n_34),
.B(n_64),
.C(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_39),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_10),
.B(n_48),
.C(n_52),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_10),
.B(n_67),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_10),
.B(n_31),
.C(n_35),
.Y(n_206)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_110),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_109),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_78),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_16),
.B(n_78),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_70),
.B2(n_72),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_123),
.C(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_20),
.A2(n_21),
.B1(n_85),
.B2(n_159),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_20),
.A2(n_21),
.B1(n_123),
.B2(n_139),
.Y(n_250)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_21),
.B(n_85),
.C(n_217),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_23),
.A2(n_33),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_206),
.Y(n_205)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_29),
.B(n_39),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_35),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_38),
.A2(n_49),
.B(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_38),
.B(n_100),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_38),
.B(n_55),
.Y(n_187)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_58),
.B1(n_59),
.B2(n_69),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_70),
.C(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_69),
.B1(n_74),
.B2(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_55),
.B(n_56),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_43),
.A2(n_55),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_50),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_104),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_44),
.A2(n_50),
.B1(n_104),
.B2(n_129),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_46),
.B(n_169),
.Y(n_168)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_51),
.B(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_90),
.B(n_103),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_55),
.A2(n_103),
.B(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_67),
.B1(n_77),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_62),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_66),
.A2(n_76),
.B(n_87),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_66),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_70),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_72),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_70),
.A2(n_72),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_70),
.A2(n_72),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_72),
.B(n_123),
.C(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_72),
.B(n_227),
.C(n_232),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_77),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_92),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_85),
.B(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_85),
.A2(n_150),
.B1(n_151),
.B2(n_159),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_105),
.B(n_106),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_94),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_105),
.B1(n_106),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_95),
.A2(n_102),
.B1(n_105),
.B2(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_99),
.A2(n_100),
.B1(n_147),
.B2(n_156),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_100),
.A2(n_127),
.B(n_157),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_102),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_130),
.B(n_261),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_112),
.B(n_115),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_122),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_116),
.A2(n_120),
.B1(n_121),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_116),
.Y(n_259)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_122),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_123),
.A2(n_139),
.B1(n_140),
.B2(n_181),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_123),
.A2(n_139),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_124),
.A2(n_125),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_126),
.A2(n_128),
.B1(n_163),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_126),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_163),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_173),
.C(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_149),
.C(n_162),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_255),
.B(n_260),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_244),
.B(n_254),
.Y(n_133)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_214),
.A3(n_239),
.B1(n_242),
.B2(n_243),
.C(n_264),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_198),
.B(n_213),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_164),
.B(n_197),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_138),
.B(n_148),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.C(n_142),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_168),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_140),
.A2(n_181),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_142),
.A2(n_143),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_160),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_155),
.C(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_191),
.B(n_196),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_177),
.B(n_190),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_175),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_204),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_182),
.B(n_189),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_220),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_186),
.B(n_188),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_200),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_203),
.C(n_207),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_222),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_219),
.CI(n_222),
.CON(n_241),
.SN(n_241)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_238),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_235),
.B2(n_236),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_236),
.C(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_253),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_248),
.C(n_251),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);


endmodule