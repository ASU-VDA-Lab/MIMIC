module real_aes_1943_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_0), .A2(n_102), .B1(n_813), .B2(n_815), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_1), .B(n_498), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_2), .A2(n_500), .B(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_3), .B(n_821), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g106 ( .A1(n_4), .A2(n_5), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_4), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_5), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_6), .B(n_209), .Y(n_535) );
INVx1_ASAP7_75t_L g141 ( .A(n_7), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_8), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_9), .B(n_209), .Y(n_584) );
INVx1_ASAP7_75t_L g179 ( .A(n_10), .Y(n_179) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_11), .A2(n_105), .B1(n_106), .B2(n_109), .C1(n_786), .C2(n_790), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_12), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_13), .Y(n_147) );
NAND2xp33_ASAP7_75t_L g576 ( .A(n_14), .B(n_206), .Y(n_576) );
INVx2_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
AOI221x1_ASAP7_75t_L g520 ( .A1(n_16), .A2(n_29), .B1(n_498), .B2(n_500), .C(n_521), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_17), .Y(n_481) );
AND3x1_ASAP7_75t_L g818 ( .A(n_17), .B(n_41), .C(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_18), .B(n_498), .Y(n_572) );
INVx1_ASAP7_75t_L g207 ( .A(n_19), .Y(n_207) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_20), .A2(n_176), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_21), .B(n_171), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_22), .A2(n_81), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_22), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_23), .B(n_209), .Y(n_509) );
AO21x1_ASAP7_75t_L g530 ( .A1(n_24), .A2(n_498), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g485 ( .A(n_25), .Y(n_485) );
INVx1_ASAP7_75t_L g204 ( .A(n_26), .Y(n_204) );
INVx1_ASAP7_75t_SL g191 ( .A(n_27), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_28), .B(n_134), .Y(n_249) );
AOI33xp33_ASAP7_75t_L g229 ( .A1(n_30), .A2(n_55), .A3(n_127), .B1(n_152), .B2(n_230), .B3(n_231), .Y(n_229) );
NAND2x1_ASAP7_75t_L g551 ( .A(n_31), .B(n_209), .Y(n_551) );
NAND2x1_ASAP7_75t_L g583 ( .A(n_32), .B(n_206), .Y(n_583) );
INVx1_ASAP7_75t_L g132 ( .A(n_33), .Y(n_132) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_34), .A2(n_88), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g173 ( .A(n_34), .B(n_88), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_35), .B(n_156), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_36), .B(n_206), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_37), .B(n_209), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_38), .B(n_206), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_39), .A2(n_500), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g140 ( .A(n_40), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g151 ( .A(n_40), .Y(n_151) );
AND2x2_ASAP7_75t_L g160 ( .A(n_40), .B(n_130), .Y(n_160) );
OR2x6_ASAP7_75t_L g483 ( .A(n_41), .B(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_42), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_43), .B(n_498), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_44), .B(n_156), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_45), .A2(n_121), .B1(n_198), .B2(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_46), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_47), .B(n_134), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_48), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_49), .B(n_206), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_50), .B(n_176), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_51), .B(n_134), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_52), .A2(n_500), .B(n_582), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_53), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_54), .B(n_206), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_56), .B(n_134), .Y(n_168) );
INVx1_ASAP7_75t_L g128 ( .A(n_57), .Y(n_128) );
INVx1_ASAP7_75t_L g136 ( .A(n_57), .Y(n_136) );
AND2x2_ASAP7_75t_L g170 ( .A(n_58), .B(n_171), .Y(n_170) );
AOI221xp5_ASAP7_75t_L g177 ( .A1(n_59), .A2(n_76), .B1(n_149), .B2(n_156), .C(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_60), .B(n_156), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_61), .B(n_209), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_62), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_63), .B(n_121), .Y(n_154) );
AOI21xp5_ASAP7_75t_SL g216 ( .A1(n_64), .A2(n_149), .B(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_65), .A2(n_500), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g201 ( .A(n_66), .Y(n_201) );
AO21x1_ASAP7_75t_L g532 ( .A1(n_67), .A2(n_500), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_68), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g167 ( .A(n_69), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_70), .B(n_498), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_71), .A2(n_149), .B(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g545 ( .A(n_72), .B(n_172), .Y(n_545) );
INVx1_ASAP7_75t_L g130 ( .A(n_73), .Y(n_130) );
INVx1_ASAP7_75t_L g138 ( .A(n_73), .Y(n_138) );
AND2x2_ASAP7_75t_L g586 ( .A(n_74), .B(n_120), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_75), .B(n_156), .Y(n_232) );
AND2x2_ASAP7_75t_L g193 ( .A(n_77), .B(n_120), .Y(n_193) );
INVx1_ASAP7_75t_L g202 ( .A(n_78), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_79), .A2(n_149), .B(n_190), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_80), .A2(n_149), .B(n_224), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g807 ( .A(n_81), .Y(n_807) );
INVx1_ASAP7_75t_L g486 ( .A(n_82), .Y(n_486) );
AND2x2_ASAP7_75t_L g495 ( .A(n_83), .B(n_120), .Y(n_495) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_84), .B(n_120), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_85), .B(n_498), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_86), .A2(n_149), .B1(n_227), .B2(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_L g531 ( .A(n_87), .B(n_198), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_89), .B(n_206), .Y(n_510) );
AND2x2_ASAP7_75t_L g554 ( .A(n_90), .B(n_120), .Y(n_554) );
INVx1_ASAP7_75t_L g218 ( .A(n_91), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_92), .B(n_209), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_93), .A2(n_500), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_94), .B(n_206), .Y(n_522) );
AND2x2_ASAP7_75t_L g233 ( .A(n_95), .B(n_120), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_96), .B(n_209), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_97), .A2(n_125), .B(n_131), .C(n_139), .Y(n_124) );
BUFx2_ASAP7_75t_L g801 ( .A(n_98), .Y(n_801) );
INVx1_ASAP7_75t_SL g812 ( .A(n_98), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_99), .A2(n_500), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_100), .B(n_134), .Y(n_219) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_797), .B(n_802), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_792), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_478), .B1(n_487), .B2(n_782), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g786 ( .A1(n_111), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
NAND3x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_357), .C(n_424), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_317), .Y(n_112) );
NOR3x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_268), .C(n_297), .Y(n_113) );
OAI221xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_182), .B1(n_221), .B2(n_236), .C(n_253), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_SL g431 ( .A1(n_115), .A2(n_195), .B(n_432), .C(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_116), .A2(n_403), .B1(n_406), .B2(n_408), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_116), .B(n_222), .Y(n_477) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_161), .Y(n_116) );
BUFx2_ASAP7_75t_L g396 ( .A(n_117), .Y(n_396) );
INVx1_ASAP7_75t_SL g409 ( .A(n_117), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_117), .B(n_264), .Y(n_451) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g234 ( .A(n_118), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g279 ( .A(n_118), .B(n_175), .Y(n_279) );
INVx1_ASAP7_75t_L g290 ( .A(n_118), .Y(n_290) );
INVx2_ASAP7_75t_L g294 ( .A(n_118), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_118), .B(n_265), .Y(n_421) );
OR2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_144), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B1(n_142), .B2(n_143), .Y(n_119) );
INVx3_ASAP7_75t_L g143 ( .A(n_120), .Y(n_143) );
INVx4_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_121), .B(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_122), .Y(n_176) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_123), .B(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g198 ( .A(n_123), .B(n_173), .Y(n_198) );
INVxp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_126), .A2(n_167), .B(n_168), .C(n_169), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g178 ( .A1(n_126), .A2(n_169), .B(n_179), .C(n_180), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_126), .A2(n_169), .B(n_191), .C(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_126), .A2(n_133), .B1(n_201), .B2(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_126), .A2(n_169), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g251 ( .A(n_126), .Y(n_251) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
AND2x2_ASAP7_75t_L g157 ( .A(n_127), .B(n_158), .Y(n_157) );
INVxp33_ASAP7_75t_L g230 ( .A(n_127), .Y(n_230) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g153 ( .A(n_128), .B(n_141), .Y(n_153) );
AND2x4_ASAP7_75t_L g209 ( .A(n_128), .B(n_137), .Y(n_209) );
INVx3_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x6_ASAP7_75t_L g206 ( .A(n_130), .B(n_135), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g498 ( .A(n_134), .B(n_140), .Y(n_498) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx5_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_163), .B(n_170), .Y(n_162) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_143), .A2(n_163), .B(n_170), .Y(n_265) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_143), .A2(n_539), .B(n_545), .Y(n_538) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_143), .A2(n_548), .B(n_554), .Y(n_547) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_143), .A2(n_548), .B(n_554), .Y(n_560) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_143), .A2(n_539), .B(n_545), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B1(n_154), .B2(n_155), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVxp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_153), .Y(n_149) );
NOR2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
AND2x6_ASAP7_75t_L g500 ( .A(n_153), .B(n_160), .Y(n_500) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g244 ( .A(n_157), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_159), .Y(n_245) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g370 ( .A(n_161), .B(n_371), .Y(n_370) );
NOR2x1_ASAP7_75t_L g161 ( .A(n_162), .B(n_174), .Y(n_161) );
INVx2_ASAP7_75t_L g273 ( .A(n_162), .Y(n_273) );
AND2x2_ASAP7_75t_L g293 ( .A(n_162), .B(n_294), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g418 ( .A(n_162), .B(n_294), .Y(n_418) );
AND2x2_ASAP7_75t_L g443 ( .A(n_162), .B(n_286), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_169), .B(n_198), .Y(n_210) );
INVx1_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_169), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_169), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_169), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_169), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_169), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_169), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_169), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_169), .A2(n_575), .B(n_576), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_169), .A2(n_583), .B(n_584), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_171), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_171), .A2(n_497), .B(n_499), .Y(n_496) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_171), .A2(n_520), .B(n_524), .Y(n_519) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_171), .A2(n_520), .B(n_524), .Y(n_590) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
INVx1_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
INVxp67_ASAP7_75t_L g296 ( .A(n_175), .Y(n_296) );
AND2x4_ASAP7_75t_L g336 ( .A(n_175), .B(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_175), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_175), .B(n_287), .Y(n_422) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_181), .Y(n_175) );
INVx2_ASAP7_75t_SL g224 ( .A(n_176), .Y(n_224) );
INVx1_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_194), .Y(n_183) );
AND2x2_ASAP7_75t_L g310 ( .A(n_184), .B(n_282), .Y(n_310) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
AND2x2_ASAP7_75t_L g266 ( .A(n_185), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g277 ( .A(n_185), .Y(n_277) );
INVx1_ASAP7_75t_L g301 ( .A(n_185), .Y(n_301) );
AND2x2_ASAP7_75t_L g304 ( .A(n_185), .B(n_196), .Y(n_304) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_185), .Y(n_326) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_193), .Y(n_185) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_186), .A2(n_580), .B(n_586), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2x1_ASAP7_75t_L g194 ( .A(n_195), .B(n_211), .Y(n_194) );
AND2x2_ASAP7_75t_L g291 ( .A(n_195), .B(n_213), .Y(n_291) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_195), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g427 ( .A(n_195), .Y(n_427) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
AND2x2_ASAP7_75t_L g282 ( .A(n_196), .B(n_241), .Y(n_282) );
NOR2x1_ASAP7_75t_SL g351 ( .A(n_196), .B(n_213), .Y(n_351) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_198), .A2(n_216), .B(n_220), .Y(n_215) );
INVx1_ASAP7_75t_SL g505 ( .A(n_198), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_198), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_198), .A2(n_572), .B(n_573), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_203), .B(n_210), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B1(n_207), .B2(n_208), .Y(n_203) );
INVxp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_211), .B(n_375), .Y(n_388) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g313 ( .A(n_212), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx4_ASAP7_75t_L g252 ( .A(n_213), .Y(n_252) );
AND2x4_ASAP7_75t_L g259 ( .A(n_213), .B(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_213), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_213), .B(n_276), .Y(n_376) );
AND2x2_ASAP7_75t_L g404 ( .A(n_213), .B(n_241), .Y(n_404) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
NAND2x1_ASAP7_75t_SL g221 ( .A(n_222), .B(n_234), .Y(n_221) );
OR2x2_ASAP7_75t_L g432 ( .A(n_222), .B(n_344), .Y(n_432) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g272 ( .A(n_223), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g337 ( .A(n_223), .Y(n_337) );
AND2x2_ASAP7_75t_L g371 ( .A(n_223), .B(n_294), .Y(n_371) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_223) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_226), .B(n_232), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g344 ( .A(n_234), .Y(n_344) );
AND2x2_ASAP7_75t_L g352 ( .A(n_234), .B(n_285), .Y(n_352) );
AND2x2_ASAP7_75t_L g469 ( .A(n_234), .B(n_272), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g423 ( .A(n_238), .B(n_364), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_238), .B(n_263), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_239), .A2(n_300), .B(n_303), .Y(n_299) );
AND2x2_ASAP7_75t_L g369 ( .A(n_239), .B(n_275), .Y(n_369) );
INVx2_ASAP7_75t_SL g456 ( .A(n_239), .Y(n_456) );
AND2x4_ASAP7_75t_SL g239 ( .A(n_240), .B(n_252), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g260 ( .A(n_241), .Y(n_260) );
INVx2_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
AND2x4_ASAP7_75t_L g314 ( .A(n_241), .B(n_267), .Y(n_314) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_247), .Y(n_241) );
NOR3xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .C(n_246), .Y(n_243) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
AND2x4_ASAP7_75t_L g346 ( .A(n_252), .B(n_260), .Y(n_346) );
OR2x2_ASAP7_75t_L g472 ( .A(n_252), .B(n_473), .Y(n_472) );
NAND4xp25_ASAP7_75t_L g253 ( .A(n_254), .B(n_258), .C(n_261), .D(n_266), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g319 ( .A(n_255), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g416 ( .A(n_255), .Y(n_416) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_256), .B(n_264), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_256), .B(n_321), .Y(n_450) );
BUFx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_259), .B(n_275), .Y(n_328) );
INVx2_ASAP7_75t_L g430 ( .A(n_259), .Y(n_430) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_259), .B(n_300), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_259), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g332 ( .A(n_263), .B(n_279), .Y(n_332) );
AND2x2_ASAP7_75t_L g400 ( .A(n_263), .B(n_336), .Y(n_400) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g285 ( .A(n_264), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_265), .Y(n_339) );
AND2x2_ASAP7_75t_L g390 ( .A(n_265), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_265), .B(n_287), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_266), .B(n_430), .Y(n_437) );
INVx1_ASAP7_75t_SL g473 ( .A(n_266), .Y(n_473) );
INVx1_ASAP7_75t_L g302 ( .A(n_267), .Y(n_302) );
AND2x2_ASAP7_75t_L g364 ( .A(n_267), .B(n_307), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_278), .B(n_280), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
AND2x2_ASAP7_75t_L g330 ( .A(n_272), .B(n_279), .Y(n_330) );
AND2x2_ASAP7_75t_L g438 ( .A(n_272), .B(n_289), .Y(n_438) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g312 ( .A(n_275), .Y(n_312) );
AND2x2_ASAP7_75t_L g345 ( .A(n_275), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g350 ( .A(n_275), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_275), .B(n_314), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_275), .B(n_450), .C(n_451), .Y(n_449) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B1(n_291), .B2(n_292), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g375 ( .A(n_282), .Y(n_375) );
AND2x2_ASAP7_75t_L g309 ( .A(n_283), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g331 ( .A(n_283), .B(n_304), .Y(n_331) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_283), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx1_ASAP7_75t_L g342 ( .A(n_285), .Y(n_342) );
AND2x2_ASAP7_75t_L g295 ( .A(n_286), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g384 ( .A(n_290), .B(n_336), .Y(n_384) );
INVx1_ASAP7_75t_L g442 ( .A(n_290), .Y(n_442) );
INVx1_ASAP7_75t_L g298 ( .A(n_292), .Y(n_298) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_293), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g429 ( .A(n_293), .B(n_336), .Y(n_429) );
AND2x2_ASAP7_75t_L g395 ( .A(n_295), .B(n_396), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_295), .B(n_464), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_308), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_300), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g356 ( .A(n_300), .B(n_305), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_300), .B(n_346), .Y(n_407) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_301), .B(n_364), .Y(n_394) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_301), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_303), .A2(n_330), .B1(n_331), .B2(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_304), .B(n_346), .Y(n_365) );
INVx1_ASAP7_75t_L g466 ( .A(n_304), .Y(n_466) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B(n_315), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_310), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g447 ( .A(n_313), .Y(n_447) );
INVx4_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
INVxp33_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g377 ( .A(n_316), .B(n_378), .Y(n_377) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_318), .B(n_333), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_329), .Y(n_318) );
INVx1_ASAP7_75t_L g367 ( .A(n_320), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
INVx1_ASAP7_75t_L g405 ( .A(n_325), .Y(n_405) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_330), .A2(n_369), .B1(n_370), .B2(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
NAND4xp25_ASAP7_75t_SL g333 ( .A(n_334), .B(n_340), .C(n_347), .D(n_353), .Y(n_333) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g355 ( .A(n_336), .Y(n_355) );
AND2x2_ASAP7_75t_L g467 ( .A(n_336), .B(n_464), .Y(n_467) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g474 ( .A(n_344), .B(n_411), .Y(n_474) );
INVx1_ASAP7_75t_L g471 ( .A(n_345), .Y(n_471) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_346), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B(n_352), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_385), .Y(n_357) );
NOR3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_373), .C(n_381), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_366), .B(n_368), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_363), .A2(n_395), .B1(n_398), .B2(n_400), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_366), .A2(n_374), .B1(n_377), .B2(n_379), .Y(n_373) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g378 ( .A(n_371), .Y(n_378) );
AND2x4_ASAP7_75t_L g389 ( .A(n_371), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_376), .Y(n_476) );
AOI31xp33_ASAP7_75t_L g475 ( .A1(n_379), .A2(n_452), .A3(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_401), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_387), .B(n_397), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_392), .B2(n_395), .Y(n_387) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_399), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_402), .B(n_412), .Y(n_401) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g413 ( .A(n_404), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_404), .A2(n_462), .B1(n_465), .B2(n_467), .Y(n_461) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_409), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_419), .B2(n_423), .Y(n_412) );
NOR2xp33_ASAP7_75t_SL g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_SL g464 ( .A(n_421), .Y(n_464) );
INVx2_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_459), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_431), .B(n_434), .C(n_448), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_430), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_435), .B(n_439), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_444), .B2(n_446), .Y(n_439) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AND2x2_ASAP7_75t_L g444 ( .A(n_442), .B(n_445), .Y(n_444) );
AO22x1_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B1(n_453), .B2(n_457), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_470), .C(n_475), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_461), .B(n_468), .Y(n_460) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI21xp33_ASAP7_75t_R g470 ( .A1(n_471), .A2(n_472), .B(n_474), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_479), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
OR2x6_ASAP7_75t_SL g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x6_ASAP7_75t_SL g785 ( .A(n_481), .B(n_483), .Y(n_785) );
OR2x2_ASAP7_75t_L g791 ( .A(n_481), .B(n_483), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_481), .B(n_482), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g817 ( .A(n_484), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_SL g788 ( .A(n_488), .Y(n_788) );
NOR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_669), .Y(n_488) );
AO211x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_514), .B(n_564), .C(n_637), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AND3x2_ASAP7_75t_L g718 ( .A(n_492), .B(n_599), .C(n_615), .Y(n_718) );
AND2x4_ASAP7_75t_L g721 ( .A(n_492), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_504), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g577 ( .A(n_493), .B(n_578), .Y(n_577) );
INVx4_ASAP7_75t_L g630 ( .A(n_493), .Y(n_630) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_493), .B(n_624), .Y(n_715) );
AND2x2_ASAP7_75t_L g758 ( .A(n_493), .B(n_579), .Y(n_758) );
INVx5_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g607 ( .A(n_494), .Y(n_607) );
AND2x2_ASAP7_75t_L g626 ( .A(n_494), .B(n_570), .Y(n_626) );
AND2x2_ASAP7_75t_L g644 ( .A(n_494), .B(n_579), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_494), .B(n_578), .Y(n_704) );
NOR2x1_ASAP7_75t_SL g731 ( .A(n_494), .B(n_504), .Y(n_731) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_504), .B(n_570), .Y(n_569) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_505), .B(n_513), .Y(n_512) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
AO21x1_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_546), .B(n_555), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_516), .A2(n_613), .B1(n_617), .B2(n_618), .Y(n_612) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
AND2x2_ASAP7_75t_L g673 ( .A(n_517), .B(n_561), .Y(n_673) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g606 ( .A(n_518), .B(n_589), .Y(n_606) );
AND2x2_ASAP7_75t_L g678 ( .A(n_518), .B(n_563), .Y(n_678) );
AND2x2_ASAP7_75t_L g697 ( .A(n_518), .B(n_663), .Y(n_697) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g556 ( .A(n_519), .Y(n_556) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_519), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_525), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g657 ( .A(n_526), .B(n_558), .Y(n_657) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
AND2x2_ASAP7_75t_L g561 ( .A(n_527), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g594 ( .A(n_527), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_527), .B(n_590), .Y(n_654) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g747 ( .A(n_528), .Y(n_747) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g589 ( .A(n_529), .Y(n_589) );
OAI21x1_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_532), .B(n_536), .Y(n_529) );
INVx1_ASAP7_75t_L g537 ( .A(n_531), .Y(n_537) );
INVx2_ASAP7_75t_L g595 ( .A(n_538), .Y(n_595) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_538), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_544), .Y(n_539) );
INVx2_ASAP7_75t_L g591 ( .A(n_546), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_546), .B(n_723), .Y(n_749) );
AND2x2_ASAP7_75t_L g768 ( .A(n_546), .B(n_758), .Y(n_768) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_SL g636 ( .A(n_547), .B(n_595), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g635 ( .A(n_556), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_556), .B(n_605), .Y(n_640) );
INVx1_ASAP7_75t_SL g767 ( .A(n_556), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_557), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g593 ( .A(n_558), .Y(n_593) );
AND2x2_ASAP7_75t_L g779 ( .A(n_558), .B(n_780), .Y(n_779) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g655 ( .A(n_559), .B(n_562), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_559), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g709 ( .A(n_559), .B(n_563), .Y(n_709) );
AND2x2_ASAP7_75t_L g740 ( .A(n_559), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g605 ( .A(n_560), .B(n_563), .Y(n_605) );
INVxp67_ASAP7_75t_L g622 ( .A(n_560), .Y(n_622) );
BUFx3_ASAP7_75t_L g663 ( .A(n_560), .Y(n_663) );
AND2x2_ASAP7_75t_L g683 ( .A(n_561), .B(n_684), .Y(n_683) );
NAND2xp33_ASAP7_75t_L g696 ( .A(n_561), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_562), .B(n_589), .Y(n_652) );
AND2x2_ASAP7_75t_L g741 ( .A(n_562), .B(n_590), .Y(n_741) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g668 ( .A(n_563), .B(n_590), .Y(n_668) );
OR3x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_612), .C(n_627), .Y(n_564) );
OAI321xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_577), .A3(n_587), .B1(n_592), .B2(n_596), .C(n_604), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_569), .Y(n_643) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_569), .Y(n_661) );
OR2x2_ASAP7_75t_L g665 ( .A(n_569), .B(n_577), .Y(n_665) );
BUFx3_ASAP7_75t_L g599 ( .A(n_570), .Y(n_599) );
AND2x2_ASAP7_75t_L g616 ( .A(n_570), .B(n_602), .Y(n_616) );
INVx1_ASAP7_75t_L g633 ( .A(n_570), .Y(n_633) );
INVx2_ASAP7_75t_L g649 ( .A(n_570), .Y(n_649) );
OR2x2_ASAP7_75t_L g688 ( .A(n_570), .B(n_578), .Y(n_688) );
INVx2_ASAP7_75t_L g676 ( .A(n_577), .Y(n_676) );
AND2x2_ASAP7_75t_L g600 ( .A(n_578), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g615 ( .A(n_578), .Y(n_615) );
AND2x4_ASAP7_75t_L g624 ( .A(n_578), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_578), .B(n_601), .Y(n_647) );
AND2x2_ASAP7_75t_L g754 ( .A(n_578), .B(n_649), .Y(n_754) );
INVx4_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_579), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_585), .Y(n_580) );
INVx1_ASAP7_75t_L g641 ( .A(n_587), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_588), .B(n_591), .Y(n_587) );
AND2x2_ASAP7_75t_L g728 ( .A(n_588), .B(n_655), .Y(n_728) );
INVx1_ASAP7_75t_SL g745 ( .A(n_588), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_588), .B(n_721), .Y(n_774) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OR2x2_ASAP7_75t_L g617 ( .A(n_589), .B(n_590), .Y(n_617) );
AND2x2_ASAP7_75t_L g710 ( .A(n_591), .B(n_606), .Y(n_710) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_595), .B(n_606), .Y(n_733) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_597), .A2(n_746), .B1(n_751), .B2(n_753), .Y(n_750) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g675 ( .A(n_598), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g770 ( .A(n_598), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g726 ( .A(n_599), .B(n_644), .Y(n_726) );
AND2x4_ASAP7_75t_L g680 ( .A(n_600), .B(n_626), .Y(n_680) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_602), .Y(n_778) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g611 ( .A(n_603), .Y(n_611) );
INVx1_ASAP7_75t_L g625 ( .A(n_603), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .C(n_607), .D(n_608), .Y(n_604) );
AND2x2_ASAP7_75t_L g762 ( .A(n_605), .B(n_747), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_605), .B(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_606), .B(n_682), .Y(n_681) );
OAI322xp33_ASAP7_75t_L g689 ( .A1(n_606), .A2(n_690), .A3(n_694), .B1(n_696), .B2(n_698), .C1(n_700), .C2(n_705), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_606), .B(n_655), .Y(n_705) );
INVx1_ASAP7_75t_L g773 ( .A(n_606), .Y(n_773) );
INVx2_ASAP7_75t_L g619 ( .A(n_607), .Y(n_619) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_610), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_611), .B(n_630), .Y(n_687) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_614), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g660 ( .A(n_615), .Y(n_660) );
AND2x2_ASAP7_75t_L g732 ( .A(n_615), .B(n_643), .Y(n_732) );
AOI31xp33_ASAP7_75t_L g618 ( .A1(n_616), .A2(n_619), .A3(n_620), .B(n_623), .Y(n_618) );
AND2x2_ASAP7_75t_L g629 ( .A(n_616), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g757 ( .A(n_616), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_SL g764 ( .A(n_616), .B(n_644), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_616), .Y(n_765) );
INVx1_ASAP7_75t_SL g723 ( .A(n_617), .Y(n_723) );
NAND3xp33_ASAP7_75t_SL g751 ( .A(n_617), .B(n_745), .C(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g651 ( .A(n_622), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_624), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g693 ( .A(n_624), .Y(n_693) );
AOI322xp5_ASAP7_75t_L g775 ( .A1(n_624), .A2(n_654), .A3(n_657), .B1(n_776), .B2(n_777), .C1(n_779), .C2(n_781), .Y(n_775) );
AND2x2_ASAP7_75t_L g781 ( .A(n_624), .B(n_630), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .B(n_634), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_630), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g776 ( .A(n_630), .B(n_663), .Y(n_776) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g702 ( .A(n_633), .Y(n_702) );
AND2x2_ASAP7_75t_L g730 ( .A(n_633), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g777 ( .A(n_633), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g682 ( .A(n_636), .Y(n_682) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
O2A1O1Ixp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B(n_642), .C(n_645), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g699 ( .A(n_644), .B(n_649), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B(n_656), .C(n_658), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_646), .A2(n_672), .B1(n_674), .B2(n_677), .C(n_679), .Y(n_671) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g691 ( .A(n_648), .Y(n_691) );
OR2x2_ASAP7_75t_L g711 ( .A(n_648), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g756 ( .A(n_651), .Y(n_756) );
INVx1_ASAP7_75t_L g780 ( .A(n_652), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_655), .Y(n_653) );
AND2x2_ASAP7_75t_L g662 ( .A(n_654), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_654), .B(n_724), .Y(n_736) );
INVx1_ASAP7_75t_L g716 ( .A(n_655), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B1(n_664), .B2(n_666), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_SL g724 ( .A(n_663), .Y(n_724) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND4xp75_ASAP7_75t_L g669 ( .A(n_670), .B(n_706), .C(n_734), .D(n_759), .Y(n_669) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_671), .B(n_689), .Y(n_670) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_SL g746 ( .A(n_678), .B(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B1(n_683), .B2(n_685), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_682), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx2_ASAP7_75t_L g722 ( .A(n_688), .Y(n_722) );
OR2x2_ASAP7_75t_L g737 ( .A(n_688), .B(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g752 ( .A(n_697), .Y(n_752) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
OAI21xp5_ASAP7_75t_SL g743 ( .A1(n_699), .A2(n_744), .B(n_746), .Y(n_743) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_719), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B1(n_714), .B2(n_716), .C(n_717), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g755 ( .A1(n_709), .A2(n_756), .B(n_757), .Y(n_755) );
INVx3_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
OAI322xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .A3(n_724), .B1(n_725), .B2(n_727), .C1(n_729), .C2(n_733), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g742 ( .A(n_730), .Y(n_742) );
INVx1_ASAP7_75t_L g738 ( .A(n_731), .Y(n_738) );
AND2x2_ASAP7_75t_L g753 ( .A(n_731), .B(n_754), .Y(n_753) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_748), .Y(n_734) );
OAI221xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_739), .B2(n_742), .C(n_743), .Y(n_735) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
OAI211xp5_ASAP7_75t_SL g748 ( .A1(n_742), .A2(n_749), .B(n_750), .C(n_755), .Y(n_748) );
INVx2_ASAP7_75t_SL g771 ( .A(n_758), .Y(n_771) );
NOR2x1_ASAP7_75t_L g759 ( .A(n_760), .B(n_769), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B1(n_765), .B2(n_766), .Y(n_760) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
OAI211xp5_ASAP7_75t_SL g769 ( .A1(n_770), .A2(n_772), .B(n_774), .C(n_775), .Y(n_769) );
CKINVDCx11_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
INVx3_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g789 ( .A(n_785), .Y(n_789) );
XOR2x2_ASAP7_75t_L g804 ( .A(n_788), .B(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_793), .A2(n_804), .B(n_808), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_R g810 ( .A(n_796), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
BUFx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_811), .Y(n_802) );
INVx1_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
BUFx4f_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_SL g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
endmodule