module real_jpeg_30206_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_29),
.B1(n_34),
.B2(n_52),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_71),
.B1(n_72),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_1),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_1),
.A2(n_29),
.B1(n_34),
.B2(n_80),
.Y(n_186)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_27),
.B(n_103),
.Y(n_160)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_71),
.B1(n_72),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_4),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_4),
.A2(n_75),
.B1(n_76),
.B2(n_112),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_112),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_4),
.A2(n_29),
.B1(n_34),
.B2(n_112),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_29),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_6),
.A2(n_39),
.B1(n_75),
.B2(n_76),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_123)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_8),
.A2(n_11),
.B(n_29),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_29),
.B1(n_34),
.B2(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_35),
.B1(n_75),
.B2(n_76),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_11),
.B(n_76),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_76),
.B(n_144),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_100),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_11),
.B(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_199),
.Y(n_202)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_13),
.A2(n_75),
.B1(n_76),
.B2(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_71),
.B1(n_72),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_15),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_78),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_15),
.A2(n_29),
.B1(n_34),
.B2(n_78),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_95),
.B2(n_113),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_53),
.B2(n_54),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_28),
.A2(n_57),
.B(n_58),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_28),
.A2(n_32),
.B1(n_57),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_28),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_36),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_28),
.A2(n_191),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_32),
.B(n_100),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_34),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_37),
.A2(n_141),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_38),
.A2(n_59),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_41),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_41),
.A2(n_48),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_41),
.A2(n_153),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_41),
.A2(n_48),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_41),
.A2(n_48),
.B1(n_152),
.B2(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_44),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_43),
.A2(n_75),
.A3(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_44),
.B(n_89),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_44),
.A2(n_47),
.B(n_100),
.C(n_177),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_49),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_48),
.B(n_100),
.Y(n_197)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_60),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_63),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_82),
.B2(n_83),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_77),
.B1(n_81),
.B2(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_74),
.B1(n_99),
.B2(n_111),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_71),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_100),
.CON(n_99),
.SN(n_99)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_75),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_100),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_91),
.B(n_93),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_88),
.B1(n_106),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_85),
.A2(n_88),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_88),
.B1(n_128),
.B2(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.C(n_108),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_97),
.B(n_101),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_115),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_118),
.B(n_119),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_129),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_125),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_129),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_232),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_228),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_215),
.B(n_227),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_168),
.B(n_214),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_154),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_137),
.B(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.C(n_150),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_138),
.A2(n_139),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_163),
.B2(n_164),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_165),
.C(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_157),
.B(n_159),
.C(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_208),
.B(n_213),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_187),
.B(n_207),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_171),
.B(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_176),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_184),
.C(n_185),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_195),
.B(n_206),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_193),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_201),
.B(n_205),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_217)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);


endmodule