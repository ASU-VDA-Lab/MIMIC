module fake_jpeg_28804_n_430 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_430);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_430;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_62),
.Y(n_99)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_55),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_19),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_82),
.Y(n_130)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_84),
.Y(n_109)
);

BUFx2_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_16),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_88),
.B(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_125),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_39),
.B1(n_66),
.B2(n_53),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_70),
.B(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_39),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_43),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_75),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_64),
.A2(n_28),
.B(n_19),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_86),
.C(n_50),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_136),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_28),
.B1(n_37),
.B2(n_47),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_150),
.B1(n_167),
.B2(n_129),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_58),
.B1(n_83),
.B2(n_68),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_135),
.A2(n_149),
.B1(n_108),
.B2(n_48),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_122),
.Y(n_136)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_139),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_145),
.C(n_97),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_76),
.C(n_73),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_156),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_71),
.B1(n_67),
.B2(n_49),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_46),
.B1(n_21),
.B2(n_33),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_96),
.B1(n_97),
.B2(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_39),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_92),
.A2(n_54),
.A3(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_109),
.B(n_54),
.C(n_27),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_164),
.Y(n_193)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_95),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_90),
.B(n_19),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_27),
.Y(n_195)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

AOI22x1_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_86),
.B1(n_107),
.B2(n_102),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_168),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_179),
.B1(n_180),
.B2(n_149),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_176),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_195),
.B(n_154),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_182),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_119),
.B1(n_87),
.B2(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_15),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_132),
.A2(n_108),
.B1(n_123),
.B2(n_113),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_191),
.B1(n_138),
.B2(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_219),
.B1(n_175),
.B2(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_138),
.B(n_145),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_205),
.B(n_173),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_133),
.B(n_140),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_147),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_214),
.B1(n_215),
.B2(n_196),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_137),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_165),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_157),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_120),
.B1(n_87),
.B2(n_119),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_120),
.B1(n_143),
.B2(n_144),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_167),
.B1(n_161),
.B2(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_188),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_231),
.B1(n_234),
.B2(n_239),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_227),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_186),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_186),
.B1(n_185),
.B2(n_191),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_188),
.B1(n_173),
.B2(n_189),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_178),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_196),
.B1(n_184),
.B2(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_200),
.B1(n_198),
.B2(n_207),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_193),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_171),
.C(n_121),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_215),
.B(n_201),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_136),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_213),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_SL g285 ( 
.A1(n_245),
.A2(n_237),
.A3(n_224),
.B1(n_103),
.B2(n_101),
.C1(n_129),
.C2(n_139),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_210),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_246),
.Y(n_273)
);

AO22x1_ASAP7_75t_SL g247 ( 
.A1(n_241),
.A2(n_211),
.B1(n_214),
.B2(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_23),
.Y(n_287)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_258),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_268),
.B1(n_222),
.B2(n_231),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_216),
.B(n_182),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_233),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_264),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_101),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_233),
.C(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_187),
.C(n_192),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_202),
.B1(n_217),
.B2(n_170),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_183),
.B1(n_148),
.B2(n_102),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_171),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_267),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_230),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_183),
.B1(n_196),
.B2(n_187),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_271),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_248),
.A2(n_232),
.B1(n_227),
.B2(n_241),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_292),
.B1(n_294),
.B2(n_253),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_298),
.B1(n_271),
.B2(n_258),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_246),
.A2(n_242),
.B(n_232),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_276),
.B(n_282),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_236),
.B(n_228),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_278),
.A2(n_265),
.B1(n_260),
.B2(n_247),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_286),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_270),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_114),
.C(n_38),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_293),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_187),
.B1(n_192),
.B2(n_121),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_255),
.B(n_152),
.CI(n_155),
.CON(n_293),
.SN(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_164),
.B1(n_162),
.B2(n_159),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_95),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_94),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_259),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_248),
.A2(n_94),
.B(n_163),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_262),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_277),
.A2(n_244),
.B1(n_247),
.B2(n_270),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_305),
.B1(n_308),
.B2(n_316),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_298),
.B1(n_282),
.B2(n_299),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_268),
.B1(n_244),
.B2(n_250),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_303),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_283),
.B(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_273),
.A2(n_261),
.B1(n_257),
.B2(n_249),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_295),
.B1(n_289),
.B2(n_272),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_257),
.B1(n_245),
.B2(n_252),
.Y(n_310)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_312),
.Y(n_337)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_324),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_274),
.A2(n_33),
.B1(n_21),
.B2(n_38),
.Y(n_318)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_123),
.B1(n_113),
.B2(n_38),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_320),
.A2(n_297),
.B1(n_280),
.B2(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_288),
.C(n_291),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_114),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_275),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_27),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_290),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_328),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_322),
.C(n_317),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_284),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_311),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_338),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_31),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_304),
.A2(n_312),
.B(n_307),
.C(n_300),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_333),
.A2(n_314),
.B1(n_23),
.B2(n_34),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_345),
.B1(n_36),
.B2(n_31),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

NOR2x1_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_320),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_293),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_36),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_292),
.B(n_278),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_346),
.A2(n_302),
.B(n_324),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_294),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_323),
.Y(n_353)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_316),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_350),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_349),
.B(n_363),
.Y(n_379)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_364),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_354),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_314),
.C(n_38),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_357),
.C(n_362),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_36),
.C(n_33),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_34),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_359),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_36),
.C(n_33),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_332),
.C(n_331),
.Y(n_363)
);

XOR2x1_ASAP7_75t_SL g364 ( 
.A(n_333),
.B(n_15),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_365),
.A2(n_340),
.B1(n_339),
.B2(n_344),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_366),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_375),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_364),
.A2(n_341),
.B(n_336),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_372),
.A2(n_358),
.B(n_345),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_360),
.A2(n_333),
.B1(n_325),
.B2(n_346),
.Y(n_374)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_356),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_380),
.Y(n_389)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_343),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_382),
.Y(n_390)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_379),
.B(n_348),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_SL g386 ( 
.A1(n_378),
.A2(n_333),
.B(n_354),
.C(n_365),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_388),
.B(n_392),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_391),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_371),
.A2(n_363),
.B(n_349),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_357),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_368),
.B(n_359),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_355),
.C(n_362),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_24),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_372),
.B(n_353),
.Y(n_394)
);

AOI21xp33_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_24),
.B(n_1),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_371),
.C(n_369),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_29),
.C(n_25),
.Y(n_410)
);

NOR3xp33_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_370),
.C(n_377),
.Y(n_396)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_382),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_399),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_384),
.A2(n_373),
.B1(n_377),
.B2(n_331),
.Y(n_399)
);

OAI21x1_ASAP7_75t_SL g400 ( 
.A1(n_394),
.A2(n_373),
.B(n_14),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_403),
.B(n_0),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_392),
.A2(n_14),
.B1(n_24),
.B2(n_23),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_401),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_3),
.C(n_4),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_410),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_402),
.A2(n_404),
.B(n_398),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_407),
.A2(n_413),
.B(n_414),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_412),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_25),
.C(n_2),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_413)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_408),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_416),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_3),
.B(n_5),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_419),
.B(n_5),
.Y(n_422)
);

OAI31xp33_ASAP7_75t_SL g420 ( 
.A1(n_412),
.A2(n_3),
.A3(n_5),
.B(n_6),
.Y(n_420)
);

AOI322xp5_ASAP7_75t_L g421 ( 
.A1(n_420),
.A2(n_25),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_SL g425 ( 
.A1(n_421),
.A2(n_422),
.B(n_418),
.C(n_415),
.Y(n_425)
);

AOI322xp5_ASAP7_75t_L g423 ( 
.A1(n_417),
.A2(n_410),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_7),
.Y(n_423)
);

AOI21xp33_ASAP7_75t_L g426 ( 
.A1(n_423),
.A2(n_424),
.B(n_8),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_425),
.B(n_426),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_7),
.Y(n_428)
);

AOI31xp67_ASAP7_75t_L g429 ( 
.A1(n_428),
.A2(n_7),
.A3(n_8),
.B(n_11),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_11),
.C(n_12),
.Y(n_430)
);


endmodule