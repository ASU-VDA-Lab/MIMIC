module real_jpeg_24793_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_215;
wire n_166;
wire n_221;
wire n_292;
wire n_176;
wire n_249;
wire n_286;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_167;
wire n_295;
wire n_128;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_1),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_25),
.B1(n_54),
.B2(n_56),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_25),
.B1(n_74),
.B2(n_75),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_5),
.A2(n_15),
.B(n_302),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_5),
.B(n_303),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_22),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_7),
.A2(n_35),
.B1(n_54),
.B2(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_35),
.B1(n_74),
.B2(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_61),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_54),
.B1(n_56),
.B2(n_61),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_61),
.B1(n_74),
.B2(n_75),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_44),
.B1(n_54),
.B2(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_44),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_10),
.A2(n_44),
.B1(n_74),
.B2(n_75),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_29),
.C(n_33),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_30),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_10),
.B(n_51),
.C(n_54),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_10),
.B(n_71),
.C(n_74),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_10),
.B(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_10),
.B(n_103),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_10),
.B(n_64),
.Y(n_252)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_295),
.B(n_299),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_77),
.B(n_294),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_18),
.B(n_37),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_18),
.B(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_18),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_40),
.B(n_41),
.Y(n_39)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_22),
.B(n_189),
.Y(n_188)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_26),
.A2(n_30),
.B1(n_42),
.B2(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_33),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_33),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_34),
.B(n_298),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_38),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_38),
.B(n_292),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_45),
.CI(n_57),
.CON(n_38),
.SN(n_38)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_40),
.A2(n_41),
.B(n_60),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_48),
.A2(n_53),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_49),
.A2(n_64),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_49),
.B(n_108),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_53),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_53),
.A2(n_107),
.B(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_56),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_54),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_65),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_58),
.B(n_126),
.C(n_134),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_58),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_134),
.B1(n_135),
.B2(n_148),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_58),
.A2(n_105),
.B1(n_148),
.B2(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_58),
.B(n_105),
.C(n_186),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_62),
.A2(n_65),
.B1(n_115),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_62),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_63),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_65),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_111),
.C(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_76),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_67),
.B(n_93),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_69),
.A2(n_93),
.B1(n_103),
.B2(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_73),
.A2(n_92),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_74),
.B(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_291),
.B(n_293),
.Y(n_77)
);

OAI211xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_136),
.B(n_150),
.C(n_290),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_120),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_120),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_98),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_100),
.C(n_109),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_89),
.B(n_94),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_94),
.B1(n_95),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_82),
.A2(n_90),
.B1(n_123),
.B2(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_84),
.B(n_196),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_88),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_85),
.B(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_87),
.A2(n_128),
.B(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_87),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_96),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_109),
.B2(n_110),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_101),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_105),
.B(n_208),
.C(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_105),
.A2(n_198),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_112),
.B1(n_144),
.B2(n_149),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_134),
.C(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_111),
.A2(n_112),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_111),
.A2(n_112),
.B1(n_168),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_160),
.C(n_168),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_112),
.B(n_140),
.C(n_144),
.Y(n_292)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_124),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_127),
.Y(n_281)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_131),
.A2(n_132),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_131),
.A2(n_132),
.B1(n_221),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_132),
.B(n_215),
.C(n_221),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_191),
.C(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_134),
.A2(n_135),
.B1(n_182),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_134),
.A2(n_135),
.B1(n_166),
.B2(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_135),
.B(n_166),
.C(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_151),
.C(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_138),
.B(n_139),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_172),
.B(n_289),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_170),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_154),
.B(n_170),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_155),
.B(n_157),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_159),
.B(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_160),
.A2(n_161),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_166),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_193),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_166),
.A2(n_179),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_166),
.B(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_168),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_284),
.B(n_288),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_211),
.B(n_270),
.C(n_283),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_200),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_175),
.B(n_200),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_185),
.B2(n_199),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_178),
.B(n_184),
.C(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_190),
.A2(n_191),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_244),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_191)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_202),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_209),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_269),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_230),
.B(n_268),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_227),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_214),
.B(n_227),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_215),
.A2(n_216),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_261),
.B(n_267),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_255),
.B(n_260),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_247),
.B(n_254),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_246),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_243),
.B(n_245),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_279),
.B2(n_280),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_280),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);


endmodule