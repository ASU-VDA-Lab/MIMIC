module fake_jpeg_28946_n_27 (n_3, n_2, n_1, n_0, n_4, n_5, n_27);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_27;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

OA22x2_ASAP7_75t_L g6 ( 
.A1(n_0),
.A2(n_3),
.B1(n_2),
.B2(n_4),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_0),
.A2(n_3),
.B1(n_2),
.B2(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_8),
.B(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_14),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_6),
.A2(n_1),
.B(n_10),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_13),
.A2(n_16),
.B(n_6),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_6),
.A2(n_7),
.B(n_9),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_10),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_8),
.CI(n_6),
.CON(n_18),
.SN(n_18)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_7),
.C(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

AO221x1_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.C(n_9),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.C(n_18),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_19),
.B(n_18),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_22),
.Y(n_27)
);


endmodule