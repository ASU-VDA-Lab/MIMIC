module fake_ariane_967_n_1669 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1669);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1669;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_48),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_21),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_113),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_69),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_45),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_77),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_41),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_100),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_90),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_68),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_88),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_142),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_42),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_103),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_57),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_22),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_22),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_46),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_0),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_32),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_134),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_43),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_86),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_95),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_16),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_139),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_9),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_25),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_70),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_67),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_129),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_53),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_33),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_66),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_48),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_1),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_11),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_106),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_96),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_118),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_80),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_9),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_120),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_24),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_5),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_75),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_62),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_99),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_25),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_16),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_30),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_47),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_131),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_19),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_132),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_7),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_46),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_28),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_1),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_65),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_21),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_3),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_23),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_152),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_5),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_43),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_108),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_64),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_23),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_127),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_18),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_11),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_63),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_112),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_12),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_24),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_38),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_19),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_42),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_18),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_151),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_135),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_83),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_17),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_73),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_12),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_84),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_10),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_34),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_29),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_52),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_15),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_30),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_3),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_155),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_153),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_109),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_93),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_122),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_119),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_49),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_140),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_117),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_125),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_31),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_190),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_193),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_218),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_254),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_2),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_233),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_156),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_210),
.B(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_267),
.Y(n_328)
);

NOR2x1_ASAP7_75t_L g329 ( 
.A(n_165),
.B(n_180),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_189),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_187),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_195),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_163),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_187),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_254),
.B(n_6),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_173),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_187),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_187),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_196),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_197),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_215),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_199),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_164),
.B(n_6),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_221),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_199),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_276),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_199),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_172),
.B(n_7),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_225),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_235),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_236),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_199),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_239),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_175),
.B(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_216),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_216),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_310),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_216),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_159),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_173),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_241),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_216),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_160),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_208),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_243),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_253),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_246),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_253),
.Y(n_374)
);

BUFx6f_ASAP7_75t_SL g375 ( 
.A(n_158),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_247),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_210),
.B(n_265),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_178),
.B(n_8),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_249),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_213),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_253),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_158),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_165),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_380),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_322),
.B(n_178),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_380),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_380),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_182),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_370),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_382),
.A2(n_198),
.B1(n_280),
.B2(n_211),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_184),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_318),
.B(n_158),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_317),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_324),
.B(n_307),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_329),
.B(n_253),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_361),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_200),
.Y(n_419)
);

BUFx8_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_356),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_332),
.B(n_203),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_321),
.B(n_180),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_382),
.B(n_171),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_339),
.B(n_207),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_324),
.B(n_307),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_307),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_377),
.B(n_319),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_374),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_345),
.B(n_202),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_341),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_343),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_433),
.A2(n_351),
.B1(n_358),
.B2(n_375),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_370),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_395),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_439),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_420),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_433),
.A2(n_375),
.B1(n_316),
.B2(n_312),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_323),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_414),
.B(n_171),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_371),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_371),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_364),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_352),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_274),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_336),
.B1(n_240),
.B2(n_174),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_396),
.B(n_353),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_392),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_354),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_369),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_417),
.A2(n_427),
.B1(n_408),
.B2(n_402),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_417),
.A2(n_161),
.B1(n_230),
.B2(n_228),
.Y(n_482)
);

BUFx6f_ASAP7_75t_SL g483 ( 
.A(n_427),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_392),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_408),
.B(n_357),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_396),
.B(n_366),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_408),
.A2(n_379),
.B1(n_376),
.B2(n_373),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_400),
.B(n_209),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_427),
.B(n_400),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_405),
.B(n_214),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_441),
.B(n_328),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_431),
.B(n_266),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_441),
.B(n_378),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_398),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_441),
.B(n_223),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_403),
.B(n_255),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_427),
.A2(n_257),
.B1(n_256),
.B2(n_251),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_420),
.B(n_274),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_417),
.A2(n_226),
.B1(n_168),
.B2(n_306),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_410),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_410),
.B(n_224),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_404),
.B(n_234),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_392),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_420),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_402),
.A2(n_288),
.B1(n_290),
.B2(n_287),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_401),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_401),
.Y(n_527)
);

AND3x2_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_222),
.C(n_188),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_411),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_390),
.B(n_237),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_427),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_404),
.B(n_244),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_227),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_427),
.B(n_341),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_432),
.B(n_248),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_415),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_392),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_390),
.B(n_268),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_432),
.B(n_277),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_409),
.A2(n_296),
.B1(n_282),
.B2(n_303),
.Y(n_547)
);

NOR2x1p5_ASAP7_75t_L g548 ( 
.A(n_395),
.B(n_281),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_415),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_392),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_409),
.B(n_348),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_403),
.A2(n_297),
.B1(n_298),
.B2(n_294),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_415),
.B(n_418),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_436),
.A2(n_297),
.B1(n_298),
.B2(n_294),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_420),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_386),
.A2(n_275),
.B1(n_289),
.B2(n_301),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_436),
.B(n_447),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_446),
.B(n_308),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_407),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_415),
.B(n_348),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_407),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_436),
.B(n_447),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_420),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_407),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_447),
.A2(n_293),
.B1(n_281),
.B2(n_287),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_407),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_407),
.B(n_157),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_407),
.B(n_157),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_406),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_406),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_384),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_416),
.B(n_291),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_446),
.B(n_291),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_426),
.B(n_288),
.C(n_290),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_418),
.B(n_355),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_418),
.B(n_355),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_416),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_384),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_407),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_426),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_416),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_407),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_407),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_413),
.B(n_292),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_425),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_419),
.B(n_424),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_419),
.B(n_359),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_R g592 ( 
.A(n_386),
.B(n_334),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_428),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_386),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_503),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_453),
.B(n_424),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_479),
.B(n_386),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_557),
.A2(n_437),
.B1(n_444),
.B2(n_428),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_453),
.B(n_162),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_517),
.B(n_342),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_557),
.A2(n_460),
.B1(n_481),
.B2(n_470),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_590),
.B(n_437),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_428),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_429),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_491),
.B(n_162),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_429),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_450),
.B(n_347),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_458),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_463),
.A2(n_293),
.B1(n_292),
.B2(n_269),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_460),
.B(n_429),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_468),
.B(n_464),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_467),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_467),
.B(n_430),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_461),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_349),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_461),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_536),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_475),
.A2(n_383),
.B(n_387),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_460),
.B(n_430),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_522),
.A2(n_383),
.B(n_387),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_508),
.B(n_362),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_542),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_460),
.B(n_532),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_555),
.A2(n_270),
.B1(n_263),
.B2(n_264),
.C(n_273),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_460),
.B(n_430),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_452),
.B(n_166),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_465),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_544),
.B(n_435),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_588),
.B(n_278),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_493),
.B(n_279),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_584),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_452),
.B(n_485),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_470),
.B(n_435),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_474),
.B(n_166),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_452),
.B(n_167),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_470),
.B(n_435),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_456),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_470),
.B(n_444),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_496),
.A2(n_229),
.B1(n_169),
.B2(n_309),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_470),
.B(n_444),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_452),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_465),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_466),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_558),
.B(n_285),
.C(n_169),
.Y(n_646)
);

AND2x4_ASAP7_75t_SL g647 ( 
.A(n_451),
.B(n_445),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_584),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_474),
.B(n_167),
.Y(n_649)
);

AOI221xp5_ASAP7_75t_L g650 ( 
.A1(n_568),
.A2(n_229),
.B1(n_309),
.B2(n_300),
.C(n_299),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_470),
.B(n_445),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_581),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_459),
.B(n_445),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_585),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_459),
.B(n_412),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_507),
.B(n_505),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_467),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_505),
.B(n_170),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_513),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_593),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_448),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_534),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_466),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_492),
.B(n_170),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_452),
.B(n_176),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_454),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_559),
.B(n_176),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_483),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_485),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_591),
.B(n_177),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_591),
.B(n_177),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_455),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_467),
.A2(n_179),
.B1(n_181),
.B2(n_183),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_485),
.B(n_384),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_521),
.B(n_537),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_574),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_462),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_485),
.B(n_179),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_521),
.B(n_181),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_485),
.B(n_519),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_471),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_537),
.B(n_183),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_557),
.A2(n_412),
.B1(n_438),
.B2(n_434),
.Y(n_684)
);

OAI22x1_ASAP7_75t_SL g685 ( 
.A1(n_573),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_472),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_519),
.B(n_520),
.Y(n_687)
);

AND2x2_ASAP7_75t_SL g688 ( 
.A(n_449),
.B(n_213),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_469),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_469),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_478),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_480),
.B(n_384),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_480),
.A2(n_283),
.B1(n_286),
.B2(n_299),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_557),
.A2(n_473),
.B1(n_594),
.B2(n_483),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_480),
.B(n_300),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_492),
.B(n_185),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_558),
.B(n_186),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_523),
.B(n_412),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_534),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_563),
.B(n_191),
.C(n_305),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_519),
.B(n_213),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_480),
.B(n_192),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_476),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_477),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_483),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_519),
.B(n_213),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_486),
.A2(n_302),
.B1(n_205),
.B2(n_206),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_574),
.B(n_412),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_538),
.B(n_421),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_519),
.B(n_213),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_538),
.A2(n_201),
.B1(n_212),
.B2(n_217),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_520),
.B(n_219),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_540),
.B(n_220),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_520),
.B(n_231),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_540),
.A2(n_546),
.B1(n_577),
.B2(n_563),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_487),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_504),
.B(n_232),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_546),
.B(n_238),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_508),
.B(n_421),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_562),
.B(n_242),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_556),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_488),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_564),
.B(n_384),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_504),
.B(n_245),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_556),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_573),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_594),
.A2(n_423),
.B1(n_438),
.B2(n_434),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_489),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_577),
.B(n_421),
.Y(n_729)
);

AND2x6_ASAP7_75t_L g730 ( 
.A(n_564),
.B(n_421),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_495),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_592),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_478),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_577),
.B(n_509),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_499),
.B(n_250),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_577),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_562),
.B(n_252),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_510),
.B(n_258),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_511),
.B(n_262),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_515),
.B(n_541),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_541),
.B(n_271),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_554),
.A2(n_387),
.B(n_388),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_562),
.B(n_304),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_484),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_484),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_539),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_533),
.B(n_13),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_561),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_578),
.A2(n_359),
.B1(n_363),
.B2(n_367),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_451),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_497),
.B(n_438),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_451),
.B(n_438),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_497),
.Y(n_753)
);

AND2x6_ASAP7_75t_L g754 ( 
.A(n_498),
.B(n_422),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_498),
.B(n_434),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_579),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_500),
.B(n_434),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_500),
.B(n_385),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_502),
.B(n_385),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_502),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_506),
.B(n_423),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_506),
.B(n_527),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_527),
.B(n_423),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_529),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_613),
.B(n_482),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_595),
.A2(n_553),
.B(n_516),
.C(n_494),
.Y(n_766)
);

AND2x2_ASAP7_75t_SL g767 ( 
.A(n_597),
.B(n_514),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_659),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_656),
.A2(n_501),
.B(n_516),
.C(n_494),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_659),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_680),
.A2(n_587),
.B(n_586),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_633),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_615),
.B(n_676),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_668),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_602),
.B(n_518),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_680),
.A2(n_587),
.B(n_586),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_596),
.B(n_523),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_687),
.A2(n_567),
.B(n_583),
.Y(n_778)
);

NAND3xp33_ASAP7_75t_L g779 ( 
.A(n_609),
.B(n_547),
.C(n_572),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_668),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_687),
.A2(n_669),
.B(n_643),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_648),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_615),
.B(n_457),
.Y(n_783)
);

NOR2x1_ASAP7_75t_R g784 ( 
.A(n_692),
.B(n_501),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_634),
.A2(n_567),
.B(n_583),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_634),
.A2(n_543),
.B(n_583),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_653),
.B(n_524),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_619),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_655),
.B(n_526),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_630),
.A2(n_551),
.B(n_490),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_606),
.A2(n_525),
.B(n_571),
.C(n_572),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_662),
.B(n_548),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_719),
.B(n_531),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_740),
.A2(n_543),
.B(n_490),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_762),
.A2(n_543),
.B(n_490),
.Y(n_795)
);

BUFx4f_ASAP7_75t_L g796 ( 
.A(n_692),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_603),
.A2(n_535),
.B(n_529),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_699),
.B(n_571),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_699),
.B(n_545),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_614),
.B(n_528),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_712),
.A2(n_551),
.B(n_560),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_734),
.A2(n_576),
.B1(n_565),
.B2(n_566),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_631),
.B(n_530),
.Y(n_803)
);

AOI21x1_ASAP7_75t_L g804 ( 
.A1(n_758),
.A2(n_535),
.B(n_530),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_623),
.B(n_552),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_614),
.B(n_549),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_747),
.A2(n_550),
.B(n_570),
.C(n_551),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_617),
.B(n_569),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_688),
.A2(n_580),
.B1(n_560),
.B2(n_569),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_712),
.A2(n_720),
.B(n_714),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_606),
.A2(n_569),
.B(n_560),
.C(n_589),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_605),
.A2(n_589),
.B(n_576),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_615),
.B(n_657),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_764),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_696),
.B(n_512),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_657),
.B(n_589),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_714),
.A2(n_387),
.B(n_383),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_636),
.B(n_512),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_649),
.B(n_512),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_720),
.A2(n_388),
.B(n_383),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_688),
.A2(n_363),
.B1(n_367),
.B2(n_368),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_632),
.A2(n_368),
.B(n_372),
.C(n_381),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_692),
.B(n_715),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_737),
.A2(n_388),
.B(n_575),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_737),
.A2(n_388),
.B(n_575),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_743),
.A2(n_582),
.B(n_575),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_664),
.B(n_512),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_659),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_601),
.A2(n_694),
.B1(n_599),
.B2(n_624),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_743),
.A2(n_582),
.B(n_575),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_625),
.A2(n_372),
.B(n_381),
.Y(n_831)
);

BUFx4f_ASAP7_75t_L g832 ( 
.A(n_647),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_697),
.B(n_576),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_764),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_726),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_709),
.B(n_667),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_708),
.B(n_512),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_652),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_670),
.B(n_512),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_611),
.A2(n_422),
.B(n_423),
.C(n_26),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_748),
.B(n_756),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_746),
.B(n_576),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_671),
.B(n_576),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_600),
.B(n_576),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_736),
.B(n_582),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_668),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_758),
.A2(n_759),
.B(n_742),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_732),
.B(n_713),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_736),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_599),
.A2(n_422),
.B(n_20),
.C(n_26),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_675),
.A2(n_422),
.B(n_442),
.C(n_425),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_759),
.A2(n_582),
.B(n_575),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_705),
.B(n_750),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_718),
.B(n_425),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_647),
.B(n_582),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_741),
.A2(n_385),
.B(n_425),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_705),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_654),
.A2(n_442),
.B(n_425),
.C(n_385),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_635),
.A2(n_385),
.B(n_425),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_660),
.B(n_442),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_650),
.B(n_14),
.C(n_20),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_620),
.A2(n_385),
.B(n_425),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_705),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_658),
.B(n_717),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_724),
.A2(n_384),
.B1(n_425),
.B2(n_442),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_622),
.A2(n_644),
.B(n_760),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_764),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_661),
.B(n_14),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_693),
.A2(n_27),
.B(n_28),
.C(n_31),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_646),
.A2(n_384),
.B1(n_425),
.B2(n_442),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_673),
.B(n_442),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_666),
.A2(n_442),
.B1(n_35),
.B2(n_36),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_695),
.B(n_442),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_672),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_702),
.B(n_34),
.Y(n_875)
);

CKINVDCx8_ASAP7_75t_R g876 ( 
.A(n_659),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_721),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_677),
.B(n_35),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_681),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_721),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_686),
.B(n_36),
.Y(n_881)
);

AO22x1_ASAP7_75t_L g882 ( 
.A1(n_752),
.A2(n_384),
.B1(n_442),
.B2(n_40),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_607),
.A2(n_645),
.B(n_629),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_703),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_604),
.B(n_384),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_638),
.A2(n_385),
.B(n_384),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_704),
.B(n_39),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_716),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_721),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_610),
.A2(n_385),
.B(n_384),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_722),
.A2(n_385),
.B(n_50),
.C(n_53),
.Y(n_891)
);

BUFx12f_ASAP7_75t_L g892 ( 
.A(n_729),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_626),
.B(n_700),
.C(n_641),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_SL g894 ( 
.A(n_604),
.B(n_384),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_711),
.B(n_49),
.Y(n_895)
);

AOI21xp33_ASAP7_75t_L g896 ( 
.A1(n_608),
.A2(n_50),
.B(n_54),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_728),
.A2(n_55),
.B(n_59),
.C(n_60),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_616),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_731),
.A2(n_61),
.B(n_76),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_679),
.B(n_154),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_598),
.B(n_82),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_618),
.A2(n_689),
.B(n_690),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_639),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_682),
.B(n_85),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_629),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_727),
.B(n_89),
.Y(n_906)
);

AOI21xp33_ASAP7_75t_L g907 ( 
.A1(n_612),
.A2(n_91),
.B(n_94),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_721),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_685),
.Y(n_909)
);

INVx3_ASAP7_75t_SL g910 ( 
.A(n_628),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_644),
.A2(n_97),
.B(n_98),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_621),
.A2(n_105),
.B1(n_121),
.B2(n_130),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_645),
.A2(n_133),
.B(n_137),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_663),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_707),
.B(n_138),
.C(n_144),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_663),
.B(n_145),
.Y(n_916)
);

AOI21xp33_ASAP7_75t_L g917 ( 
.A1(n_627),
.A2(n_147),
.B(n_640),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_735),
.B(n_738),
.C(n_739),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_639),
.B(n_683),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_689),
.A2(n_745),
.B(n_690),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_691),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_725),
.B(n_683),
.Y(n_922)
);

NOR2x2_ASAP7_75t_L g923 ( 
.A(n_691),
.B(n_753),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_733),
.B(n_745),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_733),
.A2(n_744),
.B(n_753),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_744),
.A2(n_760),
.B(n_642),
.C(n_651),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_628),
.A2(n_637),
.B(n_665),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_637),
.B(n_665),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_761),
.B(n_751),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_730),
.B(n_725),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_730),
.B(n_725),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_754),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_678),
.A2(n_757),
.B(n_755),
.C(n_698),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_730),
.B(n_684),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_730),
.B(n_678),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_749),
.B(n_701),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_754),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_730),
.B(n_754),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_730),
.B(n_754),
.Y(n_939)
);

AOI21xp33_ASAP7_75t_L g940 ( 
.A1(n_723),
.A2(n_674),
.B(n_701),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_706),
.B(n_710),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_754),
.B(n_723),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_754),
.A2(n_706),
.B(n_710),
.Y(n_943)
);

AOI33xp33_ASAP7_75t_L g944 ( 
.A1(n_674),
.A2(n_553),
.A3(n_568),
.B1(n_555),
.B2(n_538),
.B3(n_546),
.Y(n_944)
);

NOR2x1_ASAP7_75t_L g945 ( 
.A(n_656),
.B(n_467),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_619),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_636),
.A2(n_664),
.B(n_649),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_772),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_832),
.B(n_947),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_875),
.A2(n_766),
.B(n_900),
.C(n_779),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_796),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_841),
.A2(n_836),
.B(n_810),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_796),
.B(n_832),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_808),
.A2(n_928),
.B(n_799),
.C(n_893),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_803),
.A2(n_815),
.B(n_833),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_767),
.B(n_864),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_835),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_777),
.A2(n_945),
.B1(n_773),
.B2(n_765),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_785),
.A2(n_786),
.B(n_818),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_805),
.B(n_782),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_876),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_848),
.B(n_792),
.Y(n_962)
);

BUFx4f_ASAP7_75t_L g963 ( 
.A(n_863),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_892),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_788),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_787),
.A2(n_775),
.B1(n_789),
.B2(n_946),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_775),
.B(n_829),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_R g968 ( 
.A1(n_909),
.A2(n_783),
.B1(n_838),
.B2(n_874),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_903),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_879),
.A2(n_793),
.B1(n_821),
.B2(n_901),
.Y(n_970)
);

AO32x2_ASAP7_75t_L g971 ( 
.A1(n_872),
.A2(n_821),
.A3(n_809),
.B1(n_884),
.B2(n_888),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_819),
.A2(n_847),
.B(n_929),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_813),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_791),
.A2(n_769),
.B(n_944),
.C(n_918),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_800),
.B(n_798),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_868),
.A2(n_887),
.B1(n_878),
.B2(n_881),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_768),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_929),
.A2(n_790),
.B(n_795),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_827),
.B(n_910),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_853),
.B(n_774),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_840),
.A2(n_904),
.B(n_895),
.C(n_861),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_853),
.B(n_774),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_869),
.A2(n_884),
.B(n_888),
.C(n_807),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_823),
.A2(n_800),
.B1(n_806),
.B2(n_934),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_905),
.Y(n_985)
);

BUFx4f_ASAP7_75t_L g986 ( 
.A(n_853),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_844),
.B(n_885),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_932),
.B(n_780),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_914),
.B(n_898),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_921),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_771),
.A2(n_776),
.B(n_794),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_814),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_872),
.A2(n_891),
.B(n_850),
.C(n_896),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_849),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_801),
.A2(n_938),
.B(n_942),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_834),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_784),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_867),
.B(n_924),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_899),
.A2(n_843),
.B(n_927),
.C(n_842),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_768),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_860),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_942),
.A2(n_781),
.B(n_839),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_802),
.A2(n_932),
.B1(n_809),
.B2(n_906),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_899),
.A2(n_842),
.B(n_812),
.C(n_896),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_778),
.A2(n_866),
.B(n_856),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_860),
.A2(n_935),
.B1(n_806),
.B2(n_812),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_923),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_854),
.B(n_797),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_816),
.B(n_919),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_768),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_885),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_939),
.A2(n_837),
.B1(n_797),
.B2(n_931),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_915),
.A2(n_851),
.B(n_858),
.C(n_811),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_L g1014 ( 
.A1(n_831),
.A2(n_871),
.B(n_933),
.C(n_940),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_925),
.B(n_873),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_770),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_780),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_846),
.B(n_857),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_R g1019 ( 
.A(n_846),
.B(n_857),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_925),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_883),
.B(n_920),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_940),
.A2(n_926),
.B(n_930),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_804),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_770),
.B(n_908),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_SL g1025 ( 
.A1(n_912),
.A2(n_913),
.B1(n_880),
.B2(n_889),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_822),
.A2(n_897),
.B(n_936),
.C(n_912),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_902),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_SL g1028 ( 
.A(n_880),
.B(n_894),
.Y(n_1028)
);

AO32x1_ASAP7_75t_L g1029 ( 
.A1(n_937),
.A2(n_913),
.A3(n_882),
.B1(n_907),
.B2(n_859),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_828),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_877),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_877),
.B(n_908),
.Y(n_1032)
);

AOI33xp33_ASAP7_75t_L g1033 ( 
.A1(n_870),
.A2(n_865),
.A3(n_820),
.B1(n_817),
.B2(n_907),
.B3(n_862),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_855),
.B(n_922),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_917),
.B(n_943),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_916),
.A2(n_917),
.B(n_825),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_916),
.A2(n_824),
.B(n_826),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_941),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_845),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_911),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_943),
.A2(n_890),
.B(n_886),
.C(n_830),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_852),
.B(n_597),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_772),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_947),
.A2(n_597),
.B1(n_609),
.B2(n_767),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_832),
.B(n_534),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_947),
.B(n_597),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_841),
.A2(n_634),
.B(n_836),
.Y(n_1047)
);

BUFx8_ASAP7_75t_SL g1048 ( 
.A(n_772),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_832),
.B(n_517),
.Y(n_1049)
);

AOI22x1_ASAP7_75t_L g1050 ( 
.A1(n_790),
.A2(n_810),
.B1(n_927),
.B2(n_794),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_841),
.A2(n_634),
.B(n_836),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_841),
.A2(n_947),
.B(n_634),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_947),
.A2(n_597),
.B1(n_765),
.B2(n_688),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_813),
.B(n_945),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_847),
.A2(n_804),
.B(n_859),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_947),
.A2(n_597),
.B1(n_765),
.B2(n_688),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_813),
.B(n_945),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_832),
.B(n_534),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_836),
.B(n_656),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_947),
.A2(n_595),
.B(n_597),
.C(n_667),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_841),
.A2(n_634),
.B(n_836),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_841),
.A2(n_634),
.B(n_836),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_796),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_835),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_796),
.B(n_668),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_841),
.A2(n_634),
.B(n_836),
.Y(n_1066)
);

CKINVDCx14_ASAP7_75t_R g1067 ( 
.A(n_772),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_947),
.B(n_597),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_841),
.A2(n_947),
.B(n_634),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_767),
.B(n_597),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_836),
.B(n_656),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_841),
.A2(n_947),
.B(n_634),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_810),
.A2(n_927),
.B(n_831),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_947),
.A2(n_597),
.B1(n_765),
.B2(n_688),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_947),
.A2(n_595),
.B(n_597),
.C(n_667),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_947),
.A2(n_595),
.B(n_597),
.C(n_667),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_767),
.B(n_597),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_832),
.B(n_534),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_772),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_947),
.B(n_597),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_808),
.A2(n_613),
.B(n_450),
.C(n_463),
.Y(n_1081)
);

AO21x2_ASAP7_75t_L g1082 ( 
.A1(n_1036),
.A2(n_1037),
.B(n_1035),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_965),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1046),
.A2(n_1068),
.B(n_1080),
.C(n_1081),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1086)
);

OAI22x1_ASAP7_75t_L g1087 ( 
.A1(n_1044),
.A2(n_1070),
.B1(n_1077),
.B2(n_956),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1069),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_958),
.A2(n_1007),
.B1(n_984),
.B2(n_968),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_963),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_957),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_959),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_953),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_960),
.B(n_975),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1052),
.A2(n_1069),
.B(n_1072),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_1004),
.A2(n_1023),
.A3(n_950),
.B(n_999),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_995),
.A2(n_1041),
.B(n_1005),
.Y(n_1097)
);

AOI221x1_ASAP7_75t_L g1098 ( 
.A1(n_1053),
.A2(n_1074),
.B1(n_1056),
.B2(n_981),
.C(n_976),
.Y(n_1098)
);

AO32x2_ASAP7_75t_L g1099 ( 
.A1(n_1053),
.A2(n_1056),
.A3(n_1074),
.B1(n_966),
.B2(n_976),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1005),
.A2(n_991),
.B(n_978),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1050),
.A2(n_1022),
.B(n_1073),
.Y(n_1101)
);

AO21x2_ASAP7_75t_L g1102 ( 
.A1(n_955),
.A2(n_972),
.B(n_1008),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1060),
.A2(n_1076),
.B(n_1075),
.C(n_1042),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1047),
.A2(n_1066),
.B(n_1051),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

AO21x1_ASAP7_75t_L g1106 ( 
.A1(n_966),
.A2(n_970),
.B(n_1026),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1063),
.B(n_951),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1061),
.A2(n_1062),
.B(n_952),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_985),
.Y(n_1109)
);

AOI211x1_ASAP7_75t_L g1110 ( 
.A1(n_949),
.A2(n_962),
.B(n_1045),
.C(n_1078),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1003),
.A2(n_1025),
.B(n_954),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1021),
.A2(n_1027),
.B(n_1014),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_SL g1113 ( 
.A1(n_983),
.A2(n_993),
.B1(n_974),
.B2(n_970),
.C(n_1001),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_990),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1021),
.A2(n_1012),
.B(n_1013),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1003),
.A2(n_1006),
.B(n_1008),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1064),
.Y(n_1117)
);

BUFx4f_ASAP7_75t_SL g1118 ( 
.A(n_1079),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_967),
.A2(n_1040),
.B(n_1009),
.C(n_1034),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_SL g1120 ( 
.A(n_1049),
.B(n_1058),
.C(n_1010),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1006),
.A2(n_1029),
.B(n_1012),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1029),
.A2(n_1015),
.B(n_967),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1029),
.A2(n_1015),
.B(n_1020),
.Y(n_1123)
);

AOI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_1038),
.A2(n_998),
.B(n_989),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_997),
.A2(n_979),
.B1(n_987),
.B2(n_1063),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1018),
.A2(n_1028),
.B(n_988),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1032),
.A2(n_1017),
.B(n_1024),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_992),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_961),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_1033),
.A3(n_1030),
.B(n_971),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_961),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_973),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_994),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_1054),
.A2(n_1057),
.B(n_971),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_969),
.A2(n_1011),
.B(n_982),
.C(n_980),
.Y(n_1135)
);

NOR2x1_ASAP7_75t_SL g1136 ( 
.A(n_1039),
.B(n_977),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_L g1137 ( 
.A(n_1019),
.B(n_951),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_986),
.A2(n_982),
.B(n_980),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1065),
.A2(n_986),
.B(n_971),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1016),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1039),
.A2(n_977),
.B(n_1031),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1039),
.A2(n_977),
.B(n_1031),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_964),
.B(n_987),
.Y(n_1143)
);

OAI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_948),
.A2(n_1043),
.B1(n_963),
.B2(n_951),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1048),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1057),
.B(n_1068),
.C(n_1046),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1067),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1079),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1070),
.B(n_1077),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_961),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1046),
.B(n_1080),
.C(n_1068),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_1053),
.A2(n_1056),
.A3(n_1074),
.B1(n_966),
.B2(n_872),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1070),
.B(n_1077),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1069),
.Y(n_1155)
);

AOI221xp5_ASAP7_75t_SL g1156 ( 
.A1(n_983),
.A2(n_947),
.B1(n_1046),
.B2(n_1080),
.C(n_1068),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_963),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1046),
.A2(n_1068),
.B(n_1080),
.C(n_947),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_963),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_959),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1068),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1068),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1081),
.A2(n_947),
.B(n_950),
.C(n_1046),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_959),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1053),
.A2(n_1074),
.B(n_1056),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1046),
.A2(n_1068),
.B(n_1080),
.C(n_947),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1079),
.Y(n_1168)
);

OA22x2_ASAP7_75t_L g1169 ( 
.A1(n_1044),
.A2(n_1070),
.B1(n_1077),
.B2(n_715),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_961),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_965),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1036),
.A2(n_1005),
.B(n_978),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_953),
.B(n_961),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1046),
.B(n_1080),
.C(n_1068),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1052),
.A2(n_947),
.B(n_1069),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1036),
.A2(n_1004),
.A3(n_1023),
.B(n_950),
.Y(n_1177)
);

INVx3_ASAP7_75t_SL g1178 ( 
.A(n_948),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_959),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_965),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1069),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_961),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1048),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1063),
.B(n_951),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1052),
.A2(n_947),
.B(n_1069),
.Y(n_1186)
);

AOI221xp5_ASAP7_75t_SL g1187 ( 
.A1(n_983),
.A2(n_947),
.B1(n_1046),
.B2(n_1080),
.C(n_1068),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1036),
.A2(n_1005),
.B(n_978),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1052),
.A2(n_947),
.B(n_1069),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1052),
.A2(n_947),
.B(n_1069),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1068),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_SL g1193 ( 
.A1(n_1081),
.A2(n_947),
.B(n_950),
.C(n_1046),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1069),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1069),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1070),
.B(n_1077),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1052),
.A2(n_947),
.B(n_1069),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_959),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1036),
.A2(n_1004),
.A3(n_1023),
.B(n_950),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_963),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_959),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1068),
.C(n_947),
.Y(n_1202)
);

AO22x2_ASAP7_75t_L g1203 ( 
.A1(n_1053),
.A2(n_1074),
.B1(n_1056),
.B2(n_1070),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_961),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1036),
.A2(n_1004),
.A3(n_1023),
.B(n_950),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1068),
.C(n_947),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_963),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1069),
.Y(n_1208)
);

AOI21xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1046),
.A2(n_1080),
.B(n_1068),
.Y(n_1209)
);

CKINVDCx11_ASAP7_75t_R g1210 ( 
.A(n_1079),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1036),
.A2(n_1004),
.A3(n_1023),
.B(n_950),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1079),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_1129),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1117),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1169),
.A2(n_1203),
.B1(n_1173),
.B2(n_1191),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1083),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_SL g1217 ( 
.A1(n_1087),
.A2(n_1192),
.B1(n_1162),
.B2(n_1161),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1169),
.A2(n_1203),
.B1(n_1165),
.B2(n_1106),
.Y(n_1218)
);

BUFx10_ASAP7_75t_L g1219 ( 
.A(n_1184),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_SL g1220 ( 
.A(n_1090),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1168),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1210),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1200),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1161),
.A2(n_1192),
.B1(n_1162),
.B2(n_1175),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1089),
.A2(n_1154),
.B1(n_1147),
.B2(n_1143),
.Y(n_1225)
);

CKINVDCx11_ASAP7_75t_R g1226 ( 
.A(n_1212),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1183),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_1207),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1211),
.Y(n_1229)
);

INVx8_ASAP7_75t_L g1230 ( 
.A(n_1183),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1152),
.A2(n_1175),
.B1(n_1146),
.B2(n_1196),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1152),
.A2(n_1146),
.B1(n_1084),
.B2(n_1182),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1148),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1158),
.A2(n_1166),
.B1(n_1209),
.B2(n_1103),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1084),
.B(n_1086),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1149),
.A2(n_1167),
.B1(n_1182),
.B2(n_1086),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1171),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1118),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1202),
.A2(n_1206),
.B1(n_1085),
.B2(n_1111),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_1157),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_SL g1241 ( 
.A(n_1145),
.Y(n_1241)
);

BUFx2_ASAP7_75t_SL g1242 ( 
.A(n_1183),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1178),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1151),
.A2(n_1167),
.B1(n_1134),
.B2(n_1094),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1180),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1151),
.B(n_1156),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1105),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1110),
.A2(n_1091),
.B1(n_1116),
.B2(n_1119),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1120),
.A2(n_1109),
.B1(n_1128),
.B2(n_1114),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1091),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1133),
.A2(n_1124),
.B1(n_1132),
.B2(n_1125),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1131),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1131),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1125),
.A2(n_1156),
.B1(n_1187),
.B2(n_1189),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1098),
.A2(n_1139),
.B1(n_1099),
.B2(n_1153),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1187),
.A2(n_1190),
.B1(n_1186),
.B2(n_1197),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1147),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_1159),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1131),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1093),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1176),
.A2(n_1121),
.B1(n_1138),
.B2(n_1174),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1170),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1113),
.B(n_1170),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1130),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1150),
.B(n_1204),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1124),
.A2(n_1122),
.B1(n_1099),
.B2(n_1153),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1095),
.A2(n_1194),
.B1(n_1208),
.B2(n_1195),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1095),
.A2(n_1194),
.B1(n_1208),
.B2(n_1195),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1140),
.A2(n_1137),
.B1(n_1122),
.B2(n_1204),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1107),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1136),
.A2(n_1115),
.B1(n_1107),
.B2(n_1185),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1123),
.A2(n_1185),
.B1(n_1144),
.B2(n_1102),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1127),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1163),
.B(n_1193),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1123),
.A2(n_1102),
.B1(n_1126),
.B2(n_1181),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1155),
.A2(n_1181),
.B1(n_1088),
.B2(n_1135),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1141),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1142),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1112),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_SL g1280 ( 
.A1(n_1155),
.A2(n_1104),
.B(n_1108),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1172),
.A2(n_1188),
.B1(n_1104),
.B2(n_1096),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1082),
.A2(n_1188),
.B1(n_1172),
.B2(n_1101),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1211),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1082),
.A2(n_1100),
.B1(n_1097),
.B2(n_1096),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1177),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1177),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1211),
.B(n_1205),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1092),
.A2(n_1160),
.B(n_1164),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1199),
.B(n_1205),
.Y(n_1289)
);

INVx3_ASAP7_75t_SL g1290 ( 
.A(n_1179),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1198),
.A2(n_597),
.B1(n_1077),
.B2(n_1070),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1201),
.A2(n_1044),
.B1(n_1098),
.B2(n_1068),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1168),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1090),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1177),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1098),
.A2(n_1044),
.B1(n_1068),
.B2(n_1046),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_SL g1297 ( 
.A(n_1148),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1169),
.A2(n_597),
.B1(n_1077),
.B2(n_1070),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_SL g1299 ( 
.A(n_1148),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1098),
.A2(n_1044),
.B1(n_1068),
.B2(n_1046),
.Y(n_1300)
);

OAI22x1_ASAP7_75t_SL g1301 ( 
.A1(n_1184),
.A2(n_573),
.B1(n_342),
.B2(n_347),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1169),
.A2(n_597),
.B1(n_557),
.B2(n_767),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1169),
.A2(n_597),
.B1(n_557),
.B2(n_767),
.Y(n_1303)
);

BUFx10_ASAP7_75t_L g1304 ( 
.A(n_1184),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1168),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1083),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1169),
.A2(n_597),
.B1(n_1077),
.B2(n_1070),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1158),
.A2(n_1046),
.B1(n_1080),
.B2(n_1068),
.Y(n_1308)
);

OAI21xp33_ASAP7_75t_L g1309 ( 
.A1(n_1158),
.A2(n_1068),
.B(n_1046),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1117),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1091),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1169),
.A2(n_597),
.B1(n_1077),
.B2(n_1070),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1083),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1168),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1117),
.Y(n_1315)
);

BUFx4f_ASAP7_75t_L g1316 ( 
.A(n_1148),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1285),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1264),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1281),
.A2(n_1287),
.B(n_1286),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1288),
.A2(n_1268),
.B(n_1267),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1278),
.B(n_1277),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1229),
.B(n_1283),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1232),
.B(n_1246),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1302),
.A2(n_1303),
.B1(n_1298),
.B2(n_1312),
.Y(n_1324)
);

NOR2x1_ASAP7_75t_SL g1325 ( 
.A(n_1248),
.B(n_1261),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1229),
.B(n_1283),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1289),
.B(n_1224),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1224),
.B(n_1235),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1256),
.A2(n_1276),
.B(n_1282),
.Y(n_1329)
);

CKINVDCx12_ASAP7_75t_R g1330 ( 
.A(n_1225),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1295),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1295),
.Y(n_1332)
);

BUFx4f_ASAP7_75t_SL g1333 ( 
.A(n_1221),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1266),
.B(n_1255),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1216),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1237),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1245),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1239),
.A2(n_1274),
.B(n_1234),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1308),
.A2(n_1296),
.B1(n_1300),
.B2(n_1263),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1306),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1280),
.A2(n_1281),
.B(n_1292),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1279),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1230),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1266),
.B(n_1275),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1313),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1244),
.B(n_1214),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1290),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1290),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1310),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1275),
.B(n_1284),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1226),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1315),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1284),
.B(n_1282),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1244),
.B(n_1231),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1254),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1231),
.B(n_1236),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1233),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1222),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1218),
.A2(n_1272),
.B(n_1215),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1218),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1250),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1311),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1217),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1273),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1260),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1309),
.B(n_1228),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1223),
.B(n_1294),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1292),
.A2(n_1296),
.B(n_1300),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1272),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1215),
.B(n_1251),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1251),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1291),
.B(n_1312),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1269),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1298),
.A2(n_1307),
.B1(n_1291),
.B2(n_1249),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1270),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1344),
.B(n_1307),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1339),
.A2(n_1305),
.B(n_1293),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1368),
.A2(n_1230),
.B(n_1271),
.C(n_1262),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1349),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1364),
.B(n_1247),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1361),
.B(n_1257),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1335),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1349),
.B(n_1243),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1339),
.A2(n_1265),
.B(n_1227),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1368),
.A2(n_1230),
.B(n_1242),
.C(n_1259),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1338),
.A2(n_1316),
.B(n_1243),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1352),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1363),
.A2(n_1316),
.B(n_1213),
.C(n_1220),
.Y(n_1388)
);

AO22x2_ASAP7_75t_L g1389 ( 
.A1(n_1371),
.A2(n_1301),
.B1(n_1294),
.B2(n_1223),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1362),
.B(n_1228),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1338),
.A2(n_1238),
.B(n_1220),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1341),
.A2(n_1329),
.B(n_1320),
.Y(n_1392)
);

AO21x1_ASAP7_75t_L g1393 ( 
.A1(n_1323),
.A2(n_1253),
.B(n_1252),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1355),
.B(n_1253),
.C(n_1252),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1321),
.B(n_1213),
.Y(n_1395)
);

OAI211xp5_ASAP7_75t_L g1396 ( 
.A1(n_1323),
.A2(n_1241),
.B(n_1299),
.C(n_1297),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1363),
.A2(n_1240),
.B(n_1258),
.C(n_1241),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1328),
.B(n_1258),
.Y(n_1398)
);

AO32x2_ASAP7_75t_L g1399 ( 
.A1(n_1346),
.A2(n_1297),
.A3(n_1299),
.B1(n_1314),
.B2(n_1304),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1327),
.B(n_1219),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1317),
.B(n_1219),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1355),
.A2(n_1328),
.B(n_1341),
.C(n_1354),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1321),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1369),
.A2(n_1371),
.B(n_1325),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1369),
.A2(n_1325),
.B(n_1344),
.Y(n_1405)
);

AOI211xp5_ASAP7_75t_L g1406 ( 
.A1(n_1354),
.A2(n_1356),
.B(n_1366),
.C(n_1373),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1358),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1408)
);

AND2x2_ASAP7_75t_SL g1409 ( 
.A(n_1317),
.B(n_1370),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1410)
);

OAI31xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1372),
.A2(n_1373),
.A3(n_1334),
.B(n_1350),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1372),
.A2(n_1374),
.B(n_1356),
.C(n_1359),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1326),
.B(n_1375),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1331),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1372),
.A2(n_1329),
.B(n_1359),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1367),
.B(n_1337),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1331),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1329),
.A2(n_1359),
.B(n_1350),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1324),
.A2(n_1330),
.B1(n_1360),
.B2(n_1370),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1408),
.B(n_1353),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1408),
.B(n_1353),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1382),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1410),
.B(n_1353),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1379),
.B(n_1340),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1410),
.B(n_1320),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1415),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1379),
.B(n_1345),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1410),
.B(n_1342),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1392),
.B(n_1342),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1415),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1403),
.B(n_1348),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1376),
.A2(n_1360),
.B1(n_1357),
.B2(n_1319),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1414),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1376),
.A2(n_1357),
.B1(n_1319),
.B2(n_1345),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1418),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1401),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1419),
.B(n_1347),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1416),
.B(n_1413),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_SL g1440 ( 
.A(n_1401),
.B(n_1319),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1412),
.A2(n_1340),
.B1(n_1332),
.B2(n_1365),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1404),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1377),
.B(n_1347),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1420),
.A2(n_1319),
.B1(n_1333),
.B2(n_1318),
.Y(n_1444)
);

OAI211xp5_ASAP7_75t_L g1445 ( 
.A1(n_1435),
.A2(n_1402),
.B(n_1411),
.C(n_1397),
.Y(n_1445)
);

AOI31xp33_ASAP7_75t_L g1446 ( 
.A1(n_1441),
.A2(n_1402),
.A3(n_1406),
.B(n_1397),
.Y(n_1446)
);

INVxp33_ASAP7_75t_L g1447 ( 
.A(n_1443),
.Y(n_1447)
);

OAI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1441),
.A2(n_1412),
.B1(n_1378),
.B2(n_1385),
.C(n_1384),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1425),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1427),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1430),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1427),
.B(n_1387),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1431),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1431),
.Y(n_1454)
);

NAND4xp25_ASAP7_75t_L g1455 ( 
.A(n_1441),
.B(n_1398),
.C(n_1383),
.D(n_1387),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1428),
.Y(n_1458)
);

OAI31xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1443),
.A2(n_1394),
.A3(n_1386),
.B(n_1396),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1437),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1436),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1428),
.B(n_1405),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1432),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1430),
.Y(n_1464)
);

OAI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1435),
.A2(n_1378),
.B1(n_1385),
.B2(n_1391),
.C(n_1388),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1444),
.A2(n_1409),
.B1(n_1400),
.B2(n_1417),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1421),
.B(n_1409),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1437),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1437),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1428),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1421),
.B(n_1381),
.Y(n_1471)
);

AND2x4_ASAP7_75t_SL g1472 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1429),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1446),
.B(n_1393),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1474),
.B(n_1422),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1474),
.B(n_1424),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1451),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1468),
.B(n_1442),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1456),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1449),
.B(n_1434),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1467),
.B(n_1426),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1463),
.B(n_1440),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1457),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1464),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1457),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1450),
.B(n_1423),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1467),
.B(n_1426),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1458),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1458),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1468),
.Y(n_1492)
);

AOI211xp5_ASAP7_75t_L g1493 ( 
.A1(n_1448),
.A2(n_1388),
.B(n_1380),
.C(n_1399),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1446),
.B(n_1438),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1495)
);

NOR2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1455),
.B(n_1343),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1455),
.B(n_1407),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1450),
.B(n_1423),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1488),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1479),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1494),
.B(n_1470),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1488),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1498),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1498),
.Y(n_1505)
);

OAI32xp33_ASAP7_75t_L g1506 ( 
.A1(n_1494),
.A2(n_1447),
.A3(n_1448),
.B1(n_1466),
.B2(n_1462),
.Y(n_1506)
);

AOI21xp33_ASAP7_75t_L g1507 ( 
.A1(n_1475),
.A2(n_1445),
.B(n_1459),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1478),
.B(n_1453),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1479),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1479),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1478),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_1475),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1493),
.B(n_1459),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1492),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1483),
.B(n_1472),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1482),
.B(n_1452),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1489),
.B(n_1472),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1472),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1478),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1481),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1481),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1489),
.B(n_1461),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1479),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1453),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1485),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1485),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1485),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1487),
.B(n_1454),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1487),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1482),
.B(n_1452),
.Y(n_1535)
);

AND2x4_ASAP7_75t_SL g1536 ( 
.A(n_1484),
.B(n_1471),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1487),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1476),
.B(n_1460),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1482),
.B(n_1462),
.Y(n_1540)
);

AOI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1507),
.A2(n_1497),
.B(n_1493),
.C(n_1445),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1490),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1490),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1492),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1532),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1351),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1516),
.B(n_1496),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1493),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1532),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1517),
.B(n_1490),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1496),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1519),
.B(n_1484),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1536),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1529),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1532),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1538),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1511),
.Y(n_1557)
);

AND3x2_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1333),
.C(n_1390),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1496),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1515),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1517),
.B(n_1491),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1522),
.Y(n_1563)
);

NAND2x1p5_ASAP7_75t_L g1564 ( 
.A(n_1529),
.B(n_1492),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1522),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1523),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1515),
.Y(n_1567)
);

NAND2x1_ASAP7_75t_SL g1568 ( 
.A(n_1525),
.B(n_1484),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1520),
.B(n_1476),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1515),
.B(n_1495),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1506),
.B(n_1407),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1523),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1501),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1524),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1501),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1546),
.B(n_1544),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1548),
.B(n_1539),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1557),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1546),
.B(n_1520),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1557),
.Y(n_1580)
);

AOI21xp33_ASAP7_75t_L g1581 ( 
.A1(n_1541),
.A2(n_1506),
.B(n_1524),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1561),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_SL g1583 ( 
.A1(n_1541),
.A2(n_1502),
.B(n_1469),
.C(n_1535),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1554),
.B(n_1539),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1544),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1571),
.A2(n_1502),
.B(n_1525),
.Y(n_1586)
);

OAI32xp33_ASAP7_75t_L g1587 ( 
.A1(n_1552),
.A2(n_1480),
.A3(n_1535),
.B1(n_1518),
.B2(n_1540),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1567),
.B(n_1539),
.Y(n_1588)
);

OAI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1568),
.A2(n_1465),
.B1(n_1433),
.B2(n_1466),
.C(n_1444),
.Y(n_1589)
);

O2A1O1Ixp5_ASAP7_75t_L g1590 ( 
.A1(n_1553),
.A2(n_1544),
.B(n_1549),
.C(n_1545),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1499),
.Y(n_1591)
);

AOI31xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1545),
.A2(n_1540),
.A3(n_1533),
.B(n_1508),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1568),
.A2(n_1512),
.B(n_1500),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1553),
.B(n_1499),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1544),
.Y(n_1595)
);

OAI322xp33_ASAP7_75t_L g1596 ( 
.A1(n_1542),
.A2(n_1504),
.A3(n_1505),
.B1(n_1503),
.B2(n_1480),
.C1(n_1527),
.C2(n_1508),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1549),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1556),
.A2(n_1503),
.B1(n_1504),
.B2(n_1505),
.C(n_1510),
.Y(n_1598)
);

XNOR2xp5_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1389),
.Y(n_1599)
);

NAND2x2_ASAP7_75t_L g1600 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1582),
.B(n_1556),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1597),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1591),
.Y(n_1604)
);

OAI211xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1583),
.A2(n_1543),
.B(n_1553),
.C(n_1555),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_L g1606 ( 
.A(n_1583),
.B(n_1575),
.C(n_1573),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1578),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1589),
.A2(n_1570),
.B1(n_1555),
.B2(n_1547),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1569),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1585),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1600),
.A2(n_1570),
.B1(n_1550),
.B2(n_1562),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1580),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1591),
.B(n_1569),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1596),
.A2(n_1575),
.B1(n_1573),
.B2(n_1574),
.C(n_1572),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1584),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_SL g1616 ( 
.A1(n_1600),
.A2(n_1440),
.B1(n_1570),
.B2(n_1547),
.Y(n_1616)
);

OAI32xp33_ASAP7_75t_L g1617 ( 
.A1(n_1586),
.A2(n_1564),
.A3(n_1550),
.B1(n_1562),
.B2(n_1480),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1595),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1594),
.B(n_1477),
.Y(n_1619)
);

AOI32xp33_ASAP7_75t_L g1620 ( 
.A1(n_1605),
.A2(n_1611),
.A3(n_1603),
.B1(n_1608),
.B2(n_1606),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1610),
.Y(n_1621)
);

NOR2xp67_ASAP7_75t_L g1622 ( 
.A(n_1610),
.B(n_1588),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1609),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1603),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1601),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1594),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1604),
.B(n_1613),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1607),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1615),
.B(n_1579),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1619),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1625),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1625),
.B(n_1611),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_SL g1634 ( 
.A(n_1620),
.B(n_1616),
.C(n_1614),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1627),
.A2(n_1598),
.B(n_1593),
.C(n_1612),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_L g1636 ( 
.A(n_1621),
.B(n_1592),
.Y(n_1636)
);

NOR2xp67_ASAP7_75t_L g1637 ( 
.A(n_1623),
.B(n_1579),
.Y(n_1637)
);

AOI211x1_ASAP7_75t_SL g1638 ( 
.A1(n_1622),
.A2(n_1617),
.B(n_1587),
.C(n_1564),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1623),
.B(n_1551),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1628),
.B(n_1564),
.Y(n_1640)
);

OAI21xp33_ASAP7_75t_L g1641 ( 
.A1(n_1634),
.A2(n_1630),
.B(n_1631),
.Y(n_1641)
);

OAI211xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1638),
.A2(n_1626),
.B(n_1624),
.C(n_1629),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1643)
);

OAI21xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1636),
.A2(n_1559),
.B(n_1551),
.Y(n_1644)
);

NAND2xp33_ASAP7_75t_SL g1645 ( 
.A(n_1633),
.B(n_1559),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1643),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1641),
.A2(n_1632),
.B1(n_1635),
.B2(n_1599),
.Y(n_1647)
);

AOI221x1_ASAP7_75t_L g1648 ( 
.A1(n_1642),
.A2(n_1640),
.B1(n_1639),
.B2(n_1574),
.C(n_1572),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1645),
.B(n_1644),
.C(n_1563),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1641),
.B(n_1560),
.Y(n_1650)
);

O2A1O1Ixp5_ASAP7_75t_L g1651 ( 
.A1(n_1645),
.A2(n_1566),
.B(n_1565),
.C(n_1563),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1651),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1650),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1646),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1648),
.B(n_1566),
.Y(n_1655)
);

NOR2xp67_ASAP7_75t_L g1656 ( 
.A(n_1647),
.B(n_1560),
.Y(n_1656)
);

OAI322xp33_ASAP7_75t_L g1657 ( 
.A1(n_1652),
.A2(n_1649),
.A3(n_1565),
.B1(n_1480),
.B2(n_1510),
.C1(n_1526),
.C2(n_1509),
.Y(n_1657)
);

AOI221x1_ASAP7_75t_L g1658 ( 
.A1(n_1654),
.A2(n_1518),
.B1(n_1528),
.B2(n_1534),
.C(n_1530),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1656),
.A2(n_1537),
.B1(n_1509),
.B2(n_1501),
.C(n_1526),
.Y(n_1659)
);

OAI22x1_ASAP7_75t_L g1660 ( 
.A1(n_1657),
.A2(n_1653),
.B1(n_1655),
.B2(n_1518),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1660),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1659),
.B1(n_1658),
.B2(n_1537),
.Y(n_1662)
);

OA22x2_ASAP7_75t_L g1663 ( 
.A1(n_1662),
.A2(n_1518),
.B1(n_1528),
.B2(n_1534),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_1531),
.B(n_1530),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1526),
.B(n_1531),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1665),
.B(n_1389),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1666),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1389),
.B1(n_1525),
.B2(n_1500),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_R g1669 ( 
.A1(n_1668),
.A2(n_1512),
.B(n_1521),
.C(n_1399),
.Y(n_1669)
);


endmodule