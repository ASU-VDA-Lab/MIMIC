module fake_jpeg_8830_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_21),
.B(n_25),
.CON(n_41),
.SN(n_41)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_25),
.CON(n_47),
.SN(n_47)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_39),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_50),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_33),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_55),
.B1(n_35),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_64),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_33),
.B1(n_27),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_46),
.B1(n_45),
.B2(n_34),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_79),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_86),
.B(n_18),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_91),
.B1(n_31),
.B2(n_28),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_42),
.A3(n_19),
.B1(n_28),
.B2(n_39),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_89),
.A3(n_59),
.B1(n_65),
.B2(n_64),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_44),
.B(n_37),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_39),
.B1(n_36),
.B2(n_32),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_36),
.B1(n_34),
.B2(n_23),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_75),
.B1(n_34),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_25),
.B1(n_31),
.B2(n_18),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_107),
.B1(n_112),
.B2(n_45),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_49),
.B1(n_63),
.B2(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_49),
.B1(n_56),
.B2(n_50),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_114),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_63),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_70),
.B(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_84),
.B(n_31),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_86),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_79),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_125),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_71),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_90),
.A3(n_74),
.B1(n_81),
.B2(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_136),
.B(n_32),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_97),
.B1(n_77),
.B2(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_134),
.B1(n_139),
.B2(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_78),
.B1(n_89),
.B2(n_65),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_78),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_65),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_28),
.B1(n_80),
.B2(n_20),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_32),
.Y(n_161)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_149),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_108),
.B1(n_112),
.B2(n_135),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_159),
.B1(n_160),
.B2(n_166),
.Y(n_176)
);

CKINVDCx10_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_153),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_131),
.B(n_133),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_119),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_124),
.B1(n_136),
.B2(n_28),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_161),
.B(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_30),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_0),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_165),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_166)
);

AO21x2_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_130),
.B(n_136),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_156),
.B(n_159),
.C(n_163),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_120),
.C(n_125),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_179),
.C(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_174),
.B(n_175),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_185),
.B1(n_189),
.B2(n_20),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_87),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_67),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_187),
.C(n_188),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_67),
.B1(n_30),
.B2(n_27),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_67),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_151),
.C(n_143),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_153),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_165),
.C(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_206),
.B(n_209),
.Y(n_216)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_144),
.B1(n_142),
.B2(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_204),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_162),
.C(n_147),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_210),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_166),
.B(n_142),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_0),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_1),
.B(n_2),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_1),
.B(n_2),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_181),
.B1(n_178),
.B2(n_186),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_190),
.Y(n_235)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_200),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_177),
.B1(n_171),
.B2(n_180),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_222),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_188),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_185),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_202),
.C(n_205),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_210),
.B(n_209),
.Y(n_229)
);

OAI211xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_239),
.B(n_236),
.C(n_224),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_234),
.C(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_198),
.B1(n_189),
.B2(n_211),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_233),
.A2(n_229),
.B1(n_220),
.B2(n_234),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_197),
.C(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_237),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_198),
.C(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_206),
.B(n_198),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_228),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_221),
.B1(n_214),
.B2(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_224),
.C(n_227),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_217),
.C(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_219),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_248),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_249),
.A2(n_251),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_230),
.B1(n_217),
.B2(n_241),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_3),
.C(n_5),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_257),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_6),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_6),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_132),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_259),
.A2(n_242),
.B(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_263),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_246),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_252),
.A2(n_8),
.B(n_10),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_258),
.B(n_255),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_269),
.B1(n_262),
.B2(n_10),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_254),
.B(n_256),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_271),
.B(n_272),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_8),
.B(n_11),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_12),
.C(n_13),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_273),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_12),
.C(n_14),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_14),
.Y(n_276)
);


endmodule