module fake_netlist_5_349_n_180 (n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_180);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_180;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_122;
wire n_82;
wire n_142;
wire n_176;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_146;
wire n_143;
wire n_132;
wire n_83;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_29;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_147;
wire n_54;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_64;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_97;
wire n_63;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx2_ASAP7_75t_SL g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_35),
.Y(n_84)
);

OR2x6_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2x1p5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_32),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_32),
.B1(n_51),
.B2(n_8),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_71),
.B(n_72),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_53),
.B(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_70),
.B1(n_55),
.B2(n_52),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_53),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

O2A1O1Ixp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_96),
.B(n_99),
.C(n_100),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_79),
.B(n_73),
.C(n_80),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

CKINVDCx6p67_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_87),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_75),
.Y(n_108)
);

NAND2x1p5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_89),
.Y(n_109)
);

NAND4xp25_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_64),
.C(n_63),
.D(n_65),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_79),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_98),
.Y(n_114)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_92),
.B(n_100),
.Y(n_115)
);

CKINVDCx8_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_102),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AO21x2_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_104),
.B(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_103),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_112),
.C(n_110),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_119),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_112),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_132),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_88),
.B1(n_91),
.B2(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_123),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_105),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_132),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

OAI221xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_133),
.B1(n_136),
.B2(n_116),
.C(n_58),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_126),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_124),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_129),
.Y(n_147)
);

NOR2xp67_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_122),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_129),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_128),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_42),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

AOI31xp33_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_126),
.A3(n_128),
.B(n_44),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_44),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_146),
.C(n_61),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_59),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_59),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_165),
.A3(n_164),
.B1(n_159),
.B2(n_85),
.C1(n_161),
.C2(n_150),
.Y(n_168)
);

NOR4xp75_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_9),
.C(n_85),
.D(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_151),
.Y(n_170)
);

NAND4xp75_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_88),
.C(n_83),
.D(n_82),
.Y(n_171)
);

AOI211xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_151),
.B(n_124),
.C(n_122),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_30),
.B1(n_124),
.B2(n_122),
.Y(n_173)
);

NOR2x1p5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_81),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_168),
.B1(n_169),
.B2(n_125),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_54),
.B(n_132),
.C(n_93),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_173),
.Y(n_177)
);

NAND5xp2_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_101),
.C(n_95),
.D(n_109),
.E(n_28),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_178),
.B1(n_11),
.B2(n_94),
.Y(n_180)
);


endmodule