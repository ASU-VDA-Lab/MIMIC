module fake_jpeg_624_n_130 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_14),
.B(n_31),
.C(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_34),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_48),
.B(n_42),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_33),
.B(n_41),
.C(n_34),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_33),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_35),
.C(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_70),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_35),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_16),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_2),
.Y(n_88)
);

OA21x2_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_91),
.B(n_10),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_71),
.B1(n_68),
.B2(n_5),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_17),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_12),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_3),
.B(n_4),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_95),
.B(n_6),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_3),
.B(n_6),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_13),
.C(n_26),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_7),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_9),
.CI(n_10),
.CON(n_108),
.SN(n_108)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_110),
.B1(n_89),
.B2(n_25),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_9),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_20),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_108),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_122),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_119),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_120),
.B1(n_106),
.B2(n_121),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_111),
.B1(n_124),
.B2(n_110),
.Y(n_128)
);

OAI21x1_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_113),
.B(n_115),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_115),
.Y(n_130)
);


endmodule