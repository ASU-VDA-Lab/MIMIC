module fake_netlist_1_9674_n_572 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_572);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_572;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g72 ( .A(n_56), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_37), .Y(n_73) );
INVxp33_ASAP7_75t_SL g74 ( .A(n_62), .Y(n_74) );
INVxp67_ASAP7_75t_L g75 ( .A(n_39), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_58), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_63), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_19), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_36), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_30), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_41), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_68), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_46), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_70), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_4), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_42), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_52), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_29), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_33), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_43), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_44), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_24), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_32), .B(n_53), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_10), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_65), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_1), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_69), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_55), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_50), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_67), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_25), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_51), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_66), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_11), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_110), .Y(n_116) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_73), .A2(n_22), .B(n_64), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_110), .Y(n_119) );
INVx6_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_99), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_105), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_105), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_108), .Y(n_124) );
NOR2xp33_ASAP7_75t_R g125 ( .A(n_85), .B(n_20), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_82), .B(n_0), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
NOR2xp33_ASAP7_75t_R g128 ( .A(n_86), .B(n_23), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_105), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_115), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_78), .Y(n_135) );
INVx2_ASAP7_75t_SL g136 ( .A(n_83), .Y(n_136) );
INVxp67_ASAP7_75t_SL g137 ( .A(n_72), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_100), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_115), .Y(n_139) );
BUFx8_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_73), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_74), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_97), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_97), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_76), .B(n_1), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_97), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_75), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_76), .B(n_2), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_102), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_77), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_102), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_109), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_77), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_79), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_140), .Y(n_158) );
INVx4_ASAP7_75t_SL g159 ( .A(n_120), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_137), .B(n_81), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_152), .B(n_114), .Y(n_163) );
OAI22xp33_ASAP7_75t_L g164 ( .A1(n_116), .A2(n_114), .B1(n_113), .B2(n_112), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_134), .B(n_88), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_151), .B(n_113), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_152), .A2(n_112), .B1(n_98), .B2(n_91), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_120), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_116), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_140), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_117), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_149), .B(n_111), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_155), .B(n_111), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_143), .B(n_79), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_130), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_118), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_144), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_143), .B(n_95), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_118), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_140), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_127), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_132), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_155), .A2(n_95), .B1(n_84), .B2(n_106), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_127), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_120), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_141), .B(n_80), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_156), .B(n_80), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_126), .A2(n_84), .B1(n_92), .B2(n_106), .Y(n_206) );
INVx4_ASAP7_75t_SL g207 ( .A(n_133), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_136), .B(n_92), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_161), .Y(n_211) );
BUFx12f_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
NOR3xp33_ASAP7_75t_SL g213 ( .A(n_164), .B(n_121), .C(n_124), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_162), .B(n_142), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_194), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_166), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_176), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_183), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_208), .Y(n_220) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_187), .B(n_146), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_194), .Y(n_222) );
INVx5_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
OR2x2_ASAP7_75t_SL g225 ( .A(n_168), .B(n_121), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_166), .B(n_142), .Y(n_226) );
NOR2xp33_ASAP7_75t_R g227 ( .A(n_175), .B(n_119), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_174), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_179), .B(n_147), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_208), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_204), .B(n_136), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_208), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_204), .B(n_150), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_158), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_204), .B(n_128), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_168), .B(n_124), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_163), .B(n_123), .Y(n_239) );
OR2x6_ASAP7_75t_L g240 ( .A(n_175), .B(n_93), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_163), .B(n_123), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_163), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_198), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_179), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_180), .B(n_125), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_177), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_184), .B(n_122), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_179), .B(n_129), .Y(n_248) );
NAND2x1p5_ASAP7_75t_L g249 ( .A(n_178), .B(n_122), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_197), .B(n_205), .Y(n_250) );
INVxp67_ASAP7_75t_SL g251 ( .A(n_201), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_182), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_181), .B(n_148), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_169), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_195), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g258 ( .A(n_193), .B(n_3), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_185), .B(n_148), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_195), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_186), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_195), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_190), .B(n_104), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_186), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_191), .B(n_145), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_242), .A2(n_217), .B1(n_248), .B2(n_256), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_236), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_264), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_236), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_251), .B(n_192), .Y(n_270) );
AOI21x1_ASAP7_75t_L g271 ( .A1(n_250), .A2(n_167), .B(n_171), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_224), .B(n_206), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_224), .B(n_159), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_261), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_261), .A2(n_199), .B1(n_203), .B2(n_202), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_220), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_224), .B(n_159), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_219), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_230), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_235), .B(n_159), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_250), .A2(n_177), .B(n_117), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_240), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_233), .B(n_203), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_228), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_247), .A2(n_177), .B(n_117), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_223), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_227), .Y(n_292) );
OR2x6_ASAP7_75t_L g293 ( .A(n_240), .B(n_177), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_239), .B(n_188), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_241), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_212), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_240), .A2(n_188), .B1(n_199), .B2(n_202), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_246), .Y(n_298) );
AOI22xp33_ASAP7_75t_SL g299 ( .A1(n_229), .A2(n_107), .B1(n_90), .B2(n_94), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_240), .B(n_159), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_248), .B(n_157), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_246), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_227), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_212), .Y(n_304) );
CKINVDCx8_ASAP7_75t_R g305 ( .A(n_229), .Y(n_305) );
INVx3_ASAP7_75t_SL g306 ( .A(n_244), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_238), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_223), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_248), .B(n_157), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_229), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_226), .B(n_173), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_246), .Y(n_312) );
AOI22xp33_ASAP7_75t_SL g313 ( .A1(n_292), .A2(n_244), .B1(n_258), .B2(n_238), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_283), .A2(n_218), .B(n_215), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_284), .B(n_239), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_297), .A2(n_263), .B1(n_221), .B2(n_231), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_293), .A2(n_237), .B(n_209), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_280), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_268), .A2(n_253), .B(n_252), .C(n_257), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_294), .B(n_221), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_241), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_307), .A2(n_263), .B1(n_234), .B2(n_214), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_270), .B(n_263), .Y(n_326) );
INVx4_ASAP7_75t_SL g327 ( .A(n_293), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_284), .A2(n_263), .B1(n_225), .B2(n_249), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_287), .B(n_225), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_310), .A2(n_258), .B1(n_255), .B2(n_260), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_284), .B(n_211), .Y(n_331) );
OAI211xp5_ASAP7_75t_SL g332 ( .A1(n_299), .A2(n_213), .B(n_245), .C(n_101), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_277), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_281), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_310), .A2(n_262), .B1(n_260), .B2(n_249), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_262), .B1(n_210), .B2(n_259), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_288), .A2(n_117), .B(n_265), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_322), .A2(n_266), .B1(n_274), .B2(n_303), .C(n_292), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_322), .A2(n_303), .B1(n_275), .B2(n_296), .C(n_311), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_313), .A2(n_272), .B1(n_306), .B2(n_284), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_338), .B(n_272), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_340), .A2(n_312), .B(n_302), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_338), .B(n_272), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_332), .A2(n_293), .B1(n_304), .B2(n_300), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_325), .A2(n_254), .B1(n_309), .B2(n_301), .C(n_103), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_326), .B(n_262), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_321), .B(n_305), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_326), .A2(n_293), .B1(n_300), .B2(n_282), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_321), .A2(n_300), .B1(n_133), .B2(n_290), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_329), .A2(n_282), .B1(n_308), .B2(n_289), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_333), .B(n_305), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_329), .A2(n_282), .B1(n_308), .B2(n_290), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_314), .A2(n_271), .B(n_302), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_333), .B(n_290), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_316), .A2(n_279), .B1(n_273), .B2(n_223), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_316), .A2(n_328), .B1(n_335), .B2(n_337), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_318), .B(n_335), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_330), .A2(n_279), .B1(n_273), .B2(n_223), .Y(n_365) );
OAI33xp33_ASAP7_75t_L g366 ( .A1(n_363), .A2(n_93), .A3(n_101), .B1(n_103), .B2(n_104), .B3(n_337), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_363), .A2(n_315), .B1(n_339), .B2(n_336), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_345), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_345), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_341), .A2(n_315), .B1(n_334), .B2(n_323), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_350), .B(n_315), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_345), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_350), .B(n_327), .Y(n_374) );
OAI31xp33_ASAP7_75t_L g375 ( .A1(n_344), .A2(n_320), .A3(n_334), .B(n_273), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_317), .B(n_340), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_341), .A2(n_331), .B1(n_327), .B2(n_279), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_362), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_361), .A2(n_324), .B1(n_331), .B2(n_269), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_362), .B(n_327), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_362), .B(n_327), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
NOR2x1_ASAP7_75t_SL g384 ( .A(n_358), .B(n_269), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_346), .B(n_331), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_346), .B(n_109), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_109), .B(n_165), .Y(n_389) );
NOR3xp33_ASAP7_75t_SL g390 ( .A(n_342), .B(n_96), .C(n_165), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
OA222x2_ASAP7_75t_L g392 ( .A1(n_356), .A2(n_96), .B1(n_5), .B2(n_6), .C1(n_7), .C2(n_8), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_353), .B(n_198), .C(n_200), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_390), .B(n_364), .C(n_347), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_368), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_366), .A2(n_387), .B1(n_370), .B2(n_383), .C(n_356), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_388), .B(n_358), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_382), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_378), .B(n_354), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_375), .B(n_354), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_388), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_376), .A2(n_359), .B(n_349), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_377), .A2(n_351), .B1(n_343), .B2(n_353), .Y(n_405) );
OAI33xp33_ASAP7_75t_L g406 ( .A1(n_392), .A2(n_349), .A3(n_171), .B1(n_172), .B2(n_167), .B3(n_200), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_383), .B(n_351), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_378), .B(n_354), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_382), .B(n_354), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_382), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_368), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_371), .B(n_359), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_390), .A2(n_352), .B1(n_355), .B2(n_357), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_391), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_391), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_374), .B(n_359), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_380), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_382), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_369), .B(n_359), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_367), .A2(n_365), .B1(n_196), .B2(n_172), .C(n_170), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_386), .B(n_3), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_369), .Y(n_427) );
AO31x2_ASAP7_75t_L g428 ( .A1(n_379), .A2(n_170), .A3(n_298), .B(n_291), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_373), .B(n_5), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
NAND2x1_ASAP7_75t_SL g431 ( .A(n_373), .B(n_312), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_381), .B(n_6), .Y(n_433) );
AOI21x1_ASAP7_75t_L g434 ( .A1(n_429), .A2(n_385), .B(n_381), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_394), .B(n_415), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_427), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_414), .B(n_385), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
BUFx12f_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_417), .B(n_392), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_427), .Y(n_441) );
OAI33xp33_ASAP7_75t_L g442 ( .A1(n_426), .A2(n_379), .A3(n_8), .B1(n_9), .B2(n_11), .B3(n_12), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_420), .B(n_385), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_416), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_408), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_421), .B(n_375), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_427), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_406), .B(n_366), .Y(n_449) );
NAND2xp33_ASAP7_75t_SL g450 ( .A(n_400), .B(n_376), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_418), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_395), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_429), .B(n_384), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_419), .B(n_389), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_422), .B(n_393), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_425), .B(n_7), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_403), .B(n_9), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_397), .B(n_12), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_433), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_433), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_407), .B(n_13), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_396), .B(n_13), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_395), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_412), .Y(n_464) );
INVx5_ASAP7_75t_L g465 ( .A(n_400), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_422), .B(n_393), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_431), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_424), .B(n_173), .C(n_243), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_419), .B(n_14), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_432), .B(n_15), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_399), .B(n_15), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_422), .B(n_276), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_399), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_413), .B(n_17), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_436), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_470), .B(n_423), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_465), .B(n_411), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_443), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_465), .A2(n_411), .B1(n_402), .B2(n_409), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_468), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_440), .B(n_402), .Y(n_482) );
AO22x1_ASAP7_75t_L g483 ( .A1(n_465), .A2(n_410), .B1(n_408), .B2(n_401), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_435), .B(n_404), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_451), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_441), .Y(n_488) );
NAND4xp25_ASAP7_75t_SL g489 ( .A(n_458), .B(n_405), .C(n_410), .D(n_431), .Y(n_489) );
AOI21xp33_ASAP7_75t_SL g490 ( .A1(n_457), .A2(n_404), .B(n_27), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_438), .B(n_446), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_442), .B(n_18), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_465), .A2(n_428), .B1(n_278), .B2(n_269), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_428), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_449), .A2(n_428), .B(n_222), .Y(n_496) );
NAND2xp33_ASAP7_75t_L g497 ( .A(n_471), .B(n_276), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_453), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_437), .B(n_428), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_459), .B(n_28), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_460), .B(n_31), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_449), .A2(n_269), .B1(n_276), .B2(n_267), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_447), .A2(n_207), .B1(n_267), .B2(n_276), .Y(n_504) );
OAI222xp33_ASAP7_75t_L g505 ( .A1(n_464), .A2(n_35), .B1(n_38), .B2(n_45), .C1(n_47), .C2(n_49), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_472), .B(n_269), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_444), .B(n_54), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_475), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g509 ( .A1(n_462), .A2(n_57), .B(n_59), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_445), .B(n_438), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_474), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_454), .B(n_60), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_499), .B(n_446), .Y(n_513) );
XOR2xp5_ASAP7_75t_L g514 ( .A(n_489), .B(n_461), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_484), .B(n_463), .Y(n_515) );
NOR3xp33_ASAP7_75t_SL g516 ( .A(n_482), .B(n_450), .C(n_456), .Y(n_516) );
INVxp33_ASAP7_75t_L g517 ( .A(n_491), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_491), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_485), .A2(n_455), .B(n_466), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g522 ( .A1(n_508), .A2(n_439), .B1(n_466), .B2(n_455), .C1(n_448), .C2(n_467), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_476), .Y(n_523) );
CKINVDCx20_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_510), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_481), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_480), .B(n_439), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_492), .A2(n_500), .B1(n_487), .B2(n_480), .Y(n_528) );
AOI211x1_ASAP7_75t_L g529 ( .A1(n_478), .A2(n_434), .B(n_466), .C(n_455), .Y(n_529) );
BUFx4f_ASAP7_75t_SL g530 ( .A(n_478), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_511), .Y(n_531) );
XOR2xp5_ASAP7_75t_L g532 ( .A(n_477), .B(n_473), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_486), .B(n_467), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_486), .B(n_469), .Y(n_534) );
AND3x2_ASAP7_75t_L g535 ( .A(n_492), .B(n_473), .C(n_61), .Y(n_535) );
INVx6_ASAP7_75t_L g536 ( .A(n_495), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_527), .A2(n_497), .B(n_505), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_516), .A2(n_490), .B(n_488), .C(n_496), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g539 ( .A1(n_529), .A2(n_509), .B(n_488), .C(n_512), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_523), .Y(n_540) );
AND2x2_ASAP7_75t_SL g541 ( .A(n_524), .B(n_503), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_530), .B(n_494), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_528), .B(n_493), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_519), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_533), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_514), .A2(n_502), .B1(n_501), .B2(n_506), .Y(n_546) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_536), .A2(n_504), .B1(n_507), .B2(n_498), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_534), .A2(n_216), .B(n_71), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_525), .Y(n_549) );
XNOR2xp5_ASAP7_75t_L g550 ( .A(n_532), .B(n_207), .Y(n_550) );
NOR2xp33_ASAP7_75t_R g551 ( .A(n_541), .B(n_535), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_540), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_541), .B(n_522), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_537), .A2(n_549), .B1(n_542), .B2(n_544), .Y(n_554) );
AOI221x1_ASAP7_75t_L g555 ( .A1(n_543), .A2(n_534), .B1(n_533), .B2(n_521), .C(n_515), .Y(n_555) );
NOR2xp33_ASAP7_75t_R g556 ( .A(n_550), .B(n_513), .Y(n_556) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_538), .B(n_518), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_539), .B(n_548), .C(n_547), .Y(n_558) );
OAI211xp5_ASAP7_75t_SL g559 ( .A1(n_546), .A2(n_526), .B(n_520), .C(n_531), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_547), .A2(n_207), .B1(n_545), .B2(n_543), .C(n_482), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_537), .A2(n_530), .B1(n_517), .B2(n_549), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_556), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_552), .Y(n_563) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_557), .B(n_553), .Y(n_564) );
CKINVDCx16_ASAP7_75t_R g565 ( .A(n_551), .Y(n_565) );
OR4x2_ASAP7_75t_L g566 ( .A(n_565), .B(n_561), .C(n_554), .D(n_555), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_563), .Y(n_567) );
NOR2x1p5_ASAP7_75t_L g568 ( .A(n_567), .B(n_562), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_566), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_568), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_570), .A2(n_569), .B1(n_564), .B2(n_558), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_571), .A2(n_566), .B1(n_564), .B2(n_559), .C(n_560), .Y(n_572) );
endmodule