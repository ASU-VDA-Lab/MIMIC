module fake_jpeg_1804_n_227 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_8),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_16),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_0),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_86),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_22),
.B1(n_51),
.B2(n_47),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_57),
.B1(n_79),
.B2(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_80),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_95),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_65),
.B(n_71),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_67),
.B1(n_61),
.B2(n_72),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_74),
.B1(n_73),
.B2(n_72),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_75),
.C(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_106),
.Y(n_128)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_67),
.Y(n_133)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_78),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_89),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_120),
.Y(n_131)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_94),
.B1(n_105),
.B2(n_107),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_90),
.C(n_96),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_77),
.C(n_62),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_78),
.B1(n_61),
.B2(n_67),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_77),
.B1(n_68),
.B2(n_62),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_126),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_82),
.B1(n_57),
.B2(n_76),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_115),
.B1(n_109),
.B2(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_0),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_78),
.B1(n_75),
.B2(n_76),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_1),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_146),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_163),
.B1(n_4),
.B2(n_7),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_160),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_154),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_68),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_52),
.C(n_40),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_158),
.C(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_1),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx24_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_128),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_62),
.B1(n_24),
.B2(n_25),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_162),
.B(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_2),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_2),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_164),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_21),
.B1(n_44),
.B2(n_43),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_3),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_167),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_179),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_135),
.B(n_7),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_178),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_26),
.B(n_42),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_27),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_159),
.B1(n_12),
.B2(n_13),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_38),
.B(n_35),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_153),
.B(n_151),
.C(n_147),
.D(n_162),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_178),
.B(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_198),
.B1(n_187),
.B2(n_170),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_203),
.C(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_181),
.C(n_180),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_175),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_175),
.C(n_186),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_199),
.B(n_168),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_199),
.B1(n_183),
.B2(n_195),
.Y(n_211)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_212),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_185),
.B1(n_16),
.B2(n_17),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_217),
.B1(n_216),
.B2(n_212),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_215),
.A2(n_213),
.B1(n_202),
.B2(n_204),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_218),
.A3(n_217),
.B1(n_209),
.B2(n_214),
.C1(n_28),
.C2(n_30),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_31),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_32),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_15),
.B(n_17),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_18),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_19),
.Y(n_227)
);


endmodule