module fake_jpeg_12587_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_69),
.Y(n_125)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_64),
.B(n_75),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_67),
.B(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_83),
.B(n_96),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_85),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_89),
.Y(n_166)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_91),
.B(n_106),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_102),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_39),
.B(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_97),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_40),
.A2(n_1),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_98),
.B(n_1),
.Y(n_158)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_33),
.Y(n_138)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_44),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_105),
.B(n_52),
.Y(n_154)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g235 ( 
.A(n_110),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_66),
.A2(n_28),
.B1(n_43),
.B2(n_41),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_111),
.A2(n_171),
.B1(n_51),
.B2(n_35),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_138),
.Y(n_174)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_31),
.B1(n_50),
.B2(n_47),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_139),
.A2(n_168),
.B1(n_47),
.B2(n_41),
.Y(n_229)
);

BUFx16f_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_69),
.A2(n_50),
.B(n_31),
.C(n_47),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_142),
.A2(n_63),
.B(n_50),
.C(n_31),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_44),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_155),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_154),
.B(n_158),
.C(n_3),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_29),
.Y(n_155)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_77),
.B(n_29),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_65),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_88),
.A2(n_51),
.B1(n_43),
.B2(n_38),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_104),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_72),
.A2(n_43),
.B1(n_38),
.B2(n_41),
.Y(n_171)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_177),
.B(n_180),
.Y(n_284)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_126),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_112),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_188),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_42),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_182),
.B(n_185),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_108),
.C(n_101),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_198),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_37),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_53),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_190),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_70),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_189),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_53),
.Y(n_190)
);

CKINVDCx12_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_191),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_137),
.B(n_24),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_195),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_197),
.A2(n_207),
.B1(n_115),
.B2(n_152),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_142),
.B(n_59),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_37),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_146),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_42),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_203),
.B(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_24),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_61),
.B1(n_62),
.B2(n_99),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_131),
.B(n_87),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_135),
.Y(n_280)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_166),
.A2(n_35),
.B1(n_36),
.B2(n_95),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_211),
.A2(n_213),
.B1(n_226),
.B2(n_233),
.Y(n_274)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_SL g217 ( 
.A(n_164),
.B(n_50),
.Y(n_217)
);

NAND2x1p5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_134),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_107),
.B1(n_100),
.B2(n_86),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_218),
.A2(n_221),
.B1(n_223),
.B2(n_150),
.Y(n_275)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_220),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_139),
.A2(n_80),
.B1(n_78),
.B2(n_74),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_36),
.Y(n_222)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_162),
.A2(n_50),
.B1(n_47),
.B2(n_31),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_113),
.B(n_50),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_228),
.A2(n_173),
.B1(n_172),
.B2(n_157),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_234),
.B1(n_116),
.B2(n_169),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_133),
.B(n_4),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_236),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_114),
.Y(n_231)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_132),
.A2(n_38),
.B1(n_47),
.B2(n_33),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_232),
.A2(n_33),
.B1(n_122),
.B2(n_123),
.Y(n_288)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_162),
.A2(n_47),
.B1(n_33),
.B2(n_46),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_133),
.B(n_4),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_240),
.A2(n_242),
.B1(n_245),
.B2(n_248),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_181),
.A2(n_141),
.B1(n_159),
.B2(n_153),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_132),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_247),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_150),
.B1(n_124),
.B2(n_153),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_174),
.B(n_198),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_188),
.B1(n_223),
.B2(n_197),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_251),
.A2(n_199),
.B(n_205),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_196),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_263),
.Y(n_302)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_135),
.A3(n_117),
.B1(n_119),
.B2(n_145),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_260),
.A2(n_233),
.B(n_207),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_183),
.B(n_118),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_273),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_143),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_277),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_220),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_176),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_178),
.B(n_124),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_209),
.C(n_202),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_287),
.B1(n_292),
.B2(n_231),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_172),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_188),
.B(n_157),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_215),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_184),
.A2(n_147),
.B1(n_122),
.B2(n_173),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_291),
.B1(n_189),
.B2(n_205),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_207),
.A2(n_145),
.B1(n_123),
.B2(n_119),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_232),
.A2(n_33),
.B1(n_123),
.B2(n_119),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_249),
.B(n_257),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_294),
.B(n_298),
.C(n_304),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_307),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_249),
.B(n_284),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_299),
.A2(n_323),
.B1(n_326),
.B2(n_237),
.Y(n_358)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_300),
.Y(n_373)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_301),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_243),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_305),
.A2(n_313),
.B(n_12),
.Y(n_381)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_306),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_258),
.B(n_175),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_309),
.B(n_316),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_235),
.C(n_6),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_324),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_251),
.A2(n_199),
.B(n_225),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_277),
.B(n_244),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_247),
.A2(n_216),
.B1(n_194),
.B2(n_208),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_241),
.B(n_251),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_315),
.B(n_318),
.C(n_320),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_241),
.B(n_235),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_319),
.B(n_322),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_266),
.B(n_235),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_285),
.B(n_194),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_281),
.A2(n_216),
.B1(n_187),
.B2(n_210),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_252),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_176),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_337),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_281),
.A2(n_187),
.B1(n_219),
.B2(n_212),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_329),
.Y(n_356)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_239),
.B(n_214),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_239),
.B(n_206),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_335),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_334),
.Y(n_372)
);

AO22x1_ASAP7_75t_SL g335 ( 
.A1(n_277),
.A2(n_201),
.B1(n_163),
.B2(n_7),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_268),
.B(n_176),
.C(n_6),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_268),
.C(n_280),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_18),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_250),
.B(n_4),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_341),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_8),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_240),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_267),
.B1(n_261),
.B2(n_289),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_338),
.A2(n_277),
.B1(n_288),
.B2(n_268),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_347),
.A2(n_357),
.B1(n_313),
.B2(n_379),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_297),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_355),
.C(n_360),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_311),
.A2(n_245),
.B1(n_273),
.B2(n_274),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_354),
.A2(n_362),
.B1(n_336),
.B2(n_327),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_286),
.C(n_250),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_357),
.A2(n_371),
.B(n_335),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_381),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_272),
.C(n_253),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_299),
.A2(n_289),
.B1(n_261),
.B2(n_256),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_305),
.A2(n_244),
.B(n_290),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_363),
.A2(n_386),
.B(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_376),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_265),
.B1(n_262),
.B2(n_254),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_365),
.A2(n_375),
.B1(n_380),
.B2(n_301),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_290),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_378),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_237),
.B(n_265),
.Y(n_371)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_18),
.B1(n_9),
.B2(n_11),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_8),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_303),
.B(n_8),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_293),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_312),
.A2(n_12),
.B(n_13),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_350),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_394),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_417),
.B1(n_421),
.B2(n_425),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_353),
.B(n_302),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_390),
.Y(n_437)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_391),
.B(n_420),
.C(n_403),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_393),
.A2(n_371),
.B1(n_384),
.B2(n_351),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_374),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_314),
.Y(n_396)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

NOR2x1_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_315),
.Y(n_397)
);

AO21x1_ASAP7_75t_L g449 ( 
.A1(n_397),
.A2(n_424),
.B(n_382),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_398),
.A2(n_423),
.B(n_424),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_372),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_415),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_331),
.Y(n_401)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_404),
.A2(n_405),
.B1(n_348),
.B2(n_363),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_354),
.A2(n_320),
.B1(n_329),
.B2(n_318),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_321),
.Y(n_406)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_406),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_369),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_408),
.B(n_351),
.Y(n_456)
);

INVx13_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_409),
.Y(n_454)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_304),
.Y(n_412)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_412),
.Y(n_447)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

BUFx12_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g457 ( 
.A(n_414),
.Y(n_457)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_359),
.B(n_342),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_418),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_368),
.A2(n_335),
.B1(n_337),
.B2(n_306),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_361),
.B(n_334),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_317),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_419),
.B(n_366),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_355),
.B(n_300),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_365),
.A2(n_328),
.B1(n_330),
.B2(n_332),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_422),
.A2(n_386),
.B(n_385),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_346),
.A2(n_333),
.B(n_296),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_346),
.A2(n_341),
.B(n_13),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_375),
.A2(n_341),
.B1(n_14),
.B2(n_15),
.Y(n_425)
);

XNOR2x1_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_392),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_416),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_432),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_390),
.Y(n_436)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_369),
.Y(n_438)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_352),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_459),
.C(n_399),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_394),
.B(n_383),
.Y(n_440)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_442),
.A2(n_445),
.B(n_446),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_398),
.A2(n_361),
.B(n_371),
.Y(n_446)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_449),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_422),
.A2(n_373),
.B(n_384),
.Y(n_451)
);

XNOR2x2_ASAP7_75t_SL g481 ( 
.A(n_451),
.B(n_423),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_458),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_456),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_389),
.A2(n_345),
.B1(n_378),
.B2(n_344),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_345),
.C(n_344),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_473),
.C(n_475),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_436),
.B(n_397),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_461),
.B(n_471),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_440),
.B(n_396),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_465),
.B(n_476),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_399),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_427),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_SL g471 ( 
.A(n_429),
.B(n_397),
.C(n_437),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_472),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_405),
.C(n_404),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_481),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_406),
.C(n_403),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_433),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_426),
.B(n_401),
.C(n_412),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_483),
.C(n_484),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_430),
.B(n_428),
.Y(n_479)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_479),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_447),
.B(n_392),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_487),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_392),
.C(n_411),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_410),
.C(n_413),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_447),
.A2(n_417),
.B1(n_441),
.B2(n_445),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_486),
.A2(n_452),
.B1(n_444),
.B2(n_443),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_427),
.B(n_418),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_463),
.A2(n_429),
.B1(n_441),
.B2(n_431),
.Y(n_491)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_480),
.A2(n_449),
.B(n_446),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_493),
.A2(n_488),
.B(n_470),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_502),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_431),
.B1(n_451),
.B2(n_393),
.Y(n_495)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_495),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_467),
.A2(n_453),
.B1(n_442),
.B2(n_395),
.Y(n_497)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_497),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_468),
.A2(n_453),
.B1(n_395),
.B2(n_421),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_503),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_460),
.B(n_438),
.C(n_449),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_501),
.C(n_504),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_434),
.C(n_452),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_433),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_434),
.C(n_444),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_457),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_505),
.B(n_512),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_479),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_469),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_443),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_509),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_415),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_464),
.B(n_380),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_511),
.A2(n_488),
.B(n_485),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_515),
.B(n_519),
.Y(n_542)
);

XNOR2x2_ASAP7_75t_SL g516 ( 
.A(n_489),
.B(n_482),
.Y(n_516)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_516),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_522),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_510),
.A2(n_486),
.B(n_470),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_520),
.A2(n_527),
.B1(n_454),
.B2(n_364),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_483),
.C(n_487),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_475),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_526),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_497),
.Y(n_526)
);

OA21x2_ASAP7_75t_SL g527 ( 
.A1(n_506),
.A2(n_462),
.B(n_471),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_501),
.B(n_484),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_531),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_491),
.B(n_462),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_528),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_518),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_530),
.A2(n_496),
.B1(n_508),
.B2(n_502),
.Y(n_534)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_490),
.C(n_498),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_538),
.C(n_539),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_520),
.A2(n_499),
.B1(n_495),
.B2(n_498),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_537),
.A2(n_546),
.B1(n_514),
.B2(n_524),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_490),
.C(n_509),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_494),
.C(n_492),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_492),
.C(n_489),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_541),
.C(n_543),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_481),
.C(n_472),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_513),
.B(n_402),
.C(n_454),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_544),
.Y(n_558)
);

O2A1O1Ixp5_ASAP7_75t_L g546 ( 
.A1(n_515),
.A2(n_414),
.B(n_409),
.C(n_425),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_549),
.B(n_539),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_545),
.A2(n_514),
.B1(n_524),
.B2(n_523),
.Y(n_550)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_550),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_531),
.Y(n_551)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_551),
.A2(n_557),
.B(n_533),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_536),
.B(n_530),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_554),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_547),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_517),
.Y(n_564)
);

HAxp5_ASAP7_75t_SL g557 ( 
.A(n_532),
.B(n_516),
.CON(n_557),
.SN(n_557)
);

AOI221xp5_ASAP7_75t_L g559 ( 
.A1(n_535),
.A2(n_523),
.B1(n_517),
.B2(n_516),
.C(n_414),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_559),
.A2(n_541),
.B(n_543),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_561),
.B(n_555),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_553),
.A2(n_538),
.B(n_540),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_562),
.B(n_564),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_565),
.B(n_553),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_566),
.A2(n_548),
.B1(n_554),
.B2(n_558),
.Y(n_568)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_567),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_568),
.A2(n_560),
.B(n_563),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_569),
.B(n_555),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_571),
.A2(n_572),
.B(n_560),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_574),
.Y(n_576)
);

AOI322xp5_ASAP7_75t_L g575 ( 
.A1(n_573),
.A2(n_550),
.A3(n_570),
.B1(n_551),
.B2(n_549),
.C1(n_414),
.C2(n_557),
.Y(n_575)
);

AOI322xp5_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_575),
.A3(n_367),
.B1(n_341),
.B2(n_377),
.C1(n_15),
.C2(n_14),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_SL g578 ( 
.A1(n_577),
.A2(n_12),
.B(n_14),
.C(n_16),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_377),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_16),
.B(n_574),
.Y(n_580)
);


endmodule