module fake_jpeg_13522_n_189 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_26),
.B1(n_32),
.B2(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_66)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_52),
.Y(n_54)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_58),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_77),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_73),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_21),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_75),
.B(n_62),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_50),
.B1(n_48),
.B2(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_23),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_12),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_96),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_43),
.B(n_1),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_91),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_97),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_0),
.B(n_2),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_101),
.B1(n_65),
.B2(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_7),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_11),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_74),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_11),
.B1(n_70),
.B2(n_72),
.Y(n_101)
);

AO22x2_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_80),
.B1(n_74),
.B2(n_72),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_101),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_63),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_114),
.C(n_121),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_102),
.B1(n_93),
.B2(n_91),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_119),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_102),
.B(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_87),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_95),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_133),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_98),
.C(n_86),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_126),
.C(n_142),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_111),
.B1(n_118),
.B2(n_106),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_142),
.B(n_130),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_88),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_99),
.B1(n_104),
.B2(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_106),
.B1(n_113),
.B2(n_111),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_118),
.B1(n_106),
.B2(n_123),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_116),
.B(n_109),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_155),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_109),
.A3(n_116),
.B1(n_124),
.B2(n_125),
.C1(n_127),
.C2(n_136),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_143),
.C(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_131),
.C(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_163),
.C(n_164),
.Y(n_170)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_166),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_156),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_139),
.C(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_151),
.B1(n_152),
.B2(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_159),
.C(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_177),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_158),
.C(n_164),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_155),
.B(n_166),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_157),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_157),
.C(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_171),
.C(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_144),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_183),
.A2(n_179),
.B1(n_167),
.B2(n_147),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_153),
.B(n_187),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_186),
.Y(n_189)
);


endmodule