module real_jpeg_17458_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_358),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_0),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_25),
.Y(n_24)
);

AND2x4_ASAP7_75t_SL g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_45),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_59),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_4),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_4),
.B(n_281),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_5),
.Y(n_142)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_6),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_6),
.B(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_6),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_6),
.B(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_7),
.Y(n_197)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_8),
.Y(n_359)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_9),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_9),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_9),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_9),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_9),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_175),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_173),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_149),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_19),
.B(n_149),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_88),
.C(n_113),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_20),
.B(n_89),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_21),
.B(n_61),
.C(n_71),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_46),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_22),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_23),
.A2(n_36),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.Y(n_23)
);

NAND2x1p5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_24),
.A2(n_63),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_24),
.B(n_92),
.C(n_98),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_24),
.A2(n_63),
.B1(n_140),
.B2(n_218),
.Y(n_263)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_40),
.B(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_31),
.C(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_28),
.A2(n_40),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_28),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_28),
.A2(n_118),
.B1(n_214),
.B2(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_30),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_30),
.B(n_31),
.C(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_37),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_31),
.A2(n_37),
.B1(n_248),
.B2(n_252),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_36),
.A2(n_200),
.B(n_206),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_37),
.B(n_74),
.C(n_105),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_38),
.B(n_46),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_39),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_40),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_40),
.A2(n_119),
.B1(n_201),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_40),
.A2(n_78),
.B1(n_119),
.B2(n_133),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_40),
.B(n_78),
.C(n_261),
.Y(n_312)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_48),
.A2(n_49),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_48),
.A2(n_49),
.B1(n_98),
.B2(n_99),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_51),
.C(n_112),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_49),
.A2(n_99),
.B(n_194),
.C(n_227),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_50),
.Y(n_190)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_56),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_56),
.B(n_132),
.C(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_56),
.A2(n_82),
.B1(n_112),
.B2(n_132),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_56),
.A2(n_112),
.B1(n_248),
.B2(n_252),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_93),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_57),
.B(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_62),
.B(n_65),
.C(n_67),
.Y(n_162)
);

NOR2x1_ASAP7_75t_R g200 ( 
.A(n_63),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_65),
.A2(n_70),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_65),
.A2(n_70),
.B1(n_171),
.B2(n_172),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_65),
.B(n_99),
.C(n_126),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_72),
.C(n_85),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_66),
.A2(n_67),
.B1(n_143),
.B2(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_135),
.C(n_143),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_67),
.B(n_85),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_67),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_67),
.B(n_74),
.C(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_72),
.A2(n_73),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.C(n_82),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_74),
.A2(n_104),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_78),
.A2(n_82),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_121),
.B(n_129),
.Y(n_120)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_82),
.B(n_122),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_85),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_136),
.C(n_140),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_90),
.B(n_101),
.C(n_111),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_92),
.A2(n_280),
.B(n_286),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_92),
.B(n_280),
.Y(n_286)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_94),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_98),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_98),
.B(n_234),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_112),
.B(n_252),
.C(n_297),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_113),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_134),
.C(n_145),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_114),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_130),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_120),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_122),
.A2(n_123),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_126),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_125),
.A2(n_126),
.B1(n_206),
.B2(n_208),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_125),
.A2(n_126),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_126),
.A2(n_206),
.B(n_225),
.C(n_227),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_126),
.B(n_206),
.Y(n_227)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2x2_ASAP7_75t_L g342 ( 
.A(n_130),
.B(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_134),
.A2(n_145),
.B1(n_146),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_134),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_135),
.B(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_136),
.A2(n_140),
.B1(n_218),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_136),
.Y(n_309)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_140),
.Y(n_218)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_143),
.Y(n_328)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_164),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_163),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_315),
.A3(n_345),
.B1(n_351),
.B2(n_356),
.C(n_357),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_290),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_265),
.B(n_289),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_242),
.B(n_264),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_222),
.B(n_241),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_209),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_209),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_198),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_191),
.B2(n_192),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_185),
.B(n_192),
.C(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_189),
.A2(n_261),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_194),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_193),
.A2(n_194),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_233),
.B(n_235),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_219),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_219),
.B1(n_220),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_214),
.B(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_240),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_237),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_236),
.B(n_239),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_244),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_253),
.C(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_259),
.C(n_263),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_288),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_288),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_269),
.C(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_273),
.C(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_287),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_279),
.C(n_287),
.Y(n_314)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_292),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_305),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_306),
.C(n_314),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_299),
.C(n_303),
.Y(n_341)
);

XNOR2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_314),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_312),
.C(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_333),
.Y(n_315)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_316),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_331),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_331),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.C(n_329),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_329),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_325),
.B1(n_326),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

AOI31xp67_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_346),
.A3(n_352),
.B(n_355),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_336),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.C(n_342),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_337),
.A2(n_338),
.B1(n_342),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_350),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);


endmodule