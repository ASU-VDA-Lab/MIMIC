module fake_jpeg_9180_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_31),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_54),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_23),
.B1(n_35),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_34),
.B1(n_39),
.B2(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_35),
.B1(n_23),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_26),
.B1(n_31),
.B2(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_25),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_40),
.C(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_75),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_18),
.B1(n_32),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_89),
.B1(n_95),
.B2(n_106),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_46),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_18),
.B1(n_34),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_46),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_80),
.Y(n_134)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_87),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_18),
.B1(n_34),
.B2(n_24),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_86),
.B1(n_93),
.B2(n_97),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_66),
.B1(n_27),
.B2(n_29),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_19),
.B1(n_22),
.B2(n_10),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_24),
.B1(n_39),
.B2(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_42),
.B1(n_46),
.B2(n_39),
.Y(n_89)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_98),
.B1(n_105),
.B2(n_108),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_36),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_36),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_58),
.C(n_55),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_41),
.B1(n_36),
.B2(n_42),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_42),
.B1(n_41),
.B2(n_21),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_40),
.B(n_33),
.C(n_30),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_107),
.B(n_22),
.C(n_19),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_42),
.B1(n_33),
.B2(n_30),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_49),
.A2(n_27),
.B1(n_43),
.B2(n_45),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_28),
.B(n_27),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_113),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_63),
.B1(n_13),
.B2(n_14),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_92),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_108),
.B(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_29),
.B1(n_22),
.B2(n_17),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_45),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_45),
.C(n_43),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_135),
.C(n_100),
.Y(n_158)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_131),
.B1(n_102),
.B2(n_82),
.Y(n_166)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_45),
.C(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_45),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_140),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_84),
.B1(n_73),
.B2(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_147),
.B1(n_150),
.B2(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_149),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_74),
.B1(n_73),
.B2(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_130),
.B1(n_120),
.B2(n_132),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_71),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_75),
.B1(n_97),
.B2(n_93),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_167),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_113),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_100),
.B1(n_103),
.B2(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_120),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_101),
.B1(n_81),
.B2(n_99),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_81),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_99),
.B1(n_106),
.B2(n_19),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_58),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_135),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_180),
.C(n_190),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_129),
.B(n_123),
.C(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_174),
.Y(n_227)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_126),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_124),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_120),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_187),
.A2(n_197),
.B(n_203),
.Y(n_212)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_115),
.B(n_1),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_192),
.A2(n_196),
.B(n_169),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_116),
.B1(n_122),
.B2(n_111),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_203),
.B1(n_172),
.B2(n_187),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_55),
.B(n_125),
.Y(n_196)
);

CKINVDCx11_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_145),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_148),
.B(n_161),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_217),
.B(n_157),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_224),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_171),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_221),
.C(n_228),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_0),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_141),
.B(n_140),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_163),
.B1(n_161),
.B2(n_164),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_204),
.B1(n_102),
.B2(n_82),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_153),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_169),
.B(n_1),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_229),
.B(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_191),
.C(n_186),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_182),
.B(n_10),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_8),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.C(n_9),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_157),
.C(n_160),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_254),
.C(n_253),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_179),
.B1(n_173),
.B2(n_192),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_246),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_207),
.B1(n_220),
.B2(n_11),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_174),
.B1(n_204),
.B2(n_175),
.Y(n_238)
);

AOI321xp33_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_222),
.A3(n_229),
.B1(n_212),
.B2(n_205),
.C(n_208),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_242),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_211),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_228),
.C(n_221),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_9),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_9),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_253),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_15),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_1),
.C(n_2),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_10),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_11),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_14),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_264),
.C(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_244),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_270),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_260),
.A2(n_251),
.B(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_206),
.C(n_224),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_233),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_13),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_235),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_246),
.B1(n_249),
.B2(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_207),
.C(n_4),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_277),
.B(n_280),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_250),
.B1(n_239),
.B2(n_252),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_3),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_288),
.B(n_260),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_272),
.B(n_258),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_12),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_12),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_276),
.C(n_257),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_262),
.C(n_263),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_300),
.C(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_285),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_262),
.C(n_263),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_267),
.C(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_305),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_280),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_289),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_290),
.B1(n_299),
.B2(n_300),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_4),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_315),
.B1(n_4),
.B2(n_5),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_4),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_296),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_299),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_309),
.B(n_313),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_294),
.C(n_6),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_316),
.B(n_319),
.Y(n_325)
);

NAND4xp25_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_323),
.C(n_322),
.D(n_320),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_318),
.B(n_5),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_327),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

AO22x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_328),
.B1(n_326),
.B2(n_7),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_5),
.Y(n_332)
);


endmodule