module fake_netlist_5_268_n_2451 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2451);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2451;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_907;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1463;
wire n_1002;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_1412;
wire n_822;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_2243;
wire n_1684;
wire n_921;
wire n_996;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2377;
wire n_2080;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_2431;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_703;
wire n_1115;
wire n_980;
wire n_698;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_376),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_100),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_73),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_124),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_36),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_244),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_207),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_221),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_505),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_218),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_160),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_540),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_320),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_167),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_199),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_503),
.B(n_455),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_43),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_15),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_439),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_262),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_581),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_377),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_530),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_391),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_225),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_473),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_120),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_173),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_549),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_558),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_594),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_81),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_222),
.B(n_245),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_313),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_440),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_526),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_231),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_385),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_364),
.Y(n_650)
);

CKINVDCx16_ASAP7_75t_R g651 ( 
.A(n_392),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_600),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_186),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_198),
.Y(n_654)
);

BUFx5_ASAP7_75t_L g655 ( 
.A(n_309),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_9),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_591),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_446),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_575),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_534),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_249),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_429),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_579),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_383),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_283),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_137),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_199),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_573),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_117),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_205),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_196),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_590),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_272),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_48),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_583),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_332),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_306),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_269),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_460),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_545),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_229),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_130),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_487),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_246),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_92),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_340),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_20),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_431),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_402),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_544),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_483),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_65),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_177),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_360),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_41),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_50),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_35),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_116),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_48),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_492),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_256),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_496),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_77),
.Y(n_706)
);

CKINVDCx14_ASAP7_75t_R g707 ( 
.A(n_224),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_475),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_598),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_378),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_495),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_206),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_128),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_294),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_506),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_284),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_6),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_15),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_565),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_491),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_220),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_331),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_45),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_214),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_128),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_247),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_42),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_295),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_597),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_518),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_185),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_227),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_217),
.Y(n_733)
);

XNOR2x1_ASAP7_75t_L g734 ( 
.A(n_407),
.B(n_462),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_133),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_107),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_432),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_556),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_470),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_94),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_165),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_411),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_50),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_243),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_19),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_481),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_338),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_178),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_585),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_277),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_239),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_413),
.B(n_582),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_105),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_102),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_200),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_607),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_423),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_183),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_289),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_227),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_275),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_240),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_129),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_464),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_399),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_299),
.B(n_53),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_437),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_555),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_359),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_235),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_450),
.Y(n_771)
);

CKINVDCx16_ASAP7_75t_R g772 ( 
.A(n_542),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_249),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_467),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_63),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_132),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_334),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_191),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_201),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_564),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_12),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_60),
.Y(n_782)
);

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_16),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_362),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_253),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_238),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_150),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_357),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_513),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_290),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_202),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_266),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_335),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_96),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_2),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_23),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_267),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_533),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_381),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_264),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_490),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_167),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_577),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_539),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_469),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_119),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_85),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_87),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_178),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_563),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_47),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_486),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_328),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_43),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_468),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_367),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_127),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_46),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_203),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_522),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_318),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_474),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_27),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_343),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_260),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_57),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_422),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_66),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_56),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_56),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_596),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_471),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_252),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_226),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_296),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_244),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_587),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_458),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_599),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_344),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_223),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_121),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_268),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_211),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_365),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_108),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_209),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_234),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_400),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_216),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_1),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_482),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_229),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_70),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_434),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_428),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_500),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_285),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_371),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_258),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_608),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_189),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_149),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_324),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_212),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_169),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_454),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_236),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_574),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_278),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_117),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_552),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_219),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_20),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_354),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_356),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_99),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_12),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_104),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_444),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_327),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_132),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_211),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_37),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_8),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_499),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_166),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_457),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_119),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_390),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_418),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_213),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_287),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_173),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_228),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_187),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_180),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_498),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_504),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_203),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_193),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_384),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_125),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_224),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_103),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_438),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_363),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_416),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_157),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_257),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_10),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_68),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_136),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_84),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_459),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_237),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_32),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_405),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_270),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_261),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_265),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_206),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_568),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_16),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_576),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_69),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_410),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_39),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_207),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_105),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_435),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_497),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_219),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_430),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_10),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_553),
.Y(n_936)
);

CKINVDCx16_ASAP7_75t_R g937 ( 
.A(n_104),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_91),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_62),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_208),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_509),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_517),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_280),
.Y(n_943)
);

XNOR2xp5_ASAP7_75t_L g944 ( 
.A(n_174),
.B(n_447),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_535),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_425),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_92),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_409),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_605),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_393),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_17),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_87),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_580),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_210),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_238),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_97),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_165),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_251),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_588),
.Y(n_959)
);

INVxp67_ASAP7_75t_SL g960 ( 
.A(n_33),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_567),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_240),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_302),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_115),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_100),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_245),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_230),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_197),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_401),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_0),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_61),
.Y(n_971)
);

INVxp33_ASAP7_75t_L g972 ( 
.A(n_63),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_571),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_95),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_307),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_103),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_271),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_112),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_85),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_149),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_215),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_215),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_45),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_551),
.Y(n_984)
);

BUFx5_ASAP7_75t_L g985 ( 
.A(n_157),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_32),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_214),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_204),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_125),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_279),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_442),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_452),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_113),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_42),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_398),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_234),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_584),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_193),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_170),
.Y(n_999)
);

CKINVDCx16_ASAP7_75t_R g1000 ( 
.A(n_414),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_453),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_188),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_27),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_248),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_185),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_96),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_322),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_120),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_231),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_225),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_389),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_310),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_375),
.Y(n_1013)
);

INVxp33_ASAP7_75t_SL g1014 ( 
.A(n_557),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_333),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_250),
.Y(n_1016)
);

BUFx2_ASAP7_75t_SL g1017 ( 
.A(n_44),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_233),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_197),
.Y(n_1019)
);

BUFx10_ASAP7_75t_L g1020 ( 
.A(n_532),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_242),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_408),
.Y(n_1022)
);

BUFx5_ASAP7_75t_L g1023 ( 
.A(n_426),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_228),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_548),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_40),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_420),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_139),
.Y(n_1028)
);

CKINVDCx16_ASAP7_75t_R g1029 ( 
.A(n_232),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_195),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_319),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_31),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_341),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_223),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_58),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_476),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_427),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_403),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_241),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_5),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_443),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_36),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_46),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_572),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_116),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_138),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_744),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_R g1048 ( 
.A1(n_611),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_652),
.B(n_3),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_635),
.B(n_4),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_744),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_707),
.B(n_4),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_706),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_693),
.B(n_5),
.Y(n_1054)
);

OA21x2_ASAP7_75t_L g1055 ( 
.A1(n_695),
.A2(n_7),
.B(n_9),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_635),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_744),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_620),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_665),
.Y(n_1059)
);

INVx6_ASAP7_75t_L g1060 ( 
.A(n_665),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_618),
.A2(n_255),
.B(n_254),
.Y(n_1061)
);

OA21x2_ASAP7_75t_L g1062 ( 
.A1(n_695),
.A2(n_7),
.B(n_11),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_828),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_730),
.B(n_13),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_730),
.B(n_13),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_783),
.B(n_14),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_705),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_744),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_985),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_749),
.B(n_14),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_749),
.B(n_17),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_707),
.B(n_18),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_612),
.B(n_18),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_620),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_855),
.B(n_19),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_985),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_854),
.B(n_21),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_790),
.A2(n_21),
.B(n_22),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_985),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_985),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_652),
.B(n_22),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_972),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_985),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_706),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_754),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_754),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_654),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_738),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_797),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_754),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_754),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_770),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_770),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_654),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_686),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_770),
.Y(n_1096)
);

AOI22x1_ASAP7_75t_SL g1097 ( 
.A1(n_626),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_770),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_SL g1099 ( 
.A(n_640),
.B(n_26),
.Y(n_1099)
);

CKINVDCx11_ASAP7_75t_R g1100 ( 
.A(n_718),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_686),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_790),
.A2(n_28),
.B(n_29),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_763),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_741),
.B(n_28),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_621),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_797),
.Y(n_1106)
);

AND2x2_ASAP7_75t_SL g1107 ( 
.A(n_645),
.B(n_30),
.Y(n_1107)
);

BUFx8_ASAP7_75t_SL g1108 ( 
.A(n_723),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_1020),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_854),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_964),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_900),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_937),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_900),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_703),
.B(n_34),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_855),
.B(n_34),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_900),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_900),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_763),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_830),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_830),
.Y(n_1121)
);

BUFx8_ASAP7_75t_SL g1122 ( 
.A(n_823),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_873),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_655),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_964),
.B(n_35),
.Y(n_1125)
);

AND2x6_ASAP7_75t_L g1126 ( 
.A(n_636),
.B(n_259),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_902),
.B(n_37),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_873),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1016),
.B(n_38),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_879),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_965),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1131)
);

OA21x2_ASAP7_75t_L g1132 ( 
.A1(n_800),
.A2(n_44),
.B(n_47),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_655),
.Y(n_1133)
);

AOI22x1_ASAP7_75t_SL g1134 ( 
.A1(n_829),
.A2(n_52),
.B1(n_49),
.B2(n_51),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_879),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1020),
.Y(n_1136)
);

CKINVDCx11_ASAP7_75t_R g1137 ( 
.A(n_848),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_871),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_708),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1016),
.B(n_49),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_889),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1021),
.B(n_51),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1029),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_636),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_902),
.B(n_54),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_889),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_636),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_897),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_622),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_897),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_649),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_917),
.Y(n_1152)
);

CKINVDCx8_ASAP7_75t_R g1153 ( 
.A(n_1017),
.Y(n_1153)
);

CKINVDCx16_ASAP7_75t_R g1154 ( 
.A(n_651),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1021),
.B(n_55),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_972),
.A2(n_58),
.B1(n_55),
.B2(n_57),
.Y(n_1156)
);

INVx5_ASAP7_75t_L g1157 ( 
.A(n_649),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_960),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_662),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_809),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_649),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_614),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_702),
.A2(n_64),
.B1(n_59),
.B2(n_62),
.Y(n_1163)
);

BUFx8_ASAP7_75t_L g1164 ( 
.A(n_716),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_910),
.B(n_64),
.Y(n_1165)
);

AND2x2_ASAP7_75t_SL g1166 ( 
.A(n_772),
.B(n_65),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1000),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_628),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_771),
.B(n_67),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_792),
.B(n_70),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_888),
.B(n_71),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_703),
.B(n_71),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_677),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_613),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_927),
.B(n_72),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_SL g1176 ( 
.A1(n_909),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1036),
.B(n_74),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_809),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_619),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_677),
.Y(n_1180)
);

OAI22x1_ASAP7_75t_SL g1181 ( 
.A1(n_912),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1181)
);

OA22x2_ASAP7_75t_SL g1182 ( 
.A1(n_960),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_615),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_677),
.Y(n_1184)
);

AND2x6_ASAP7_75t_L g1185 ( 
.A(n_784),
.B(n_263),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_644),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_784),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_910),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_610),
.B(n_82),
.Y(n_1189)
);

CKINVDCx6p67_ASAP7_75t_R g1190 ( 
.A(n_1100),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1154),
.B(n_1014),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1090),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1047),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1060),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1099),
.B(n_766),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1091),
.Y(n_1196)
);

AND2x6_ASAP7_75t_L g1197 ( 
.A(n_1052),
.B(n_784),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1092),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1119),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1117),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1105),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1137),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1067),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1051),
.B(n_1057),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1064),
.B(n_860),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1113),
.A2(n_755),
.B1(n_986),
.B2(n_926),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1068),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1072),
.B(n_650),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1059),
.B(n_761),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1149),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1068),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1085),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1085),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1093),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1131),
.A2(n_755),
.B1(n_1024),
.B2(n_1019),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1093),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1096),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1108),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1098),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1112),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1183),
.B(n_780),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1114),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1071),
.A2(n_752),
.B(n_860),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1109),
.B(n_969),
.Y(n_1225)
);

AND3x2_ASAP7_75t_L g1226 ( 
.A(n_1169),
.B(n_1171),
.C(n_1170),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1118),
.B(n_991),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1075),
.B(n_991),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1143),
.A2(n_701),
.B1(n_743),
.B2(n_623),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1168),
.B(n_780),
.Y(n_1230)
);

BUFx10_ASAP7_75t_L g1231 ( 
.A(n_1060),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1086),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1151),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1136),
.B(n_1166),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1119),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1151),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1153),
.B(n_992),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1120),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1120),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1163),
.A2(n_806),
.B1(n_819),
.B2(n_802),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1125),
.A2(n_904),
.B1(n_956),
.B2(n_1040),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1126),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1152),
.B(n_631),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1121),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1173),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1116),
.B(n_800),
.Y(n_1246)
);

NOR2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1088),
.B(n_869),
.Y(n_1247)
);

INVxp33_ASAP7_75t_SL g1248 ( 
.A(n_1053),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1058),
.B(n_869),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1089),
.B(n_931),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1180),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1121),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1180),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1126),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1128),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1127),
.B(n_810),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1128),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1148),
.Y(n_1258)
);

INVx8_ASAP7_75t_L g1259 ( 
.A(n_1162),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1150),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1074),
.B(n_931),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1150),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1145),
.B(n_810),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1106),
.B(n_936),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1079),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1135),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1080),
.B(n_639),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1069),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1175),
.B(n_936),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1174),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1179),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1061),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1144),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_L g1274 ( 
.A(n_1177),
.B(n_1035),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1076),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1083),
.B(n_1049),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1122),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1087),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1165),
.B(n_812),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1094),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1056),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1110),
.B(n_812),
.Y(n_1282)
);

INVxp67_ASAP7_75t_R g1283 ( 
.A(n_1048),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1184),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1095),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1049),
.B(n_663),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1081),
.B(n_616),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1187),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_1084),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1101),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1139),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1124),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1103),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1123),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1081),
.B(n_617),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1130),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1141),
.B(n_1158),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1133),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1158),
.B(n_668),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1146),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1115),
.B(n_638),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1115),
.B(n_1172),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1172),
.B(n_890),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1160),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1189),
.B(n_648),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1178),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_L g1307 ( 
.A(n_1073),
.B(n_1045),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1063),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1063),
.B(n_678),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1138),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1104),
.B(n_656),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_SL g1312 ( 
.A(n_1129),
.B(n_1140),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1147),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1188),
.A2(n_878),
.B1(n_924),
.B2(n_847),
.Y(n_1314)
);

BUFx4f_ASAP7_75t_L g1315 ( 
.A(n_1126),
.Y(n_1315)
);

NOR2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1050),
.B(n_773),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1142),
.B(n_661),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1111),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1157),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1157),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1157),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1161),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1161),
.B(n_680),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1111),
.B(n_681),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1161),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1055),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1155),
.B(n_1039),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1062),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1062),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1078),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1102),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1054),
.B(n_890),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1102),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1132),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1082),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_L g1336 ( 
.A(n_1156),
.B(n_980),
.C(n_957),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1182),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1139),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1066),
.B(n_734),
.C(n_667),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1186),
.A2(n_630),
.B(n_629),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1185),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1185),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1159),
.A2(n_633),
.B(n_632),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1167),
.B(n_684),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1077),
.B(n_671),
.C(n_666),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1077),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1164),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1164),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1176),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1181),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1097),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1134),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1134),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1058),
.B(n_672),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1090),
.B(n_689),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1090),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1090),
.B(n_690),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1154),
.B(n_682),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1105),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1090),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1064),
.B(n_634),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1090),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1090),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1064),
.B(n_641),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1067),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1105),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1090),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1047),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1090),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1047),
.Y(n_1370)
);

AND2x2_ASAP7_75t_SL g1371 ( 
.A(n_1107),
.B(n_625),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1090),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1060),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1047),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1183),
.B(n_709),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1090),
.B(n_711),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1090),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1090),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1047),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1154),
.B(n_683),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1090),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1090),
.B(n_714),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1119),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1047),
.Y(n_1384)
);

NAND3xp33_ASAP7_75t_L g1385 ( 
.A(n_1099),
.B(n_688),
.C(n_685),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1060),
.Y(n_1386)
);

INVxp33_ASAP7_75t_L g1387 ( 
.A(n_1183),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1090),
.B(n_720),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1119),
.Y(n_1389)
);

NAND2xp33_ASAP7_75t_L g1390 ( 
.A(n_1052),
.B(n_1032),
.Y(n_1390)
);

INVxp33_ASAP7_75t_L g1391 ( 
.A(n_1183),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1154),
.B(n_694),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1047),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1047),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1052),
.B(n_699),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1090),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1119),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1090),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1183),
.B(n_729),
.Y(n_1399)
);

CKINVDCx14_ASAP7_75t_R g1400 ( 
.A(n_1053),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1047),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1154),
.B(n_713),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1047),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1090),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1108),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1047),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1090),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1064),
.B(n_642),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1183),
.B(n_742),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1105),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_L g1411 ( 
.A(n_1052),
.B(n_717),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1090),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1090),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1047),
.Y(n_1414)
);

NOR2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1067),
.B(n_624),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1060),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1060),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1154),
.B(n_721),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1064),
.B(n_647),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1047),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1099),
.B(n_725),
.C(n_724),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1047),
.Y(n_1422)
);

XOR2xp5_ASAP7_75t_L g1423 ( 
.A(n_1154),
.B(n_646),
.Y(n_1423)
);

INVxp33_ASAP7_75t_L g1424 ( 
.A(n_1183),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1154),
.B(n_733),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1064),
.B(n_657),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1125),
.A2(n_1042),
.B1(n_1043),
.B2(n_1030),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1125),
.A2(n_1046),
.B1(n_637),
.B2(n_643),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1090),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1154),
.B(n_735),
.Y(n_1430)
);

INVxp33_ASAP7_75t_L g1431 ( 
.A(n_1183),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1047),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1047),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1154),
.B(n_736),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1047),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_L g1436 ( 
.A(n_1052),
.B(n_748),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1067),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1154),
.B(n_753),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1090),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1047),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1090),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1099),
.A2(n_664),
.B1(n_676),
.B2(n_659),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1047),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1090),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1278),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1212),
.B(n_746),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1280),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1297),
.B(n_758),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1212),
.B(n_747),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1266),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1205),
.B(n_760),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1373),
.B(n_691),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1285),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1290),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1205),
.B(n_778),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1228),
.B(n_757),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1233),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1228),
.B(n_779),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1195),
.B(n_782),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1373),
.B(n_1417),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1302),
.B(n_764),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1417),
.B(n_722),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1361),
.B(n_786),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1361),
.B(n_787),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1385),
.B(n_728),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1339),
.A2(n_774),
.B1(n_820),
.B2(n_768),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1339),
.A2(n_796),
.B1(n_811),
.B2(n_791),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1236),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1302),
.B(n_769),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1385),
.B(n_867),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1371),
.A2(n_997),
.B1(n_1013),
.B2(n_946),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1308),
.B(n_814),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1276),
.A2(n_660),
.B(n_658),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1332),
.B(n_785),
.Y(n_1474)
);

NOR2xp67_ASAP7_75t_L g1475 ( 
.A(n_1242),
.B(n_793),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_L g1476 ( 
.A(n_1197),
.B(n_1025),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1421),
.B(n_1332),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1246),
.B(n_801),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1293),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1294),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1296),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1266),
.B(n_1299),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1256),
.B(n_803),
.Y(n_1483)
);

NAND2xp33_ASAP7_75t_L g1484 ( 
.A(n_1197),
.B(n_784),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1256),
.B(n_805),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1263),
.A2(n_726),
.B1(n_727),
.B2(n_627),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1263),
.A2(n_696),
.B(n_715),
.C(n_687),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1279),
.B(n_816),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1201),
.B(n_858),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1364),
.B(n_818),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1347),
.B(n_1027),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1364),
.B(n_836),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1359),
.B(n_821),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1300),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1270),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1387),
.B(n_944),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1366),
.B(n_1309),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1249),
.B(n_653),
.Y(n_1498)
);

AO22x2_ASAP7_75t_L g1499 ( 
.A1(n_1337),
.A2(n_675),
.B1(n_697),
.B2(n_670),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1326),
.A2(n_817),
.B(n_877),
.C(n_745),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1251),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_SL g1502 ( 
.A(n_1347),
.B(n_1210),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1271),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1408),
.B(n_841),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1324),
.B(n_832),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1273),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1261),
.B(n_698),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1442),
.B(n_864),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1253),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1408),
.A2(n_1034),
.B1(n_884),
.B2(n_712),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1303),
.B(n_824),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1442),
.B(n_845),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1265),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1419),
.B(n_1426),
.C(n_1427),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1391),
.B(n_1424),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1419),
.B(n_842),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1204),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1277),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1303),
.B(n_825),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_SL g1520 ( 
.A(n_1338),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1267),
.B(n_833),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1267),
.B(n_835),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1431),
.B(n_840),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1199),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1426),
.B(n_1286),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1312),
.A2(n_731),
.B1(n_732),
.B2(n_700),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1210),
.B(n_849),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1268),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1273),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1275),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1292),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1298),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1230),
.B(n_846),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1355),
.B(n_852),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1316),
.B(n_1247),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1192),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1357),
.B(n_876),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1335),
.A2(n_853),
.B1(n_862),
.B2(n_850),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1357),
.B(n_880),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1376),
.B(n_886),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1376),
.B(n_898),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1382),
.B(n_899),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1383),
.B(n_1389),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1382),
.B(n_908),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1344),
.A2(n_892),
.B1(n_894),
.B2(n_885),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1354),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1388),
.B(n_915),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1410),
.B(n_1305),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1388),
.B(n_921),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1427),
.B(n_923),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1208),
.B(n_895),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1196),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1198),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1397),
.Y(n_1554)
);

AND2x4_ASAP7_75t_SL g1555 ( 
.A(n_1231),
.B(n_788),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1428),
.B(n_963),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1200),
.Y(n_1557)
);

BUFx5_ASAP7_75t_L g1558 ( 
.A(n_1328),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1233),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1222),
.B(n_896),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1203),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1284),
.Y(n_1562)
);

AND2x4_ASAP7_75t_SL g1563 ( 
.A(n_1231),
.B(n_788),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1356),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1360),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1234),
.A2(n_990),
.B1(n_1001),
.B2(n_977),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1362),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1375),
.B(n_1044),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1323),
.B(n_1007),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1241),
.B(n_1028),
.C(n_911),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1224),
.B(n_1015),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1363),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1399),
.B(n_1041),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1409),
.B(n_1237),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1367),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1344),
.A2(n_913),
.B1(n_916),
.B2(n_901),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1206),
.A2(n_938),
.B1(n_967),
.B2(n_928),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1369),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1372),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1365),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1377),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1358),
.B(n_929),
.Y(n_1582)
);

INVxp33_ASAP7_75t_L g1583 ( 
.A(n_1282),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1259),
.B(n_1291),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1321),
.B(n_669),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1322),
.B(n_673),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1329),
.A2(n_740),
.B1(n_762),
.B2(n_751),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1245),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1325),
.B(n_674),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1241),
.B(n_930),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1219),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1380),
.B(n_933),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1209),
.B(n_935),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1378),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1288),
.B(n_679),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1245),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1392),
.B(n_951),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1313),
.B(n_692),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1207),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1381),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1396),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1398),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1211),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1336),
.A2(n_776),
.B1(n_781),
.B2(n_775),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1395),
.A2(n_966),
.B1(n_968),
.B2(n_962),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1225),
.B(n_970),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1319),
.B(n_704),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1437),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1315),
.B(n_971),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1390),
.A2(n_982),
.B1(n_983),
.B2(n_974),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1320),
.B(n_710),
.Y(n_1611)
);

OAI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1282),
.A2(n_1336),
.B1(n_1411),
.B2(n_1436),
.C(n_1327),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1255),
.Y(n_1613)
);

BUFx4f_ASAP7_75t_L g1614 ( 
.A(n_1259),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1243),
.B(n_719),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1240),
.B(n_989),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1206),
.A2(n_999),
.B1(n_1003),
.B2(n_994),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1217),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1318),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1240),
.B(n_1004),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1404),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1407),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1412),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1402),
.B(n_1005),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1218),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_SL g1626 ( 
.A(n_1289),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1243),
.B(n_737),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1221),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1418),
.B(n_1009),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1216),
.A2(n_1018),
.B1(n_1026),
.B2(n_1010),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1281),
.B(n_794),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1413),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1223),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1345),
.A2(n_807),
.B1(n_808),
.B2(n_795),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1194),
.B(n_826),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1386),
.B(n_834),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1314),
.B(n_788),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1216),
.A2(n_851),
.B1(n_863),
.B2(n_844),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1429),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1226),
.B(n_1235),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1330),
.A2(n_1331),
.B1(n_1334),
.B2(n_1333),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1314),
.B(n_815),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1229),
.B(n_815),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1423),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1214),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1226),
.B(n_865),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1229),
.B(n_815),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1343),
.A2(n_868),
.B1(n_874),
.B2(n_866),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1214),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1439),
.B(n_750),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1405),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_L g1652 ( 
.A(n_1341),
.B(n_1025),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1416),
.B(n_1025),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1255),
.Y(n_1654)
);

BUFx8_ASAP7_75t_L g1655 ( 
.A(n_1351),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1220),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1220),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1370),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1370),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1441),
.B(n_756),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1444),
.B(n_759),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1345),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1233),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1232),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1317),
.B(n_882),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1269),
.A2(n_767),
.B(n_765),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_L g1667 ( 
.A(n_1342),
.B(n_1025),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1250),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1248),
.B(n_739),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1191),
.B(n_1038),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1425),
.B(n_777),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1430),
.B(n_1037),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1264),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1414),
.Y(n_1674)
);

INVx8_ASAP7_75t_L g1675 ( 
.A(n_1259),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1420),
.B(n_883),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1434),
.B(n_789),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1415),
.Y(n_1678)
);

INVxp33_ASAP7_75t_L g1679 ( 
.A(n_1346),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1438),
.B(n_798),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1443),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1238),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1254),
.B(n_799),
.Y(n_1683)
);

INVx4_ASAP7_75t_L g1684 ( 
.A(n_1254),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1287),
.B(n_804),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1311),
.A2(n_1295),
.B1(n_1301),
.B2(n_1340),
.Y(n_1686)
);

INVxp33_ASAP7_75t_L g1687 ( 
.A(n_1227),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1641),
.A2(n_1274),
.B(n_1307),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1525),
.B(n_1272),
.Y(n_1689)
);

BUFx12f_ASAP7_75t_L g1690 ( 
.A(n_1584),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1687),
.B(n_1400),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1495),
.Y(n_1692)
);

AO32x2_ASAP7_75t_L g1693 ( 
.A1(n_1686),
.A2(n_1545),
.A3(n_1471),
.B1(n_1538),
.B2(n_1684),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1503),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1457),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1583),
.B(n_1343),
.Y(n_1696)
);

AO21x1_ASAP7_75t_L g1697 ( 
.A1(n_1477),
.A2(n_822),
.B(n_813),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1446),
.B(n_827),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1683),
.A2(n_1306),
.B(n_1304),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1548),
.B(n_1239),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1521),
.A2(n_1522),
.B(n_1534),
.Y(n_1702)
);

A2O1A1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1514),
.A2(n_837),
.B(n_838),
.C(n_831),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1543),
.B(n_1244),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1490),
.A2(n_839),
.B(n_856),
.C(n_843),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1445),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1662),
.A2(n_859),
.B1(n_861),
.B2(n_857),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1449),
.B(n_870),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1451),
.B(n_1289),
.Y(n_1709)
);

AOI21xp33_ASAP7_75t_L g1710 ( 
.A1(n_1492),
.A2(n_1349),
.B(n_875),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1537),
.A2(n_881),
.B(n_872),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1460),
.B(n_1252),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1539),
.A2(n_893),
.B(n_891),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1482),
.B(n_1257),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1543),
.B(n_1258),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1447),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1612),
.A2(n_1458),
.B1(n_1455),
.B2(n_1504),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1453),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1554),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1516),
.B(n_1348),
.Y(n_1720)
);

AND2x2_ASAP7_75t_SL g1721 ( 
.A(n_1466),
.B(n_1352),
.Y(n_1721)
);

OAI321xp33_ASAP7_75t_L g1722 ( 
.A1(n_1643),
.A2(n_914),
.A3(n_903),
.B1(n_922),
.B2(n_905),
.C(n_887),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1454),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1546),
.B(n_1310),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1619),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1479),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1540),
.A2(n_907),
.B(n_906),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1558),
.B(n_918),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1456),
.A2(n_920),
.B1(n_925),
.B2(n_919),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1541),
.A2(n_934),
.B(n_932),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1542),
.A2(n_942),
.B(n_941),
.Y(n_1731)
);

AO21x1_ASAP7_75t_L g1732 ( 
.A1(n_1671),
.A2(n_945),
.B(n_943),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1448),
.B(n_1260),
.Y(n_1733)
);

AO32x2_ASAP7_75t_L g1734 ( 
.A1(n_1499),
.A2(n_1023),
.A3(n_947),
.B1(n_952),
.B2(n_940),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1536),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1647),
.A2(n_948),
.B1(n_950),
.B2(n_949),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1552),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1533),
.B(n_1450),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1544),
.A2(n_958),
.B(n_953),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1560),
.B(n_1262),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1457),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1558),
.B(n_959),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1608),
.Y(n_1743)
);

BUFx8_ASAP7_75t_L g1744 ( 
.A(n_1626),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1547),
.A2(n_973),
.B(n_961),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1631),
.B(n_1283),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1549),
.A2(n_984),
.B(n_975),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1480),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1461),
.A2(n_1011),
.B(n_995),
.Y(n_1749)
);

CKINVDCx10_ASAP7_75t_R g1750 ( 
.A(n_1626),
.Y(n_1750)
);

CKINVDCx10_ASAP7_75t_R g1751 ( 
.A(n_1520),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1469),
.A2(n_1022),
.B(n_1012),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1571),
.A2(n_1033),
.B(n_1031),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1481),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1553),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1557),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1515),
.B(n_1193),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1457),
.Y(n_1758)
);

INVxp67_ASAP7_75t_SL g1759 ( 
.A(n_1506),
.Y(n_1759)
);

NOR2xp67_ASAP7_75t_SL g1760 ( 
.A(n_1637),
.B(n_1642),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1459),
.A2(n_954),
.B1(n_955),
.B2(n_939),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1494),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1677),
.A2(n_1440),
.B1(n_1213),
.B2(n_1215),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_SL g1764 ( 
.A(n_1614),
.B(n_1190),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1613),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1564),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1565),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1567),
.Y(n_1768)
);

AO21x1_ASAP7_75t_L g1769 ( 
.A1(n_1685),
.A2(n_978),
.B(n_976),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1669),
.B(n_1368),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1582),
.B(n_1374),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1465),
.B(n_1379),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1569),
.A2(n_1519),
.B(n_1511),
.Y(n_1773)
);

OAI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1551),
.A2(n_981),
.B(n_979),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1478),
.B(n_1384),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1483),
.B(n_1393),
.Y(n_1776)
);

OAI321xp33_ASAP7_75t_L g1777 ( 
.A1(n_1634),
.A2(n_996),
.A3(n_988),
.B1(n_998),
.B2(n_993),
.C(n_987),
.Y(n_1777)
);

NAND2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1614),
.B(n_1529),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1485),
.B(n_1394),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1654),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1470),
.A2(n_1435),
.B1(n_1403),
.B2(n_1406),
.Y(n_1781)
);

CKINVDCx10_ASAP7_75t_R g1782 ( 
.A(n_1520),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1640),
.B(n_1401),
.Y(n_1783)
);

INVx5_ASAP7_75t_L g1784 ( 
.A(n_1675),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1488),
.B(n_1422),
.Y(n_1785)
);

A2O1A1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1500),
.A2(n_1006),
.B(n_1008),
.C(n_1002),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1474),
.A2(n_1433),
.B(n_1432),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1572),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1575),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1513),
.B(n_1615),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1627),
.A2(n_1475),
.B(n_1517),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1578),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1574),
.B(n_1202),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1472),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1508),
.B(n_1353),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1580),
.B(n_1353),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1646),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1592),
.B(n_1350),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1502),
.B(n_83),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1597),
.B(n_83),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1635),
.B(n_84),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1648),
.A2(n_89),
.B(n_86),
.C(n_88),
.Y(n_1802)
);

CKINVDCx10_ASAP7_75t_R g1803 ( 
.A(n_1584),
.Y(n_1803)
);

O2A1O1Ixp5_ASAP7_75t_L g1804 ( 
.A1(n_1473),
.A2(n_274),
.B(n_276),
.C(n_273),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1512),
.B(n_86),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1624),
.B(n_88),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1648),
.A2(n_282),
.B1(n_286),
.B2(n_281),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1579),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1595),
.A2(n_291),
.B(n_288),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1475),
.A2(n_293),
.B(n_292),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_SL g1811 ( 
.A(n_1675),
.B(n_89),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1581),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1629),
.B(n_90),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1587),
.A2(n_93),
.B1(n_90),
.B2(n_91),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1665),
.A2(n_298),
.B(n_297),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1487),
.A2(n_97),
.B(n_94),
.C(n_95),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1535),
.B(n_98),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1535),
.B(n_98),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1528),
.B(n_300),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1594),
.Y(n_1820)
);

OR2x6_ASAP7_75t_L g1821 ( 
.A(n_1675),
.B(n_99),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1530),
.B(n_301),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1636),
.B(n_101),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1590),
.A2(n_107),
.B(n_101),
.C(n_106),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1526),
.A2(n_304),
.B(n_303),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1531),
.B(n_305),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1532),
.B(n_308),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1600),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1559),
.Y(n_1829)
);

AOI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1598),
.A2(n_312),
.B(n_311),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1523),
.B(n_106),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1666),
.A2(n_315),
.B(n_314),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1561),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1601),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1568),
.A2(n_317),
.B(n_316),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1524),
.B(n_321),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1559),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1550),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_1838)
);

INVx5_ASAP7_75t_L g1839 ( 
.A(n_1559),
.Y(n_1839)
);

NOR2xp67_ASAP7_75t_L g1840 ( 
.A(n_1518),
.B(n_609),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1679),
.B(n_109),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1573),
.A2(n_1505),
.B(n_1609),
.Y(n_1842)
);

O2A1O1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1556),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1452),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1566),
.B(n_111),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1498),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1498),
.A2(n_325),
.B1(n_326),
.B2(n_323),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1674),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1576),
.A2(n_114),
.B(n_118),
.Y(n_1849)
);

BUFx12f_ASAP7_75t_L g1850 ( 
.A(n_1584),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1668),
.B(n_121),
.Y(n_1851)
);

AOI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1607),
.A2(n_330),
.B(n_329),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1602),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1621),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1489),
.B(n_122),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1622),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1562),
.B(n_336),
.Y(n_1857)
);

O2A1O1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1616),
.A2(n_1620),
.B(n_1680),
.C(n_1672),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1623),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1507),
.A2(n_1497),
.B1(n_1670),
.B2(n_1673),
.Y(n_1860)
);

NAND2x1p5_ASAP7_75t_L g1861 ( 
.A(n_1674),
.B(n_337),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1610),
.B(n_122),
.Y(n_1862)
);

NOR2xp67_ASAP7_75t_L g1863 ( 
.A(n_1644),
.B(n_339),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1476),
.A2(n_345),
.B(n_342),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1493),
.B(n_123),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1632),
.Y(n_1866)
);

O2A1O1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1467),
.A2(n_126),
.B(n_123),
.C(n_124),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1664),
.B(n_346),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_1527),
.B(n_347),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1639),
.B(n_348),
.Y(n_1870)
);

O2A1O1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1585),
.A2(n_131),
.B(n_127),
.C(n_129),
.Y(n_1871)
);

NAND3xp33_ASAP7_75t_L g1872 ( 
.A(n_1577),
.B(n_1630),
.C(n_1617),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1496),
.A2(n_350),
.B1(n_351),
.B2(n_349),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_1591),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1681),
.B(n_352),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1484),
.A2(n_355),
.B(n_353),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1468),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1611),
.B(n_358),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1577),
.A2(n_134),
.B1(n_131),
.B2(n_133),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1663),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1676),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1698),
.B(n_1499),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1692),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1874),
.Y(n_1884)
);

AOI221x1_ASAP7_75t_L g1885 ( 
.A1(n_1717),
.A2(n_1650),
.B1(n_1661),
.B2(n_1660),
.C(n_1589),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1738),
.B(n_1462),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_SL g1887 ( 
.A1(n_1825),
.A2(n_1586),
.B(n_1604),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1695),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1695),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1689),
.B(n_1605),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1743),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1694),
.Y(n_1892)
);

CKINVDCx11_ASAP7_75t_R g1893 ( 
.A(n_1690),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1702),
.A2(n_1667),
.B(n_1652),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1688),
.A2(n_1630),
.B1(n_1617),
.B2(n_1638),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1753),
.A2(n_1570),
.B(n_1593),
.Y(n_1896)
);

BUFx6f_ASAP7_75t_L g1897 ( 
.A(n_1741),
.Y(n_1897)
);

INVx4_ASAP7_75t_L g1898 ( 
.A(n_1784),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1790),
.B(n_1678),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1696),
.A2(n_1491),
.B1(n_1606),
.B2(n_1638),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1806),
.A2(n_1682),
.B1(n_1501),
.B2(n_1509),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1712),
.B(n_1555),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1735),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1699),
.B(n_1510),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1710),
.B(n_1674),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1706),
.Y(n_1906)
);

OAI21x1_ASAP7_75t_SL g1907 ( 
.A1(n_1815),
.A2(n_1486),
.B(n_1588),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1832),
.A2(n_1645),
.B(n_1596),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1719),
.B(n_1599),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_SL g1910 ( 
.A(n_1799),
.B(n_1651),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1708),
.B(n_1563),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1872),
.A2(n_1618),
.B(n_1603),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1813),
.A2(n_1656),
.B1(n_1657),
.B2(n_1649),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1773),
.A2(n_1628),
.B(n_1625),
.Y(n_1914)
);

AOI21xp33_ASAP7_75t_L g1915 ( 
.A1(n_1709),
.A2(n_1633),
.B(n_1658),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1741),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1794),
.B(n_1659),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1716),
.Y(n_1918)
);

INVx4_ASAP7_75t_L g1919 ( 
.A(n_1784),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1791),
.A2(n_1653),
.B(n_361),
.Y(n_1920)
);

AO31x2_ASAP7_75t_L g1921 ( 
.A1(n_1697),
.A2(n_1732),
.A3(n_1703),
.B(n_1728),
.Y(n_1921)
);

BUFx8_ASAP7_75t_L g1922 ( 
.A(n_1850),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1844),
.A2(n_368),
.B1(n_369),
.B2(n_366),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1718),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1775),
.A2(n_372),
.B(n_370),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1742),
.A2(n_374),
.B(n_373),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1723),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1737),
.Y(n_1928)
);

BUFx4f_ASAP7_75t_L g1929 ( 
.A(n_1778),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1760),
.B(n_134),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1858),
.A2(n_1805),
.B(n_1855),
.Y(n_1931)
);

AOI221x1_ASAP7_75t_L g1932 ( 
.A1(n_1810),
.A2(n_386),
.B1(n_606),
.B2(n_604),
.C(n_603),
.Y(n_1932)
);

AND3x4_ASAP7_75t_L g1933 ( 
.A(n_1783),
.B(n_1655),
.C(n_135),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1881),
.B(n_135),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1795),
.A2(n_1655),
.B1(n_379),
.B2(n_380),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_SL g1936 ( 
.A(n_1764),
.B(n_382),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1726),
.Y(n_1937)
);

OAI21x1_ASAP7_75t_L g1938 ( 
.A1(n_1700),
.A2(n_602),
.B(n_387),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1787),
.A2(n_601),
.B(n_388),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1776),
.B(n_136),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1748),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1779),
.B(n_137),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1785),
.B(n_138),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1865),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1860),
.B(n_394),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1842),
.A2(n_1804),
.B(n_1752),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1797),
.A2(n_396),
.B1(n_397),
.B2(n_395),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1754),
.Y(n_1948)
);

AO31x2_ASAP7_75t_L g1949 ( 
.A1(n_1769),
.A2(n_142),
.A3(n_140),
.B(n_141),
.Y(n_1949)
);

A2O1A1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1831),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_1744),
.Y(n_1951)
);

AO31x2_ASAP7_75t_L g1952 ( 
.A1(n_1705),
.A2(n_1729),
.A3(n_1807),
.B(n_1772),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1762),
.B(n_143),
.Y(n_1953)
);

AO31x2_ASAP7_75t_L g1954 ( 
.A1(n_1786),
.A2(n_146),
.A3(n_144),
.B(n_145),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1857),
.B(n_145),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1755),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1800),
.B(n_146),
.C(n_147),
.Y(n_1957)
);

OA21x2_ASAP7_75t_L g1958 ( 
.A1(n_1749),
.A2(n_406),
.B(n_404),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1857),
.B(n_412),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1714),
.B(n_1756),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_SL g1961 ( 
.A1(n_1835),
.A2(n_417),
.B(n_415),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1711),
.A2(n_421),
.B(n_419),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1870),
.A2(n_595),
.B(n_424),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1766),
.B(n_147),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1767),
.B(n_148),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1768),
.B(n_148),
.Y(n_1966)
);

A2O1A1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1849),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1833),
.B(n_151),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1788),
.B(n_152),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1746),
.B(n_1841),
.Y(n_1970)
);

A2O1A1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1774),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1868),
.A2(n_436),
.B(n_433),
.Y(n_1972)
);

OA21x2_ASAP7_75t_L g1973 ( 
.A1(n_1713),
.A2(n_445),
.B(n_441),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1765),
.B(n_448),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1814),
.A2(n_1736),
.B1(n_1862),
.B2(n_1845),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1771),
.A2(n_451),
.B(n_449),
.Y(n_1976)
);

AO21x1_ASAP7_75t_L g1977 ( 
.A1(n_1838),
.A2(n_153),
.B(n_154),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1840),
.B(n_456),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1808),
.Y(n_1979)
);

NAND3xp33_ASAP7_75t_L g1980 ( 
.A(n_1720),
.B(n_155),
.C(n_156),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1789),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1757),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1792),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1828),
.B(n_156),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1758),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1878),
.A2(n_463),
.B(n_461),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1796),
.B(n_158),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1727),
.A2(n_466),
.B(n_465),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1691),
.B(n_158),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1853),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1725),
.B(n_159),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1856),
.B(n_159),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1730),
.A2(n_1739),
.B(n_1731),
.Y(n_1993)
);

AOI21xp33_ASAP7_75t_L g1994 ( 
.A1(n_1721),
.A2(n_160),
.B(n_161),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1801),
.B(n_161),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1823),
.B(n_162),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1812),
.B(n_162),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1819),
.A2(n_477),
.B(n_472),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1780),
.B(n_478),
.Y(n_1999)
);

OAI21x1_ASAP7_75t_L g2000 ( 
.A1(n_1822),
.A2(n_480),
.B(n_479),
.Y(n_2000)
);

A2O1A1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1843),
.A2(n_163),
.B(n_164),
.C(n_166),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1745),
.A2(n_485),
.B(n_484),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1820),
.Y(n_2003)
);

INVx5_ASAP7_75t_L g2004 ( 
.A(n_1784),
.Y(n_2004)
);

INVx5_ASAP7_75t_L g2005 ( 
.A(n_1758),
.Y(n_2005)
);

INVx3_ASAP7_75t_L g2006 ( 
.A(n_1758),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1834),
.B(n_163),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1854),
.B(n_168),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1747),
.A2(n_489),
.B(n_488),
.Y(n_2009)
);

OAI21x1_ASAP7_75t_L g2010 ( 
.A1(n_1826),
.A2(n_593),
.B(n_494),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1733),
.A2(n_592),
.B1(n_589),
.B2(n_586),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1859),
.B(n_168),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1839),
.B(n_493),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1827),
.A2(n_578),
.B(n_570),
.Y(n_2014)
);

OAI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1931),
.A2(n_1886),
.B1(n_1890),
.B2(n_1895),
.Y(n_2015)
);

OAI21x1_ASAP7_75t_L g2016 ( 
.A1(n_1908),
.A2(n_1852),
.B(n_1830),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1970),
.B(n_1740),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1982),
.B(n_1798),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1883),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1891),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1903),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1902),
.B(n_1724),
.Y(n_2022)
);

AO31x2_ASAP7_75t_L g2023 ( 
.A1(n_1932),
.A2(n_1707),
.A3(n_1802),
.B(n_1761),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1946),
.A2(n_1839),
.B(n_1759),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1900),
.A2(n_1701),
.B1(n_1847),
.B2(n_1869),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1928),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1884),
.Y(n_2027)
);

BUFx12f_ASAP7_75t_L g2028 ( 
.A(n_1893),
.Y(n_2028)
);

INVx4_ASAP7_75t_L g2029 ( 
.A(n_2005),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1956),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1899),
.B(n_1836),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_R g2032 ( 
.A(n_2004),
.B(n_1817),
.Y(n_2032)
);

NAND3xp33_ASAP7_75t_L g2033 ( 
.A(n_1896),
.B(n_1818),
.C(n_1851),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1892),
.Y(n_2034)
);

NAND3x1_ASAP7_75t_L g2035 ( 
.A(n_1882),
.B(n_1793),
.C(n_1750),
.Y(n_2035)
);

OAI21x1_ASAP7_75t_L g2036 ( 
.A1(n_1914),
.A2(n_1809),
.B(n_1877),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1989),
.B(n_1704),
.Y(n_2037)
);

CKINVDCx6p67_ASAP7_75t_R g2038 ( 
.A(n_1951),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1960),
.B(n_1866),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1906),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1975),
.A2(n_1879),
.B1(n_1875),
.B2(n_1863),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1910),
.B(n_1911),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_SL g2043 ( 
.A(n_1945),
.B(n_1837),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1955),
.B(n_1770),
.Y(n_2044)
);

NOR2x1_ASAP7_75t_R g2045 ( 
.A(n_2004),
.B(n_1751),
.Y(n_2045)
);

AO21x2_ASAP7_75t_L g2046 ( 
.A1(n_1907),
.A2(n_1876),
.B(n_1864),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1904),
.A2(n_1824),
.B(n_1722),
.Y(n_2047)
);

AOI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_1994),
.A2(n_1777),
.B1(n_1867),
.B2(n_1846),
.C(n_1871),
.Y(n_2048)
);

AO22x2_ASAP7_75t_L g2049 ( 
.A1(n_1980),
.A2(n_1734),
.B1(n_1693),
.B2(n_1811),
.Y(n_2049)
);

OAI21x1_ASAP7_75t_L g2050 ( 
.A1(n_1894),
.A2(n_1829),
.B(n_1861),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1938),
.A2(n_1781),
.B(n_1816),
.Y(n_2051)
);

OAI21x1_ASAP7_75t_L g2052 ( 
.A1(n_1939),
.A2(n_1873),
.B(n_1763),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1963),
.A2(n_1693),
.B(n_1837),
.Y(n_2053)
);

AO21x2_ASAP7_75t_L g2054 ( 
.A1(n_1887),
.A2(n_1693),
.B(n_1734),
.Y(n_2054)
);

AO21x1_ASAP7_75t_L g2055 ( 
.A1(n_1920),
.A2(n_1930),
.B(n_1962),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_1922),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1918),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1917),
.B(n_1715),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1979),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1924),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1995),
.A2(n_1880),
.B1(n_1848),
.B2(n_1837),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1972),
.A2(n_1848),
.B(n_1839),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1909),
.Y(n_2063)
);

O2A1O1Ixp33_ASAP7_75t_SL g2064 ( 
.A1(n_2001),
.A2(n_1821),
.B(n_569),
.C(n_566),
.Y(n_2064)
);

AO31x2_ASAP7_75t_L g2065 ( 
.A1(n_1977),
.A2(n_169),
.A3(n_170),
.B(n_171),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_2000),
.A2(n_527),
.B(n_562),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_1968),
.Y(n_2067)
);

AOI21x1_ASAP7_75t_L g2068 ( 
.A1(n_1885),
.A2(n_1821),
.B(n_561),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1888),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1927),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_2010),
.A2(n_560),
.B(n_559),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1940),
.A2(n_550),
.B(n_547),
.Y(n_2072)
);

OA21x2_ASAP7_75t_L g2073 ( 
.A1(n_1912),
.A2(n_546),
.B(n_541),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_1888),
.Y(n_2074)
);

AOI22x1_ASAP7_75t_L g2075 ( 
.A1(n_1993),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_2075)
);

AO21x1_ASAP7_75t_L g2076 ( 
.A1(n_1988),
.A2(n_2009),
.B(n_2002),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1990),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1937),
.A2(n_1803),
.B1(n_1782),
.B2(n_538),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1889),
.Y(n_2079)
);

OAI21x1_ASAP7_75t_L g2080 ( 
.A1(n_1926),
.A2(n_537),
.B(n_536),
.Y(n_2080)
);

OR2x6_ASAP7_75t_L g2081 ( 
.A(n_1898),
.B(n_172),
.Y(n_2081)
);

AO21x2_ASAP7_75t_L g2082 ( 
.A1(n_1978),
.A2(n_531),
.B(n_528),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_SL g2083 ( 
.A1(n_1936),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_2083)
);

OAI21x1_ASAP7_75t_L g2084 ( 
.A1(n_1998),
.A2(n_525),
.B(n_524),
.Y(n_2084)
);

INVx8_ASAP7_75t_L g2085 ( 
.A(n_2005),
.Y(n_2085)
);

O2A1O1Ixp33_ASAP7_75t_SL g2086 ( 
.A1(n_1971),
.A2(n_523),
.B(n_521),
.C(n_520),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1941),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2003),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1948),
.Y(n_2089)
);

AOI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1942),
.A2(n_516),
.B(n_515),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1943),
.B(n_179),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1981),
.Y(n_2092)
);

BUFx4_ASAP7_75t_R g2093 ( 
.A(n_1929),
.Y(n_2093)
);

OAI21x1_ASAP7_75t_L g2094 ( 
.A1(n_2014),
.A2(n_514),
.B(n_512),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1983),
.Y(n_2095)
);

NAND2x1p5_ASAP7_75t_L g2096 ( 
.A(n_2005),
.B(n_501),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1974),
.B(n_1999),
.Y(n_2097)
);

AOI21x1_ASAP7_75t_L g2098 ( 
.A1(n_1913),
.A2(n_511),
.B(n_510),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1964),
.Y(n_2099)
);

NAND2x1p5_ASAP7_75t_L g2100 ( 
.A(n_2004),
.B(n_507),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1889),
.B(n_508),
.Y(n_2101)
);

OA21x2_ASAP7_75t_L g2102 ( 
.A1(n_1965),
.A2(n_1992),
.B(n_1984),
.Y(n_2102)
);

OA21x2_ASAP7_75t_L g2103 ( 
.A1(n_2053),
.A2(n_1969),
.B(n_1966),
.Y(n_2103)
);

INVx4_ASAP7_75t_L g2104 ( 
.A(n_2085),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_2027),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2040),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2040),
.Y(n_2107)
);

AOI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2015),
.A2(n_1967),
.B1(n_1950),
.B2(n_1944),
.C(n_1957),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2092),
.Y(n_2109)
);

NAND3xp33_ASAP7_75t_SL g2110 ( 
.A(n_2041),
.B(n_1935),
.C(n_1996),
.Y(n_2110)
);

CKINVDCx6p67_ASAP7_75t_R g2111 ( 
.A(n_2028),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2019),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2034),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2057),
.Y(n_2114)
);

OR2x6_ASAP7_75t_L g2115 ( 
.A(n_2085),
.B(n_1897),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_2018),
.B(n_1987),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2060),
.Y(n_2117)
);

OA21x2_ASAP7_75t_L g2118 ( 
.A1(n_2016),
.A2(n_2007),
.B(n_2012),
.Y(n_2118)
);

BUFx2_ASAP7_75t_L g2119 ( 
.A(n_2020),
.Y(n_2119)
);

OAI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_2047),
.A2(n_1961),
.B(n_1925),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2070),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2087),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2074),
.Y(n_2123)
);

OR2x2_ASAP7_75t_L g2124 ( 
.A(n_2017),
.B(n_1934),
.Y(n_2124)
);

AOI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_2076),
.A2(n_1905),
.B1(n_1953),
.B2(n_1959),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_2069),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2089),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2095),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_2063),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_2029),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2088),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2099),
.B(n_1952),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2021),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2067),
.B(n_1901),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2026),
.Y(n_2135)
);

INVx3_ASAP7_75t_L g2136 ( 
.A(n_2029),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_2079),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2031),
.B(n_1991),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_2042),
.A2(n_1933),
.B1(n_2008),
.B2(n_1997),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2058),
.B(n_1915),
.Y(n_2140)
);

BUFx2_ASAP7_75t_SL g2141 ( 
.A(n_2056),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2030),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_2059),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2077),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2039),
.B(n_1952),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_2038),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2022),
.B(n_1897),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2050),
.Y(n_2148)
);

AND2x6_ASAP7_75t_L g2149 ( 
.A(n_2101),
.B(n_2011),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2101),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2102),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2037),
.B(n_1916),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2091),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2033),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2032),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2065),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2065),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_2097),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2036),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2065),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2075),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_2097),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2044),
.B(n_2006),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2075),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2049),
.B(n_1985),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_2082),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2049),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2064),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2068),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2048),
.A2(n_1923),
.B1(n_1947),
.B2(n_1976),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2093),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2054),
.B(n_1916),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_2096),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2086),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_2100),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_2139),
.B(n_2025),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2124),
.B(n_2081),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2151),
.Y(n_2178)
);

INVx4_ASAP7_75t_L g2179 ( 
.A(n_2115),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_2130),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_2158),
.B(n_1919),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_2119),
.Y(n_2182)
);

HB1xp67_ASAP7_75t_L g2183 ( 
.A(n_2172),
.Y(n_2183)
);

BUFx2_ASAP7_75t_L g2184 ( 
.A(n_2126),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2134),
.B(n_2081),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2106),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2154),
.B(n_2043),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2107),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_2105),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2138),
.B(n_2083),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_2115),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2112),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2121),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2113),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2158),
.B(n_2061),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2153),
.B(n_2023),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2116),
.B(n_2078),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2116),
.B(n_1954),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2147),
.B(n_2023),
.Y(n_2199)
);

INVx4_ASAP7_75t_L g2200 ( 
.A(n_2115),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2114),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2140),
.B(n_2163),
.Y(n_2202)
);

AOI222xp33_ASAP7_75t_L g2203 ( 
.A1(n_2110),
.A2(n_2072),
.B1(n_2045),
.B2(n_2043),
.C1(n_2035),
.C2(n_2052),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2152),
.B(n_1954),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2145),
.B(n_2023),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2150),
.B(n_1949),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2109),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_2165),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2143),
.B(n_1921),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2143),
.B(n_1949),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2133),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2139),
.B(n_2013),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2117),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2122),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2171),
.B(n_1921),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2127),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2128),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2131),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2123),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2145),
.B(n_2024),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2162),
.B(n_2084),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2135),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_2162),
.B(n_2094),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2171),
.B(n_2090),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2132),
.B(n_2055),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2132),
.B(n_2073),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2144),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2142),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2165),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2108),
.B(n_2051),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2108),
.B(n_2046),
.Y(n_2231)
);

BUFx4f_ASAP7_75t_L g2232 ( 
.A(n_2111),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2167),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2123),
.B(n_2090),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2170),
.A2(n_2098),
.B1(n_1973),
.B2(n_1958),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2169),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_2156),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2157),
.Y(n_2238)
);

BUFx2_ASAP7_75t_L g2239 ( 
.A(n_2137),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2155),
.B(n_1958),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2160),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2155),
.B(n_1973),
.Y(n_2242)
);

BUFx2_ASAP7_75t_L g2243 ( 
.A(n_2129),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2146),
.B(n_2066),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2175),
.B(n_2071),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_2161),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2183),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2183),
.B(n_2199),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2202),
.B(n_2173),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_2176),
.B(n_2110),
.Y(n_2250)
);

INVx2_ASAP7_75t_SL g2251 ( 
.A(n_2182),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_2237),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2190),
.B(n_2173),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2215),
.B(n_2125),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2188),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2188),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_2191),
.B(n_2104),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2236),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2186),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2233),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2216),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2229),
.B(n_2125),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2204),
.B(n_2149),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2198),
.B(n_2149),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2212),
.B(n_2149),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2236),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2208),
.B(n_2164),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2191),
.B(n_2130),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2208),
.B(n_2149),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2177),
.B(n_2136),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2224),
.B(n_2136),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2197),
.B(n_2168),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2216),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2207),
.B(n_2141),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2196),
.B(n_2174),
.Y(n_2275)
);

INVx2_ASAP7_75t_SL g2276 ( 
.A(n_2182),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2217),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2192),
.B(n_2118),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2237),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2205),
.B(n_2118),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2192),
.B(n_2103),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2217),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2193),
.B(n_2103),
.Y(n_2283)
);

BUFx2_ASAP7_75t_L g2284 ( 
.A(n_2184),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_2219),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2238),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_2239),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2243),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2193),
.B(n_2120),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2241),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2246),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2185),
.B(n_2120),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2209),
.B(n_2159),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2246),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2194),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2205),
.B(n_2170),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2189),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2201),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2176),
.B(n_2148),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2213),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2214),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2187),
.B(n_2166),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2218),
.Y(n_2303)
);

OR2x2_ASAP7_75t_L g2304 ( 
.A(n_2248),
.B(n_2220),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_2268),
.B(n_2179),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2286),
.Y(n_2306)
);

INVx3_ASAP7_75t_L g2307 ( 
.A(n_2268),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2290),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2295),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2247),
.B(n_2271),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2250),
.B(n_2210),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2269),
.B(n_2220),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2260),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2250),
.B(n_2222),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2298),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_2269),
.B(n_2225),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_2285),
.B(n_2234),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2300),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2292),
.B(n_2227),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2267),
.B(n_2302),
.Y(n_2320)
);

AND2x2_ASAP7_75t_SL g2321 ( 
.A(n_2265),
.B(n_2232),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2285),
.B(n_2178),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2252),
.Y(n_2323)
);

OR2x2_ASAP7_75t_L g2324 ( 
.A(n_2267),
.B(n_2225),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2301),
.Y(n_2325)
);

INVxp67_ASAP7_75t_L g2326 ( 
.A(n_2287),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2257),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2264),
.B(n_2263),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2252),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_2284),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2270),
.B(n_2206),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2258),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2253),
.B(n_2240),
.Y(n_2333)
);

OR2x2_ASAP7_75t_L g2334 ( 
.A(n_2302),
.B(n_2226),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2289),
.B(n_2187),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2259),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2279),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2293),
.B(n_2226),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2266),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_2279),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2288),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2291),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2249),
.B(n_2242),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2266),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2274),
.B(n_2244),
.Y(n_2345)
);

OAI22xp33_ASAP7_75t_SL g2346 ( 
.A1(n_2314),
.A2(n_2262),
.B1(n_2231),
.B2(n_2230),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2310),
.B(n_2251),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2310),
.B(n_2345),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2309),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2306),
.Y(n_2350)
);

OR2x2_ASAP7_75t_L g2351 ( 
.A(n_2312),
.B(n_2320),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2306),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2308),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2315),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2308),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2318),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2317),
.B(n_2294),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2331),
.B(n_2276),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2334),
.B(n_2280),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_2317),
.B(n_2303),
.Y(n_2360)
);

HB1xp67_ASAP7_75t_L g2361 ( 
.A(n_2340),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2304),
.B(n_2316),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2343),
.B(n_2333),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_2341),
.B(n_2297),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2338),
.B(n_2280),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2313),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2323),
.B(n_2262),
.Y(n_2367)
);

INVxp67_ASAP7_75t_L g2368 ( 
.A(n_2325),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2336),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2311),
.B(n_2272),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_2329),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2361),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2362),
.B(n_2330),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2351),
.B(n_2335),
.Y(n_2374)
);

INVx3_ASAP7_75t_L g2375 ( 
.A(n_2360),
.Y(n_2375)
);

INVx1_ASAP7_75t_SL g2376 ( 
.A(n_2347),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2361),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2350),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2348),
.B(n_2326),
.Y(n_2379)
);

A2O1A1Ixp33_ASAP7_75t_L g2380 ( 
.A1(n_2370),
.A2(n_2321),
.B(n_2232),
.C(n_2254),
.Y(n_2380)
);

AOI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2370),
.A2(n_2203),
.B1(n_2195),
.B2(n_2319),
.Y(n_2381)
);

AOI322xp5_ASAP7_75t_L g2382 ( 
.A1(n_2363),
.A2(n_2328),
.A3(n_2296),
.B1(n_2342),
.B2(n_2337),
.C1(n_2231),
.C2(n_2322),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_2364),
.B(n_2327),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2352),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2373),
.B(n_2383),
.Y(n_2385)
);

AOI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_2381),
.A2(n_2360),
.B1(n_2346),
.B2(n_2357),
.Y(n_2386)
);

INVxp33_ASAP7_75t_L g2387 ( 
.A(n_2374),
.Y(n_2387)
);

OAI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2381),
.A2(n_2368),
.B(n_2346),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2378),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2382),
.B(n_2368),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2384),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2375),
.B(n_2358),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2372),
.B(n_2357),
.Y(n_2393)
);

OAI221xp5_ASAP7_75t_L g2394 ( 
.A1(n_2388),
.A2(n_2380),
.B1(n_2376),
.B2(n_2375),
.C(n_2377),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2390),
.A2(n_2367),
.B(n_2366),
.Y(n_2395)
);

OAI211xp5_ASAP7_75t_L g2396 ( 
.A1(n_2386),
.A2(n_2371),
.B(n_2369),
.C(n_2324),
.Y(n_2396)
);

NAND5xp2_ASAP7_75t_SL g2397 ( 
.A(n_2392),
.B(n_2379),
.C(n_2283),
.D(n_2281),
.E(n_2278),
.Y(n_2397)
);

O2A1O1Ixp5_ASAP7_75t_L g2398 ( 
.A1(n_2387),
.A2(n_2354),
.B(n_2349),
.C(n_2356),
.Y(n_2398)
);

AOI211xp5_ASAP7_75t_L g2399 ( 
.A1(n_2385),
.A2(n_2391),
.B(n_2389),
.C(n_2393),
.Y(n_2399)
);

AOI21xp5_ASAP7_75t_L g2400 ( 
.A1(n_2388),
.A2(n_2371),
.B(n_2359),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2388),
.A2(n_2355),
.B(n_2353),
.Y(n_2401)
);

NOR2x1_ASAP7_75t_L g2402 ( 
.A(n_2394),
.B(n_2257),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2395),
.B(n_2365),
.Y(n_2403)
);

NOR3x1_ASAP7_75t_L g2404 ( 
.A(n_2396),
.B(n_2296),
.C(n_2275),
.Y(n_2404)
);

AOI211xp5_ASAP7_75t_L g2405 ( 
.A1(n_2400),
.A2(n_1986),
.B(n_2322),
.C(n_2230),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2398),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2399),
.Y(n_2407)
);

NAND3xp33_ASAP7_75t_L g2408 ( 
.A(n_2401),
.B(n_2273),
.C(n_2261),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2407),
.B(n_2307),
.Y(n_2409)
);

OAI211xp5_ASAP7_75t_SL g2410 ( 
.A1(n_2405),
.A2(n_2397),
.B(n_2307),
.C(n_2327),
.Y(n_2410)
);

NOR2xp67_ASAP7_75t_L g2411 ( 
.A(n_2408),
.B(n_179),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2402),
.B(n_2305),
.Y(n_2412)
);

NOR3x1_ASAP7_75t_L g2413 ( 
.A(n_2409),
.B(n_2406),
.C(n_2403),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2411),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2412),
.B(n_2179),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2410),
.B(n_2404),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2414),
.Y(n_2417)
);

XNOR2xp5_ASAP7_75t_L g2418 ( 
.A(n_2416),
.B(n_181),
.Y(n_2418)
);

NOR2x1_ASAP7_75t_L g2419 ( 
.A(n_2415),
.B(n_2200),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2413),
.Y(n_2420)
);

INVxp67_ASAP7_75t_L g2421 ( 
.A(n_2414),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2414),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2417),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2420),
.A2(n_2200),
.B1(n_2282),
.B2(n_2277),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2422),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2418),
.B(n_181),
.Y(n_2426)
);

AOI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2421),
.A2(n_2344),
.B1(n_2339),
.B2(n_2332),
.Y(n_2427)
);

NOR4xp25_ASAP7_75t_L g2428 ( 
.A(n_2419),
.B(n_2228),
.C(n_183),
.D(n_184),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2428),
.B(n_182),
.Y(n_2429)
);

AOI22xp33_ASAP7_75t_L g2430 ( 
.A1(n_2423),
.A2(n_2255),
.B1(n_2256),
.B2(n_2223),
.Y(n_2430)
);

OAI22xp5_ASAP7_75t_SL g2431 ( 
.A1(n_2426),
.A2(n_2181),
.B1(n_2195),
.B2(n_186),
.Y(n_2431)
);

OAI21x1_ASAP7_75t_L g2432 ( 
.A1(n_2425),
.A2(n_2098),
.B(n_2180),
.Y(n_2432)
);

OA21x2_ASAP7_75t_L g2433 ( 
.A1(n_2424),
.A2(n_2080),
.B(n_2062),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_2429),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2433),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2431),
.A2(n_2430),
.B(n_2427),
.Y(n_2436)
);

OAI22x1_ASAP7_75t_L g2437 ( 
.A1(n_2432),
.A2(n_2181),
.B1(n_2211),
.B2(n_2180),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_SL g2438 ( 
.A1(n_2429),
.A2(n_182),
.B1(n_184),
.B2(n_187),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2429),
.B(n_188),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2438),
.B(n_2221),
.Y(n_2440)
);

OAI331xp33_ASAP7_75t_L g2441 ( 
.A1(n_2435),
.A2(n_189),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.B3(n_194),
.C1(n_195),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2439),
.Y(n_2442)
);

NAND2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2434),
.B(n_190),
.Y(n_2443)
);

AOI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2436),
.A2(n_2235),
.B(n_2245),
.Y(n_2444)
);

AO22x2_ASAP7_75t_L g2445 ( 
.A1(n_2442),
.A2(n_2440),
.B1(n_2441),
.B2(n_2444),
.Y(n_2445)
);

XOR2xp5_ASAP7_75t_L g2446 ( 
.A(n_2443),
.B(n_2437),
.Y(n_2446)
);

OAI21xp33_ASAP7_75t_L g2447 ( 
.A1(n_2442),
.A2(n_2299),
.B(n_2275),
.Y(n_2447)
);

OR5x1_ASAP7_75t_L g2448 ( 
.A(n_2441),
.B(n_192),
.C(n_194),
.D(n_196),
.E(n_200),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2446),
.B(n_2448),
.Y(n_2449)
);

XNOR2x1_ASAP7_75t_L g2450 ( 
.A(n_2449),
.B(n_2445),
.Y(n_2450)
);

AOI21xp33_ASAP7_75t_L g2451 ( 
.A1(n_2450),
.A2(n_2447),
.B(n_202),
.Y(n_2451)
);


endmodule