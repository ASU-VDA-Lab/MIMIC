module fake_aes_10577_n_657 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_657);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_657;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g91 ( .A(n_78), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_45), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_10), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_71), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_41), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_46), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
INVx2_ASAP7_75t_SL g101 ( .A(n_60), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_56), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_83), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_90), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_7), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_66), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_54), .B(n_86), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_88), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_80), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_48), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
INVxp33_ASAP7_75t_L g116 ( .A(n_59), .Y(n_116) );
BUFx10_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_26), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_10), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_24), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_23), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_69), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_13), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_50), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_34), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_28), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_4), .Y(n_129) );
INVxp33_ASAP7_75t_SL g130 ( .A(n_77), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_65), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_47), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_19), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_117), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_95), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_101), .B(n_0), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_101), .B(n_0), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_95), .B(n_106), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_126), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_106), .B(n_1), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
CKINVDCx6p67_ASAP7_75t_R g144 ( .A(n_91), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_116), .B(n_2), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_98), .B(n_2), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_117), .B(n_3), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_119), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_100), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_96), .B(n_3), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_120), .B(n_4), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_102), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_100), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
INVx1_ASAP7_75t_SL g162 ( .A(n_159), .Y(n_162) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
INVx8_ASAP7_75t_L g164 ( .A(n_154), .Y(n_164) );
INVx2_ASAP7_75t_SL g165 ( .A(n_144), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
INVxp67_ASAP7_75t_L g167 ( .A(n_159), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_135), .B(n_117), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_154), .B(n_120), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_154), .B(n_103), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_160), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_160), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_144), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
AND3x1_ASAP7_75t_L g180 ( .A(n_149), .B(n_133), .C(n_121), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_134), .B(n_108), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_135), .B(n_151), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_159), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_146), .B(n_96), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_146), .B(n_104), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_148), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
OAI22xp33_ASAP7_75t_SL g194 ( .A1(n_142), .A2(n_133), .B1(n_121), .B2(n_130), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_190), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_185), .B(n_145), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_185), .B(n_145), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_165), .B(n_145), .Y(n_199) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_163), .B(n_149), .Y(n_200) );
NOR2xp33_ASAP7_75t_SL g201 ( .A(n_165), .B(n_93), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_169), .B(n_151), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_172), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_169), .B(n_144), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_163), .A2(n_138), .B(n_136), .Y(n_206) );
BUFx12f_ASAP7_75t_L g207 ( .A(n_178), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_186), .Y(n_209) );
OR2x6_ASAP7_75t_L g210 ( .A(n_164), .B(n_149), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_164), .Y(n_212) );
OR2x6_ASAP7_75t_L g213 ( .A(n_164), .B(n_139), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_180), .B(n_157), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_167), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_175), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_186), .B(n_157), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_195), .B(n_141), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
INVxp67_ASAP7_75t_L g224 ( .A(n_188), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_163), .B(n_117), .Y(n_226) );
NOR2xp67_ASAP7_75t_L g227 ( .A(n_181), .B(n_141), .Y(n_227) );
INVx5_ASAP7_75t_L g228 ( .A(n_171), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_187), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_176), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_171), .B(n_150), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_177), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_180), .A2(n_137), .B1(n_150), .B2(n_152), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_163), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_170), .B(n_152), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_171), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_171), .Y(n_238) );
NAND2x1p5_ASAP7_75t_L g239 ( .A(n_181), .B(n_183), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_179), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_202), .B(n_171), .Y(n_242) );
OAI221xp5_ASAP7_75t_L g243 ( .A1(n_233), .A2(n_194), .B1(n_182), .B2(n_147), .C(n_158), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_196), .A2(n_183), .B(n_187), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_204), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_215), .A2(n_171), .B1(n_170), .B2(n_194), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_211), .B(n_178), .Y(n_248) );
INVx4_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_211), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_204), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_213), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_206), .A2(n_179), .B(n_171), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_196), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_197), .B(n_171), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_213), .A2(n_170), .B1(n_195), .B2(n_99), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g259 ( .A(n_233), .B(n_137), .C(n_138), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_225), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_213), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_220), .B(n_191), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_212), .B(n_170), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_225), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_228), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_205), .A2(n_187), .B(n_191), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_210), .B(n_189), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_212), .B(n_112), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_198), .B(n_189), .Y(n_270) );
HAxp5_ASAP7_75t_L g271 ( .A(n_220), .B(n_125), .CON(n_271), .SN(n_271) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_200), .B(n_104), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_208), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_213), .A2(n_161), .B1(n_142), .B2(n_158), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_213), .A2(n_161), .B1(n_139), .B2(n_147), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_224), .B(n_109), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_215), .A2(n_156), .B1(n_143), .B2(n_129), .Y(n_277) );
CKINVDCx6p67_ASAP7_75t_R g278 ( .A(n_210), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_236), .B(n_143), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_230), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_210), .B(n_107), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_210), .A2(n_143), .B1(n_156), .B2(n_110), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_236), .B(n_156), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_241), .Y(n_286) );
INVx6_ASAP7_75t_L g287 ( .A(n_249), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_249), .B(n_210), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_263), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_272), .B(n_200), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_263), .B(n_214), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_245), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_199), .B(n_240), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_272), .B(n_200), .Y(n_294) );
OAI222xp33_ASAP7_75t_L g295 ( .A1(n_258), .A2(n_203), .B1(n_209), .B2(n_215), .C1(n_226), .C2(n_221), .Y(n_295) );
BUFx4f_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_245), .Y(n_297) );
OAI22xp33_ASAP7_75t_L g298 ( .A1(n_247), .A2(n_201), .B1(n_217), .B2(n_215), .Y(n_298) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_274), .A2(n_226), .B1(n_236), .B2(n_201), .Y(n_299) );
BUFx12f_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_236), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_270), .B(n_222), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_256), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_278), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_272), .A2(n_239), .B1(n_222), .B2(n_227), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_276), .B(n_239), .Y(n_307) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_245), .Y(n_308) );
AOI32xp33_ASAP7_75t_L g309 ( .A1(n_243), .A2(n_124), .A3(n_105), .B1(n_132), .B2(n_115), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_268), .A2(n_239), .B1(n_227), .B2(n_237), .Y(n_310) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_275), .A2(n_235), .B(n_238), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_245), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_245), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_250), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g315 ( .A1(n_247), .A2(n_237), .B1(n_207), .B2(n_235), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_254), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_261), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_259), .A2(n_268), .B1(n_265), .B2(n_261), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_268), .A2(n_218), .B1(n_207), .B2(n_231), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_265), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_298), .A2(n_282), .B1(n_259), .B2(n_262), .Y(n_323) );
AO31x2_ASAP7_75t_L g324 ( .A1(n_306), .A2(n_280), .A3(n_253), .B(n_246), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g325 ( .A1(n_289), .A2(n_271), .B1(n_282), .B2(n_280), .C1(n_277), .C2(n_257), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_288), .B(n_254), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_288), .B(n_262), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_299), .A2(n_282), .B1(n_284), .B2(n_207), .Y(n_328) );
OAI21xp33_ASAP7_75t_SL g329 ( .A1(n_309), .A2(n_246), .B(n_273), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_291), .A2(n_271), .B1(n_242), .B2(n_250), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_286), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_302), .B(n_252), .Y(n_332) );
AOI31xp67_ASAP7_75t_L g333 ( .A1(n_286), .A2(n_140), .A3(n_155), .B(n_273), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_290), .B(n_271), .Y(n_334) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_290), .A2(n_253), .B1(n_252), .B2(n_285), .C(n_279), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_299), .A2(n_264), .B1(n_251), .B2(n_250), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_295), .A2(n_267), .B1(n_244), .B2(n_255), .C(n_240), .Y(n_337) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_318), .A2(n_155), .B(n_140), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_296), .B(n_228), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_299), .A2(n_251), .B1(n_269), .B2(n_218), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_293), .A2(n_248), .B(n_234), .Y(n_341) );
NAND2xp33_ASAP7_75t_SL g342 ( .A(n_294), .B(n_260), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
AOI21x1_ASAP7_75t_L g344 ( .A1(n_317), .A2(n_155), .B(n_140), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_294), .A2(n_251), .B1(n_218), .B2(n_234), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_320), .A2(n_230), .B1(n_208), .B2(n_216), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_315), .A2(n_216), .B1(n_219), .B2(n_232), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_216), .B1(n_219), .B2(n_232), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_303), .A2(n_140), .B(n_155), .Y(n_351) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_307), .A2(n_156), .B(n_94), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_321), .B(n_219), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_334), .B(n_332), .Y(n_355) );
NOR3xp33_ASAP7_75t_L g356 ( .A(n_330), .B(n_105), .C(n_131), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_329), .A2(n_296), .B1(n_288), .B2(n_316), .Y(n_358) );
OAI332xp33_ASAP7_75t_SL g359 ( .A1(n_327), .A2(n_343), .A3(n_348), .B1(n_334), .B2(n_310), .B3(n_325), .C1(n_11), .C2(n_12), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_352), .A2(n_123), .B(n_131), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_343), .B(n_292), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_325), .A2(n_300), .B1(n_296), .B2(n_316), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_329), .A2(n_337), .B(n_323), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_328), .A2(n_301), .B1(n_319), .B2(n_305), .C(n_311), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_348), .B(n_292), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_331), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_335), .A2(n_305), .B1(n_113), .B2(n_114), .C(n_128), .Y(n_367) );
OAI33xp33_ASAP7_75t_L g368 ( .A1(n_353), .A2(n_113), .A3(n_122), .B1(n_123), .B2(n_124), .B3(n_127), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_331), .B(n_313), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_347), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_335), .A2(n_287), .B1(n_314), .B2(n_132), .C(n_122), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_340), .A2(n_114), .B(n_127), .C(n_115), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_337), .A2(n_128), .B1(n_314), .B2(n_223), .C(n_232), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_324), .Y(n_374) );
AOI331xp33_ASAP7_75t_L g375 ( .A1(n_336), .A2(n_111), .A3(n_6), .B1(n_7), .B2(n_8), .B3(n_9), .C1(n_11), .Y(n_375) );
NOR3xp33_ASAP7_75t_L g376 ( .A(n_352), .B(n_312), .C(n_118), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_333), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_326), .A2(n_300), .B1(n_287), .B2(n_313), .Y(n_380) );
OAI31xp33_ASAP7_75t_L g381 ( .A1(n_342), .A2(n_312), .A3(n_308), .B(n_223), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_345), .B1(n_346), .B2(n_350), .C(n_353), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_357), .B(n_366), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_379), .Y(n_384) );
NOR3xp33_ASAP7_75t_L g385 ( .A(n_364), .B(n_339), .C(n_326), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_357), .B(n_324), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_324), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_366), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_366), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_377), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_362), .A2(n_126), .B(n_338), .C(n_351), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_377), .Y(n_392) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_367), .A2(n_341), .B(n_333), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
AOI33xp33_ASAP7_75t_L g395 ( .A1(n_358), .A2(n_326), .A3(n_6), .B1(n_8), .B2(n_9), .B3(n_13), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_327), .B1(n_326), .B2(n_287), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_379), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_374), .B(n_324), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_355), .B(n_324), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_369), .B(n_324), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_355), .B(n_338), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_369), .B(n_344), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_327), .B1(n_338), .B2(n_297), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_338), .Y(n_410) );
INVx4_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_361), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_363), .B(n_351), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_364), .B(n_344), .C(n_341), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_361), .B(n_327), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_365), .B(n_351), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_354), .B(n_327), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_367), .B(n_381), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_403), .B(n_381), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
NOR2x1_ASAP7_75t_SL g422 ( .A(n_396), .B(n_372), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_403), .B(n_380), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_400), .B(n_5), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_400), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_417), .B(n_5), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_412), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_405), .B(n_360), .Y(n_428) );
NAND4xp25_ASAP7_75t_L g429 ( .A(n_395), .B(n_356), .C(n_373), .D(n_372), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_391), .A2(n_360), .B(n_376), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_412), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g432 ( .A(n_395), .B(n_368), .C(n_373), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_418), .B(n_382), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_397), .Y(n_434) );
XNOR2x2_ASAP7_75t_L g435 ( .A(n_396), .B(n_375), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_418), .B(n_382), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_406), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_405), .B(n_360), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_417), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_385), .A2(n_359), .B(n_351), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_411), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_397), .B(n_14), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_388), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_416), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_405), .B(n_148), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_384), .Y(n_448) );
BUFx6f_ASAP7_75t_SL g449 ( .A(n_408), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_385), .B(n_359), .C(n_15), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_401), .B(n_153), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_404), .B(n_297), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_398), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_401), .B(n_153), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_388), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_401), .B(n_153), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_409), .A2(n_297), .B(n_228), .Y(n_457) );
OR2x6_ASAP7_75t_L g458 ( .A(n_404), .B(n_297), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_416), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_416), .B(n_14), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_410), .B(n_153), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_383), .B(n_16), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_418), .B(n_16), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_415), .B(n_17), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_406), .Y(n_466) );
NOR3xp33_ASAP7_75t_SL g467 ( .A(n_393), .B(n_399), .C(n_402), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_410), .B(n_153), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_443), .B(n_406), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_451), .B(n_404), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_421), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_433), .B(n_399), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_433), .A2(n_414), .B1(n_410), .B2(n_415), .C(n_413), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_437), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_446), .B(n_425), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_451), .B(n_404), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_420), .B(n_404), .Y(n_479) );
NOR2xp33_ASAP7_75t_SL g480 ( .A(n_465), .B(n_413), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_459), .B(n_389), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_436), .B(n_386), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_454), .B(n_456), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_454), .B(n_386), .Y(n_485) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_424), .B(n_411), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_434), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_456), .B(n_407), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_436), .B(n_386), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_428), .B(n_387), .Y(n_492) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_467), .A2(n_414), .B(n_409), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_428), .B(n_387), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_437), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_423), .B(n_390), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_439), .B(n_387), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_438), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_447), .B(n_390), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_445), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_455), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
AND4x1_ASAP7_75t_L g503 ( .A(n_465), .B(n_393), .C(n_18), .D(n_19), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_440), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_447), .B(n_461), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_466), .B(n_392), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_439), .B(n_383), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_462), .B(n_383), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_462), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_450), .B(n_415), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_458), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_468), .B(n_392), .Y(n_512) );
AO211x2_ASAP7_75t_L g513 ( .A1(n_419), .A2(n_429), .B(n_441), .C(n_435), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_464), .A2(n_411), .B1(n_415), .B2(n_407), .Y(n_514) );
NAND4xp25_ASAP7_75t_SL g515 ( .A(n_432), .B(n_394), .C(n_402), .D(n_398), .Y(n_515) );
XOR2xp5_ASAP7_75t_L g516 ( .A(n_422), .B(n_415), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_468), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_452), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_463), .B(n_394), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_426), .B(n_407), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_453), .Y(n_521) );
OAI322xp33_ASAP7_75t_L g522 ( .A1(n_435), .A2(n_411), .A3(n_153), .B1(n_398), .B2(n_407), .C1(n_22), .C2(n_23), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_444), .B(n_407), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_444), .B(n_408), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_448), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_448), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_442), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_492), .B(n_452), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_513), .A2(n_449), .B1(n_452), .B2(n_442), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_484), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_500), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_501), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_502), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_510), .A2(n_430), .B(n_457), .C(n_408), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_479), .B(n_411), .Y(n_536) );
XNOR2xp5_ASAP7_75t_L g537 ( .A(n_516), .B(n_458), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_513), .A2(n_510), .B(n_493), .Y(n_538) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_479), .B(n_17), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_476), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_489), .A2(n_449), .B1(n_408), .B2(n_153), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_472), .B(n_408), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_470), .B(n_18), .Y(n_543) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_487), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_472), .B(n_20), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_494), .B(n_153), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_482), .B(n_20), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_491), .B(n_21), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_497), .B(n_21), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_503), .B(n_22), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_483), .Y(n_552) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_489), .B(n_24), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_504), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_498), .B(n_25), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_497), .B(n_27), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_507), .B(n_29), .Y(n_557) );
XNOR2x1_ASAP7_75t_L g558 ( .A(n_469), .B(n_30), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_515), .A2(n_266), .B(n_260), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_480), .A2(n_281), .B(n_228), .C(n_260), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_473), .A2(n_166), .B1(n_173), .B2(n_174), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_481), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_506), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_507), .B(n_31), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_485), .B(n_33), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_485), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_508), .B(n_35), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_470), .B(n_478), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_508), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_38), .Y(n_570) );
XOR2xp5_ASAP7_75t_L g571 ( .A(n_505), .B(n_39), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_512), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_517), .Y(n_574) );
NAND3xp33_ASAP7_75t_SL g575 ( .A(n_469), .B(n_40), .C(n_42), .Y(n_575) );
AOI321xp33_ASAP7_75t_L g576 ( .A1(n_486), .A2(n_193), .A3(n_192), .B1(n_168), .B2(n_223), .C(n_53), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_489), .B(n_266), .Y(n_577) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_478), .B(n_43), .Y(n_578) );
OAI21xp33_ASAP7_75t_SL g579 ( .A1(n_498), .A2(n_49), .B(n_51), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_525), .B(n_52), .Y(n_580) );
NAND2xp33_ASAP7_75t_L g581 ( .A(n_511), .B(n_266), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_490), .Y(n_582) );
XOR2x2_ASAP7_75t_SL g583 ( .A(n_511), .B(n_55), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_521), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_518), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_522), .A2(n_266), .B(n_260), .C(n_166), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_526), .Y(n_587) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_519), .A2(n_281), .B(n_266), .C(n_260), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_527), .Y(n_589) );
AOI22xp5_ASAP7_75t_SL g590 ( .A1(n_527), .A2(n_57), .B1(n_58), .B2(n_61), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_524), .B(n_62), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_471), .B(n_64), .Y(n_592) );
XNOR2xp5_ASAP7_75t_L g593 ( .A(n_514), .B(n_67), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_474), .B(n_68), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_514), .A2(n_229), .B1(n_75), .B2(n_76), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_475), .B(n_72), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_520), .B(n_81), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_523), .A2(n_495), .B(n_475), .C(n_193), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_522), .A2(n_168), .B1(n_193), .B2(n_192), .C(n_184), .Y(n_599) );
OAI32xp33_ASAP7_75t_L g600 ( .A1(n_469), .A2(n_82), .A3(n_84), .B1(n_85), .B2(n_87), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_SL g601 ( .A1(n_510), .A2(n_192), .B(n_168), .C(n_89), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g602 ( .A1(n_472), .A2(n_166), .A3(n_173), .B1(n_174), .B2(n_184), .C1(n_229), .C2(n_510), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_488), .Y(n_603) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_516), .B(n_229), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_489), .B(n_229), .Y(n_605) );
XOR2x2_ASAP7_75t_L g606 ( .A(n_516), .B(n_229), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_477), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_477), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_510), .A2(n_166), .B(n_173), .C(n_174), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_538), .A2(n_539), .B1(n_543), .B2(n_547), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_551), .A2(n_545), .B(n_579), .C(n_550), .Y(n_611) );
AOI32xp33_ASAP7_75t_L g612 ( .A1(n_558), .A2(n_553), .A3(n_578), .B1(n_543), .B2(n_552), .Y(n_612) );
AOI21xp5_ASAP7_75t_SL g613 ( .A1(n_558), .A2(n_560), .B(n_536), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_530), .A2(n_544), .B1(n_535), .B2(n_551), .C(n_536), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_575), .B(n_549), .C(n_547), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_603), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_566), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_540), .A2(n_563), .B1(n_562), .B2(n_548), .C(n_572), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g619 ( .A1(n_530), .A2(n_535), .B1(n_542), .B2(n_537), .C(n_571), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_531), .A2(n_608), .B1(n_607), .B2(n_534), .C(n_533), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_546), .B(n_569), .Y(n_621) );
NAND4xp75_ASAP7_75t_L g622 ( .A(n_605), .B(n_556), .C(n_564), .D(n_557), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_602), .B(n_575), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_582), .A2(n_573), .B1(n_574), .B2(n_568), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_577), .B(n_593), .Y(n_626) );
AOI22x1_ASAP7_75t_SL g627 ( .A1(n_583), .A2(n_585), .B1(n_606), .B2(n_532), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_529), .B(n_554), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_560), .A2(n_609), .B(n_541), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_627), .A2(n_568), .B1(n_528), .B2(n_589), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_619), .A2(n_604), .B1(n_565), .B2(n_561), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_612), .A2(n_599), .B(n_576), .C(n_567), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_614), .A2(n_595), .B(n_581), .C(n_600), .Y(n_633) );
NOR2x1_ASAP7_75t_L g634 ( .A(n_613), .B(n_555), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_610), .A2(n_599), .B(n_555), .C(n_588), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_626), .A2(n_601), .B1(n_590), .B2(n_587), .C(n_584), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_611), .B(n_570), .C(n_597), .D(n_591), .Y(n_637) );
AOI31xp33_ASAP7_75t_L g638 ( .A1(n_624), .A2(n_598), .A3(n_559), .B(n_580), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_615), .A2(n_594), .B(n_592), .C(n_596), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_636), .B(n_629), .C(n_616), .Y(n_640) );
NOR3xp33_ASAP7_75t_SL g641 ( .A(n_632), .B(n_622), .C(n_618), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_634), .B(n_620), .C(n_628), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_638), .A2(n_621), .B(n_617), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_637), .B(n_625), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_631), .B(n_623), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_640), .A2(n_630), .B1(n_635), .B2(n_633), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_641), .A2(n_639), .B1(n_623), .B2(n_174), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_645), .B(n_623), .C(n_229), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_648), .Y(n_649) );
NOR3x1_ASAP7_75t_L g650 ( .A(n_647), .B(n_644), .C(n_642), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_646), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_649), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_651), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_652), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_653), .B(n_651), .Y(n_655) );
XNOR2x1_ASAP7_75t_L g656 ( .A(n_655), .B(n_650), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_654), .B(n_643), .Y(n_657) );
endmodule