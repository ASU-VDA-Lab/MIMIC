module fake_jpeg_27005_n_82 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx13_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_6),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_5),
.B1(n_10),
.B2(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_5),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_48),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B1(n_42),
.B2(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_75),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_28),
.C(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_30),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_35),
.C(n_60),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_77),
.A3(n_55),
.B1(n_40),
.B2(n_50),
.C1(n_61),
.C2(n_57),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_55),
.B(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_56),
.C(n_53),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_61),
.Y(n_82)
);


endmodule