module fake_jpeg_17166_n_143 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_43),
.B1(n_48),
.B2(n_34),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_66),
.B1(n_68),
.B2(n_2),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_45),
.B1(n_49),
.B2(n_37),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_44),
.B1(n_33),
.B2(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_74),
.Y(n_94)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_73),
.B1(n_59),
.B2(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_41),
.B(n_46),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_35),
.B(n_4),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_38),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_1),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_3),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_3),
.Y(n_113)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_83),
.B1(n_79),
.B2(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_110),
.B1(n_103),
.B2(n_95),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_77),
.C(n_78),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_94),
.B1(n_76),
.B2(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_116),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_112),
.B1(n_96),
.B2(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_99),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_99),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_111),
.Y(n_127)
);

INVxp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_105),
.C(n_108),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_123),
.B1(n_122),
.B2(n_124),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_125),
.B(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.Y(n_133)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_6),
.B(n_8),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_9),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_10),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_16),
.B(n_20),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_21),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_22),
.B(n_24),
.Y(n_143)
);


endmodule