module fake_jpeg_15119_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_9),
.B(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_1),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_51),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_41),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_48),
.B1(n_47),
.B2(n_43),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_65),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_48),
.B1(n_45),
.B2(n_49),
.Y(n_64)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_49),
.B1(n_45),
.B2(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_50),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_2),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_68),
.C(n_62),
.Y(n_90)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_62),
.B1(n_73),
.B2(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_96),
.B1(n_81),
.B2(n_87),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_94),
.B(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_74),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_16),
.B1(n_37),
.B2(n_36),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_13),
.B(n_33),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_103),
.B1(n_90),
.B2(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_75),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_81),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_95),
.C(n_91),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_96),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_108),
.B1(n_107),
.B2(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_11),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_10),
.B(n_38),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_28),
.B(n_23),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.C(n_86),
.Y(n_116)
);

AO221x1_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_117)
);

AOI31xp33_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_3),
.A3(n_7),
.B(n_8),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_8),
.Y(n_119)
);


endmodule