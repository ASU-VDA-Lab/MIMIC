module fake_ibex_649_n_2340 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2340);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2340;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_2183;
wire n_1859;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_2219;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_864;
wire n_608;
wire n_412;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_443;
wire n_1683;
wire n_436;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1941;
wire n_1707;
wire n_2064;
wire n_1679;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2251;
wire n_722;
wire n_2012;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_415;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_424;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_2337;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_924;
wire n_2331;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_566;
wire n_416;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_19),
.B(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_123),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_126),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_316),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_358),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

INVx4_ASAP7_75t_R g418 ( 
.A(n_313),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_343),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_190),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_48),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_387),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_336),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_4),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_2),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_3),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_205),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_18),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_321),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_153),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_164),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_291),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_325),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_299),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_44),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_259),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_266),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_84),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_172),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_288),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_314),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_72),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_394),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_108),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_363),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_302),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_65),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_250),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_295),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_85),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_233),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_285),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_376),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_335),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_89),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_60),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_258),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_362),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_12),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_212),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_2),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_399),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_146),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_1),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_353),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_115),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_319),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_377),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_76),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_46),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_214),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_402),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_315),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_232),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_33),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_142),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_307),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_298),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_263),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_300),
.Y(n_486)
);

BUFx5_ASAP7_75t_L g487 ( 
.A(n_251),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_225),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_368),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_365),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_107),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_310),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_84),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_346),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_158),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_229),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_222),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_345),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_227),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_72),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_5),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_111),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_328),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_284),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_53),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_158),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_391),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_367),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_224),
.Y(n_510)
);

INVxp33_ASAP7_75t_SL g511 ( 
.A(n_283),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_290),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_190),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_375),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_47),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_388),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_247),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_208),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_369),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_337),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_364),
.B(n_34),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_224),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_274),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_95),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_359),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_40),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_306),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_157),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_219),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_166),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_101),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_88),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_322),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_303),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_371),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_344),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_330),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_145),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_274),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_20),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_141),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_333),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_280),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_L g545 ( 
.A(n_338),
.B(n_329),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_392),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_357),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_177),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_114),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_59),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_204),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_13),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_265),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_106),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_127),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_311),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_45),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_203),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_334),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_386),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_31),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_326),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_1),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_222),
.Y(n_565)
);

CKINVDCx6p67_ASAP7_75t_R g566 ( 
.A(n_201),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_63),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_74),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_331),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_312),
.Y(n_570)
);

CKINVDCx14_ASAP7_75t_R g571 ( 
.A(n_188),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_233),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_28),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_372),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_354),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_7),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g577 ( 
.A(n_92),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_162),
.Y(n_578)
);

BUFx5_ASAP7_75t_L g579 ( 
.A(n_55),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_339),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_74),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_184),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_100),
.B(n_86),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_187),
.Y(n_584)
);

BUFx2_ASAP7_75t_SL g585 ( 
.A(n_155),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_297),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_209),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_246),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_173),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_348),
.B(n_151),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_305),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_201),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_378),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_157),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_218),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_176),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_144),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_106),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g599 ( 
.A(n_196),
.B(n_254),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_163),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_205),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_361),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_154),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_384),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_6),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_393),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_225),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_167),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_55),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_54),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_217),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_396),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_400),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_252),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_52),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_320),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_167),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_113),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_104),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_198),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_27),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_166),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_56),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_9),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_219),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_112),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_129),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_149),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_408),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_324),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_355),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_189),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_296),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_236),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_56),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_374),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_264),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_356),
.Y(n_638)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_120),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_294),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_397),
.Y(n_641)
);

BUFx2_ASAP7_75t_SL g642 ( 
.A(n_244),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_47),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_113),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_382),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_19),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_162),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_383),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_152),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_87),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_120),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_182),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_340),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_101),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_192),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_250),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_258),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_304),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_352),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_360),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_131),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_57),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_67),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_30),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_8),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_147),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_65),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_179),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_11),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_241),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_323),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_193),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_104),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_189),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_159),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_327),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_385),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_12),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_151),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_220),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_191),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_155),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_389),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_373),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_61),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_196),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_191),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_301),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_231),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_14),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_434),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_510),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_423),
.B(n_411),
.Y(n_693)
);

OAI22x1_ASAP7_75t_SL g694 ( 
.A1(n_421),
.A2(n_4),
.B1(n_0),
.B2(n_3),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_430),
.B(n_687),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_510),
.A2(n_6),
.B1(n_0),
.B2(n_5),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_429),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_429),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_487),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_429),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_423),
.B(n_410),
.Y(n_701)
);

OA21x2_ASAP7_75t_L g702 ( 
.A1(n_444),
.A2(n_281),
.B(n_279),
.Y(n_702)
);

AOI22x1_ASAP7_75t_SL g703 ( 
.A1(n_421),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_703)
);

INVx6_ASAP7_75t_L g704 ( 
.A(n_648),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_575),
.Y(n_705)
);

BUFx12f_ASAP7_75t_L g706 ( 
.A(n_434),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_527),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_527),
.B(n_10),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_429),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_435),
.B(n_15),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_496),
.B(n_15),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_487),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_562),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_571),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_434),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_648),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_507),
.B(n_16),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_571),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_507),
.B(n_21),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_426),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_479),
.B(n_282),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_515),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_437),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_487),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_SL g725 ( 
.A(n_425),
.B(n_407),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_624),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_489),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_672),
.B(n_22),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_548),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_428),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_447),
.B(n_25),
.Y(n_731)
);

INVx5_ASAP7_75t_L g732 ( 
.A(n_437),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_620),
.B(n_26),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_548),
.B(n_687),
.Y(n_734)
);

CKINVDCx6p67_ASAP7_75t_R g735 ( 
.A(n_648),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_487),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_493),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_588),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_558),
.A2(n_639),
.B1(n_577),
.B2(n_440),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_422),
.B(n_29),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_601),
.B(n_29),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_537),
.B(n_30),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_601),
.B(n_31),
.Y(n_743)
);

BUFx8_ASAP7_75t_SL g744 ( 
.A(n_454),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_521),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_449),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_444),
.B(n_32),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_487),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_490),
.A2(n_287),
.B(n_286),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_635),
.Y(n_750)
);

INVx6_ASAP7_75t_L g751 ( 
.A(n_579),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_416),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_635),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_427),
.B(n_33),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_663),
.Y(n_755)
);

BUFx12f_ASAP7_75t_L g756 ( 
.A(n_439),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_439),
.A2(n_540),
.B1(n_632),
.B2(n_440),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_420),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_540),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_431),
.B(n_34),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_490),
.B(n_35),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_453),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_579),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_449),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_455),
.Y(n_765)
);

OAI22x1_ASAP7_75t_SL g766 ( 
.A1(n_454),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_453),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_579),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_579),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_494),
.B(n_36),
.Y(n_770)
);

BUFx8_ASAP7_75t_SL g771 ( 
.A(n_498),
.Y(n_771)
);

OAI21x1_ASAP7_75t_L g772 ( 
.A1(n_504),
.A2(n_292),
.B(n_289),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_521),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_503),
.Y(n_774)
);

NOR2x1_ASAP7_75t_L g775 ( 
.A(n_517),
.B(n_293),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_SL g776 ( 
.A1(n_498),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_455),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_517),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_524),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_455),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_704),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_752),
.B(n_646),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_692),
.B(n_466),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_712),
.Y(n_784)
);

CKINVDCx6p67_ASAP7_75t_R g785 ( 
.A(n_691),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_724),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_736),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_704),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_696),
.B(n_714),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_695),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_711),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_748),
.B(n_505),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_763),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_768),
.B(n_505),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_769),
.Y(n_795)
);

INVx6_ASAP7_75t_L g796 ( 
.A(n_695),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_717),
.B(n_526),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_698),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_751),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_698),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_719),
.B(n_526),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_741),
.B(n_574),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_752),
.B(n_646),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_759),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_SL g805 ( 
.A(n_708),
.B(n_420),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_709),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_743),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_715),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_693),
.B(n_579),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_755),
.B(n_669),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_751),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_727),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_734),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_749),
.A2(n_417),
.B(n_415),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_723),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_716),
.B(n_511),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_726),
.B(n_713),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_726),
.B(n_466),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_713),
.B(n_566),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_715),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_753),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_738),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_705),
.B(n_419),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_745),
.B(n_773),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_566),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_746),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_762),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_757),
.B(n_413),
.Y(n_830)
);

BUFx4f_ASAP7_75t_L g831 ( 
.A(n_706),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_696),
.B(n_585),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_756),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_746),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_710),
.B(n_586),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_744),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_762),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_722),
.B(n_432),
.Y(n_838)
);

AND3x2_ASAP7_75t_L g839 ( 
.A(n_725),
.B(n_595),
.C(n_438),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_757),
.B(n_579),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_764),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_764),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_775),
.B(n_613),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_765),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_729),
.B(n_633),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_772),
.A2(n_660),
.B(n_633),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_765),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_701),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_777),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_750),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_701),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_728),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_777),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_701),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_725),
.B(n_660),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_780),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_731),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_742),
.B(n_671),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_780),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_721),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_697),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_697),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_742),
.B(n_671),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_697),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_700),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_771),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_702),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_700),
.Y(n_868)
);

NOR2x1p5_ASAP7_75t_L g869 ( 
.A(n_758),
.B(n_525),
.Y(n_869)
);

INVx8_ASAP7_75t_L g870 ( 
.A(n_721),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_700),
.Y(n_871)
);

AO22x2_ASAP7_75t_L g872 ( 
.A1(n_703),
.A2(n_714),
.B1(n_718),
.B2(n_737),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_767),
.B(n_436),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_732),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_732),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_732),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_739),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_702),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_721),
.Y(n_879)
);

OA22x2_ASAP7_75t_L g880 ( 
.A1(n_707),
.A2(n_441),
.B1(n_450),
.B2(n_433),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_774),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_778),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

AND2x4_ASAP7_75t_SL g884 ( 
.A(n_739),
.B(n_424),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_740),
.Y(n_885)
);

OR2x6_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_776),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_740),
.A2(n_456),
.B(n_443),
.Y(n_887)
);

NOR2x1p5_ASAP7_75t_L g888 ( 
.A(n_754),
.B(n_554),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_754),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_760),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_747),
.B(n_636),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_761),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_733),
.B(n_761),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_760),
.B(n_455),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_707),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_770),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_720),
.B(n_524),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_L g898 ( 
.A(n_720),
.B(n_534),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_730),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_730),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_737),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_776),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_694),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_766),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_692),
.B(n_636),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_704),
.B(n_457),
.Y(n_906)
);

AND3x2_ASAP7_75t_L g907 ( 
.A(n_759),
.B(n_468),
.C(n_459),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_695),
.B(n_559),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_SL g909 ( 
.A(n_708),
.B(n_424),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_776),
.A2(n_619),
.B1(n_622),
.B2(n_584),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_711),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_699),
.Y(n_912)
);

BUFx6f_ASAP7_75t_SL g913 ( 
.A(n_711),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_704),
.B(n_464),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_699),
.Y(n_915)
);

INVxp67_ASAP7_75t_R g916 ( 
.A(n_726),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_699),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_711),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_699),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_704),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_726),
.B(n_458),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_711),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_711),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_711),
.B(n_547),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_759),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_854),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_890),
.B(n_638),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_898),
.A2(n_499),
.B1(n_508),
.B2(n_461),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_790),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_885),
.B(n_640),
.Y(n_930)
);

NAND2x1_ASAP7_75t_L g931 ( 
.A(n_924),
.B(n_418),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_890),
.B(n_640),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_890),
.B(n_641),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_889),
.B(n_852),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_781),
.B(n_653),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_916),
.B(n_414),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_820),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_790),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_893),
.B(n_469),
.Y(n_939)
);

BUFx8_ASAP7_75t_L g940 ( 
.A(n_827),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_785),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_809),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_781),
.B(n_788),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_896),
.B(n_471),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_899),
.A2(n_499),
.B1(n_508),
.B2(n_461),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_815),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_896),
.B(n_477),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_796),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_796),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_920),
.B(n_509),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_883),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_891),
.B(n_446),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_883),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_898),
.A2(n_543),
.B1(n_591),
.B2(n_528),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_804),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_782),
.B(n_448),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_803),
.B(n_452),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_881),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_888),
.B(n_472),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_796),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_908),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_925),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_870),
.B(n_476),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_840),
.A2(n_543),
.B1(n_591),
.B2(n_528),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_783),
.B(n_483),
.Y(n_965)
);

OAI22xp33_ASAP7_75t_L g966 ( 
.A1(n_789),
.A2(n_584),
.B1(n_622),
.B2(n_619),
.Y(n_966)
);

INVx8_ASAP7_75t_L g967 ( 
.A(n_870),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_905),
.B(n_484),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_908),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_819),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_818),
.B(n_630),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_910),
.B(n_610),
.C(n_533),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_908),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_825),
.A2(n_475),
.B(n_506),
.C(n_478),
.Y(n_974)
);

BUFx5_ASAP7_75t_L g975 ( 
.A(n_848),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_791),
.B(n_486),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_808),
.B(n_631),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_821),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_921),
.B(n_857),
.Y(n_979)
);

NOR2x1p5_ASAP7_75t_L g980 ( 
.A(n_785),
.B(n_442),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_831),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_831),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_SL g983 ( 
.A(n_913),
.B(n_658),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_807),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_814),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_882),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_832),
.B(n_789),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_811),
.B(n_445),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_823),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_911),
.B(n_918),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_860),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_814),
.B(n_451),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_879),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_807),
.B(n_480),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_829),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_829),
.Y(n_996)
);

NOR2x1p5_ASAP7_75t_L g997 ( 
.A(n_836),
.B(n_460),
.Y(n_997)
);

AO221x1_ASAP7_75t_L g998 ( 
.A1(n_872),
.A2(n_676),
.B1(n_658),
.B2(n_668),
.C(n_551),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_829),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_822),
.B(n_516),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_807),
.B(n_492),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_814),
.B(n_462),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_923),
.B(n_495),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_923),
.B(n_922),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_833),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_899),
.A2(n_676),
.B1(n_668),
.B2(n_583),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_832),
.B(n_642),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_837),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_805),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_830),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_837),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_839),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_848),
.B(n_535),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_837),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_851),
.B(n_538),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_824),
.B(n_557),
.Y(n_1016)
);

INVx8_ASAP7_75t_L g1017 ( 
.A(n_870),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_851),
.B(n_580),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_850),
.B(n_593),
.Y(n_1019)
);

INVxp33_ASAP7_75t_L g1020 ( 
.A(n_906),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_833),
.B(n_590),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_909),
.Y(n_1022)
);

OR2x6_ASAP7_75t_SL g1023 ( 
.A(n_836),
.B(n_463),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_797),
.B(n_612),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_861),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_851),
.B(n_629),
.Y(n_1026)
);

NOR2x1p5_ASAP7_75t_L g1027 ( 
.A(n_866),
.B(n_465),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_835),
.B(n_512),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_801),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_802),
.B(n_858),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_810),
.B(n_470),
.C(n_467),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_802),
.B(n_514),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_884),
.B(n_473),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_900),
.A2(n_474),
.B1(n_482),
.B2(n_481),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_826),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_924),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_903),
.B(n_38),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_884),
.B(n_485),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_858),
.B(n_519),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_863),
.B(n_488),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_863),
.B(n_491),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_892),
.B(n_497),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_864),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_914),
.B(n_520),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_913),
.B(n_877),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_892),
.B(n_500),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_913),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_901),
.A2(n_549),
.B1(n_553),
.B2(n_541),
.C(n_531),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_892),
.B(n_544),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_902),
.B(n_682),
.C(n_502),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_845),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_855),
.B(n_887),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_845),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_897),
.B(n_501),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_873),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_792),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_838),
.B(n_550),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_816),
.B(n_560),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_843),
.B(n_513),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_867),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_799),
.B(n_518),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_865),
.Y(n_1062)
);

INVxp33_ASAP7_75t_L g1063 ( 
.A(n_900),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_L g1064 ( 
.A(n_902),
.B(n_895),
.C(n_904),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_792),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_799),
.B(n_523),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_868),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_813),
.B(n_530),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_813),
.B(n_532),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_794),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_897),
.B(n_561),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_816),
.B(n_563),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_904),
.B(n_39),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_794),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_868),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_866),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_907),
.B(n_569),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_880),
.B(n_539),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_894),
.B(n_570),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_919),
.B(n_542),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_784),
.B(n_606),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_784),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_880),
.B(n_552),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_862),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_871),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_846),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_786),
.B(n_556),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_871),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_787),
.B(n_616),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_875),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_875),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_L g1092 ( 
.A(n_867),
.B(n_565),
.C(n_564),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_789),
.B(n_832),
.Y(n_1093)
);

BUFx8_ASAP7_75t_L g1094 ( 
.A(n_872),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_876),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_832),
.B(n_573),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_869),
.B(n_599),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_872),
.B(n_589),
.C(n_576),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_793),
.B(n_645),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_793),
.B(n_677),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_795),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_795),
.B(n_683),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_912),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_886),
.B(n_592),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_912),
.B(n_684),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_878),
.B(n_688),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_886),
.B(n_598),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_SL g1108 ( 
.A(n_886),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_915),
.B(n_559),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_862),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_917),
.A2(n_568),
.B1(n_572),
.B2(n_567),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_874),
.B(n_667),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_874),
.B(n_690),
.Y(n_1113)
);

O2A1O1Ixp5_ASAP7_75t_L g1114 ( 
.A1(n_798),
.A2(n_522),
.B(n_690),
.C(n_679),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_812),
.Y(n_1115)
);

BUFx5_ASAP7_75t_L g1116 ( 
.A(n_812),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_R g1117 ( 
.A(n_985),
.B(n_958),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_934),
.B(n_600),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_978),
.B(n_603),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_934),
.B(n_605),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_987),
.A2(n_582),
.B1(n_587),
.B2(n_578),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1112),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1036),
.B(n_608),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1010),
.B(n_970),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_SL g1125 ( 
.A(n_967),
.B(n_545),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1086),
.A2(n_806),
.B(n_800),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_R g1127 ( 
.A(n_941),
.B(n_615),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1036),
.B(n_679),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_986),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1112),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_927),
.B(n_932),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1113),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_927),
.B(n_617),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_987),
.B(n_594),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_L g1135 ( 
.A(n_945),
.B(n_966),
.C(n_1006),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_932),
.B(n_618),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1058),
.A2(n_412),
.B(n_596),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_933),
.B(n_621),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_933),
.B(n_626),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_967),
.B(n_547),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1058),
.A2(n_607),
.B(n_597),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_926),
.B(n_627),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_974),
.A2(n_611),
.B(n_614),
.C(n_609),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_955),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1113),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_930),
.B(n_628),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_945),
.B(n_649),
.Y(n_1147)
);

BUFx2_ASAP7_75t_R g1148 ( 
.A(n_1023),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_987),
.A2(n_643),
.B1(n_644),
.B2(n_637),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_962),
.B(n_656),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_984),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_982),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_951),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1072),
.A2(n_650),
.B(n_647),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1106),
.A2(n_654),
.B(n_655),
.C(n_651),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1055),
.B(n_657),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_967),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1017),
.B(n_659),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1020),
.B(n_662),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_988),
.B(n_673),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_979),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_1017),
.B(n_659),
.Y(n_1162)
);

CKINVDCx8_ASAP7_75t_R g1163 ( 
.A(n_1076),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1004),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1035),
.B(n_678),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1045),
.B(n_661),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1029),
.B(n_664),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_953),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1064),
.A2(n_666),
.B1(n_670),
.B2(n_665),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_939),
.A2(n_675),
.B(n_680),
.C(n_674),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1004),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1054),
.A2(n_685),
.B1(n_686),
.B2(n_681),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_936),
.B(n_689),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_940),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1007),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1030),
.B(n_529),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1030),
.B(n_551),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_990),
.B(n_555),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_939),
.B(n_937),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_964),
.B(n_40),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1017),
.Y(n_1181)
);

BUFx4f_ASAP7_75t_L g1182 ( 
.A(n_1007),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1114),
.A2(n_623),
.B(n_625),
.C(n_581),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_944),
.A2(n_834),
.B(n_828),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_992),
.B(n_581),
.Y(n_1185)
);

NOR2xp67_ASAP7_75t_L g1186 ( 
.A(n_981),
.B(n_41),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_944),
.A2(n_842),
.B(n_841),
.Y(n_1187)
);

CKINVDCx6p67_ASAP7_75t_R g1188 ( 
.A(n_1005),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1093),
.A2(n_625),
.B1(n_634),
.B2(n_623),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1002),
.B(n_623),
.Y(n_1190)
);

OAI21xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1007),
.A2(n_41),
.B(n_42),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1009),
.B(n_1022),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_947),
.A2(n_842),
.B(n_841),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_947),
.A2(n_847),
.B(n_844),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_940),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_928),
.A2(n_634),
.B1(n_652),
.B2(n_625),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1098),
.A2(n_652),
.B1(n_634),
.B2(n_546),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1079),
.A2(n_652),
.B(n_634),
.C(n_546),
.Y(n_1198)
);

BUFx4f_ASAP7_75t_L g1199 ( 
.A(n_1012),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1039),
.A2(n_652),
.B(n_546),
.C(n_602),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_942),
.B(n_42),
.Y(n_1201)
);

BUFx4f_ASAP7_75t_L g1202 ( 
.A(n_1097),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_946),
.B(n_43),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_961),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_969),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1107),
.B(n_43),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_973),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_983),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1032),
.B(n_44),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_954),
.A2(n_546),
.B1(n_602),
.B2(n_536),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1032),
.B(n_1071),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1039),
.A2(n_602),
.B1(n_604),
.B2(n_536),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1085),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1033),
.B(n_46),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1040),
.B(n_48),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1047),
.B(n_49),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1084),
.Y(n_1217)
);

AO21x1_ASAP7_75t_L g1218 ( 
.A1(n_1049),
.A2(n_853),
.B(n_849),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_994),
.A2(n_1003),
.B(n_1001),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_994),
.A2(n_859),
.B(n_856),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1038),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1041),
.B(n_49),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1057),
.B(n_50),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1057),
.B(n_50),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_968),
.B(n_51),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_989),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1044),
.B(n_51),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1034),
.B(n_52),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_929),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1104),
.B(n_53),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_L g1231 ( 
.A(n_1097),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1001),
.A2(n_859),
.B(n_856),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1111),
.A2(n_58),
.B(n_54),
.C(n_57),
.Y(n_1233)
);

CKINVDCx6p67_ASAP7_75t_R g1234 ( 
.A(n_1108),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1082),
.B(n_59),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_817),
.B1(n_63),
.B2(n_60),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1078),
.B(n_62),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_938),
.B(n_62),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_948),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_949),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1111),
.A2(n_67),
.B(n_64),
.C(n_66),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1028),
.B(n_66),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_980),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1028),
.B(n_1080),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1084),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_960),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1101),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1056),
.A2(n_71),
.B(n_68),
.C(n_70),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1096),
.B(n_71),
.Y(n_1249)
);

NOR2x1_ASAP7_75t_R g1250 ( 
.A(n_998),
.B(n_1083),
.Y(n_1250)
);

NOR2x1p5_ASAP7_75t_L g1251 ( 
.A(n_931),
.B(n_73),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1025),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1087),
.B(n_73),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1021),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_959),
.B(n_75),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_971),
.B(n_75),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1073),
.B(n_76),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_965),
.B(n_77),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_952),
.B(n_77),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1065),
.A2(n_1074),
.B(n_1070),
.Y(n_1260)
);

NAND2x1p5_ASAP7_75t_L g1261 ( 
.A(n_991),
.B(n_78),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_935),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_956),
.B(n_79),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1099),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1264)
);

OAI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1024),
.A2(n_80),
.B(n_81),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1109),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_991),
.B(n_82),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_957),
.B(n_82),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1048),
.B(n_83),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1059),
.B(n_83),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1031),
.A2(n_309),
.B(n_308),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1103),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_977),
.B(n_943),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1092),
.A2(n_318),
.B(n_317),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1049),
.A2(n_90),
.B(n_91),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_976),
.B(n_90),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1037),
.B(n_91),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_995),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_972),
.B(n_93),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1043),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1042),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1051),
.B(n_1053),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_950),
.B(n_94),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1050),
.B(n_94),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1099),
.A2(n_342),
.B(n_341),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_997),
.B(n_1027),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1061),
.B(n_95),
.Y(n_1287)
);

BUFx8_ASAP7_75t_L g1288 ( 
.A(n_1108),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_996),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_993),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_L g1291 ( 
.A(n_999),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1102),
.A2(n_349),
.B(n_347),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1008),
.Y(n_1293)
);

AOI33xp33_ASAP7_75t_L g1294 ( 
.A1(n_1011),
.A2(n_96),
.A3(n_97),
.B1(n_98),
.B2(n_99),
.B3(n_100),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1102),
.A2(n_351),
.B(n_350),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1046),
.B(n_98),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1000),
.B(n_99),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1014),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1016),
.B(n_102),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1066),
.B(n_1068),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1077),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1019),
.B(n_105),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1088),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1090),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1081),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1089),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1306)
);

NOR3xp33_ASAP7_75t_L g1307 ( 
.A(n_1069),
.B(n_110),
.C(n_111),
.Y(n_1307)
);

BUFx8_ASAP7_75t_L g1308 ( 
.A(n_1062),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1100),
.B(n_110),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1105),
.B(n_114),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_963),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1013),
.B(n_117),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1091),
.B(n_118),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1060),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1095),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1015),
.B(n_124),
.Y(n_1317)
);

BUFx4f_ASAP7_75t_L g1318 ( 
.A(n_1110),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1018),
.B(n_124),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1115),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1116),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1026),
.B(n_125),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1094),
.B(n_127),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_975),
.A2(n_128),
.B(n_129),
.C(n_130),
.Y(n_1324)
);

INVx4_ASAP7_75t_L g1325 ( 
.A(n_975),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1116),
.B(n_128),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1094),
.A2(n_380),
.B(n_379),
.Y(n_1327)
);

NAND3x1_ASAP7_75t_L g1328 ( 
.A(n_1148),
.B(n_132),
.C(n_133),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1164),
.B(n_133),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1226),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1171),
.B(n_134),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_SL g1332 ( 
.A1(n_1327),
.A2(n_134),
.B(n_135),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1161),
.B(n_135),
.Y(n_1333)
);

BUFx4f_ASAP7_75t_SL g1334 ( 
.A(n_1308),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1179),
.B(n_136),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1176),
.A2(n_1177),
.B(n_1244),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1188),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1273),
.B(n_136),
.C(n_137),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1182),
.B(n_137),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1126),
.A2(n_1183),
.B(n_1184),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1308),
.Y(n_1341)
);

CKINVDCx9p33_ASAP7_75t_R g1342 ( 
.A(n_1124),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1122),
.B(n_138),
.Y(n_1343)
);

AND3x4_ASAP7_75t_L g1344 ( 
.A(n_1135),
.B(n_138),
.C(n_139),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1191),
.A2(n_139),
.B(n_140),
.C(n_142),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1144),
.Y(n_1346)
);

AOI21xp33_ASAP7_75t_L g1347 ( 
.A1(n_1159),
.A2(n_140),
.B(n_143),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1216),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1275),
.A2(n_143),
.A3(n_144),
.B(n_146),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1218),
.A2(n_147),
.A3(n_148),
.B(n_149),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1153),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1168),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1147),
.B(n_148),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1130),
.B(n_150),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1132),
.A2(n_405),
.B(n_403),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1321),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1145),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1118),
.B(n_154),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1197),
.B(n_1166),
.C(n_1307),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1120),
.B(n_156),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1195),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1303),
.A2(n_1266),
.B1(n_1182),
.B2(n_1154),
.Y(n_1362)
);

NAND3x1_ASAP7_75t_L g1363 ( 
.A(n_1323),
.B(n_160),
.C(n_161),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1216),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1212),
.A2(n_165),
.A3(n_168),
.B(n_169),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1172),
.B(n_168),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1260),
.A2(n_169),
.B(n_170),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1303),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1211),
.B(n_173),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1173),
.B(n_174),
.Y(n_1370)
);

AOI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1119),
.A2(n_174),
.B(n_175),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1221),
.B(n_175),
.Y(n_1372)
);

NAND2x1_ASAP7_75t_L g1373 ( 
.A(n_1217),
.B(n_176),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1121),
.B(n_178),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1217),
.B(n_179),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1141),
.A2(n_1154),
.B(n_1282),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1180),
.B(n_180),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1141),
.A2(n_180),
.B(n_181),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1327),
.A2(n_183),
.B(n_185),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1150),
.B(n_185),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1157),
.B(n_186),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1137),
.A2(n_186),
.B(n_187),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1201),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1203),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1206),
.B(n_1134),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1134),
.B(n_194),
.Y(n_1386)
);

INVx6_ASAP7_75t_SL g1387 ( 
.A(n_1277),
.Y(n_1387)
);

AOI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1250),
.A2(n_195),
.B(n_197),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1155),
.B(n_1214),
.Y(n_1389)
);

AOI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1143),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.C(n_200),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1169),
.B(n_202),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1170),
.B(n_203),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1149),
.A2(n_1262),
.B1(n_1235),
.B2(n_1230),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1229),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1165),
.B(n_206),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1304),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1185),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1269),
.B(n_207),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1149),
.B(n_1249),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1133),
.B(n_209),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1136),
.B(n_210),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1140),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1174),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1160),
.B(n_211),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1138),
.B(n_212),
.Y(n_1405)
);

OAI21xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1251),
.A2(n_213),
.B(n_214),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1300),
.B(n_213),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1204),
.B(n_215),
.Y(n_1408)
);

BUFx8_ASAP7_75t_L g1409 ( 
.A(n_1286),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1156),
.B(n_1192),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1259),
.A2(n_1268),
.B(n_1263),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1223),
.A2(n_216),
.B1(n_218),
.B2(n_220),
.Y(n_1412)
);

AND3x4_ASAP7_75t_L g1413 ( 
.A(n_1152),
.B(n_221),
.C(n_223),
.Y(n_1413)
);

AND2x6_ASAP7_75t_SL g1414 ( 
.A(n_1163),
.B(n_221),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1140),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1279),
.B(n_226),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1224),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_1128),
.Y(n_1418)
);

AOI221x1_ASAP7_75t_L g1419 ( 
.A1(n_1265),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.C(n_232),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1205),
.B(n_234),
.Y(n_1420)
);

OAI22x1_ASAP7_75t_L g1421 ( 
.A1(n_1257),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1196),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1140),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1146),
.B(n_239),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1190),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1234),
.B(n_240),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1207),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1129),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1225),
.B(n_242),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1285),
.A2(n_242),
.B(n_243),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1287),
.B(n_243),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1287),
.B(n_245),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1215),
.A2(n_248),
.B(n_249),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1258),
.B(n_251),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1178),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1233),
.A2(n_252),
.B(n_253),
.C(n_255),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1278),
.A2(n_253),
.B(n_255),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1202),
.B(n_256),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1199),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1289),
.Y(n_1440)
);

OAI22x1_ASAP7_75t_L g1441 ( 
.A1(n_1257),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1175),
.B(n_257),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1222),
.A2(n_262),
.B(n_263),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1167),
.B(n_1237),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1293),
.A2(n_262),
.B(n_264),
.Y(n_1445)
);

INVx6_ASAP7_75t_SL g1446 ( 
.A(n_1277),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1128),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1298),
.A2(n_1313),
.B(n_1242),
.Y(n_1448)
);

OAI321xp33_ASAP7_75t_L g1449 ( 
.A1(n_1196),
.A2(n_267),
.A3(n_268),
.B1(n_269),
.B2(n_270),
.C(n_271),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1213),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1228),
.B(n_269),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1181),
.B(n_272),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1187),
.A2(n_1194),
.B(n_1193),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_SL g1454 ( 
.A(n_1301),
.B(n_273),
.C(n_275),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1227),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1321),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1238),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1253),
.A2(n_276),
.B(n_277),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1139),
.B(n_278),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1252),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1281),
.B(n_278),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1321),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1255),
.B(n_1284),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1245),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1299),
.B(n_1209),
.Y(n_1465)
);

AOI21xp33_ASAP7_75t_L g1466 ( 
.A1(n_1254),
.A2(n_1256),
.B(n_1297),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1208),
.B(n_1243),
.Y(n_1467)
);

O2A1O1Ixp5_ASAP7_75t_L g1468 ( 
.A1(n_1326),
.A2(n_1274),
.B(n_1271),
.C(n_1296),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1220),
.A2(n_1232),
.B(n_1270),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1202),
.B(n_1231),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1240),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1151),
.B(n_1246),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1280),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1210),
.A2(n_1283),
.B1(n_1231),
.B2(n_1319),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1305),
.B(n_1276),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1200),
.A2(n_1198),
.A3(n_1236),
.B(n_1189),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1241),
.A2(n_1294),
.B(n_1311),
.C(n_1264),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_SL g1478 ( 
.A(n_1316),
.B(n_1162),
.C(n_1158),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1302),
.B(n_1312),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1199),
.B(n_1291),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1239),
.B(n_1142),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1314),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1309),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1325),
.B(n_1123),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1291),
.B(n_1318),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1310),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_SL g1487 ( 
.A(n_1127),
.B(n_1288),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1288),
.Y(n_1488)
);

BUFx10_ASAP7_75t_L g1489 ( 
.A(n_1317),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1210),
.B(n_1322),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1290),
.Y(n_1491)
);

AO31x2_ASAP7_75t_L g1492 ( 
.A1(n_1236),
.A2(n_1324),
.A3(n_1248),
.B(n_1247),
.Y(n_1492)
);

INVx5_ASAP7_75t_L g1493 ( 
.A(n_1320),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1272),
.A2(n_1306),
.A3(n_1267),
.B(n_1261),
.Y(n_1494)
);

NOR2x1_ASAP7_75t_SL g1495 ( 
.A(n_1306),
.B(n_1320),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1320),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1117),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1158),
.A2(n_1162),
.B1(n_1125),
.B2(n_1186),
.Y(n_1498)
);

INVx4_ASAP7_75t_L g1499 ( 
.A(n_1318),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1164),
.B(n_934),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1226),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1226),
.Y(n_1502)
);

AO31x2_ASAP7_75t_L g1503 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1164),
.B(n_934),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1153),
.Y(n_1505)
);

BUFx12f_ASAP7_75t_L g1506 ( 
.A(n_1174),
.Y(n_1506)
);

INVx8_ASAP7_75t_L g1507 ( 
.A(n_1140),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1308),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1164),
.B(n_934),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1164),
.B(n_934),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1308),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_L g1512 ( 
.A(n_1174),
.Y(n_1512)
);

AO31x2_ASAP7_75t_L g1513 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1183),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1219),
.A2(n_1052),
.B(n_1131),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1226),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1175),
.B(n_987),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1161),
.B(n_970),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1161),
.B(n_970),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1164),
.B(n_934),
.Y(n_1520)
);

AO21x2_ASAP7_75t_L g1521 ( 
.A1(n_1137),
.A2(n_1183),
.B(n_1072),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1219),
.A2(n_1052),
.B(n_1131),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1183),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1191),
.C(n_1233),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1164),
.B(n_934),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1179),
.B(n_1093),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1217),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1164),
.B(n_934),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1217),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1161),
.B(n_970),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1164),
.B(n_934),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1183),
.Y(n_1532)
);

AO31x2_ASAP7_75t_L g1533 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1161),
.B(n_945),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1161),
.B(n_970),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1308),
.Y(n_1536)
);

AO21x1_ASAP7_75t_L g1537 ( 
.A1(n_1285),
.A2(n_1295),
.B(n_1292),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1174),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1195),
.B(n_945),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1161),
.B(n_970),
.Y(n_1540)
);

AO31x2_ASAP7_75t_L g1541 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1217),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1161),
.B(n_970),
.Y(n_1543)
);

OAI22x1_ASAP7_75t_L g1544 ( 
.A1(n_1216),
.A2(n_964),
.B1(n_758),
.B2(n_954),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1183),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_SL g1546 ( 
.A(n_1148),
.B(n_945),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1164),
.B(n_934),
.Y(n_1547)
);

AO31x2_ASAP7_75t_L g1548 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1164),
.B(n_934),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1164),
.B(n_934),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1174),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1188),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1164),
.B(n_934),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1164),
.B(n_934),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1226),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1164),
.B(n_934),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1315),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1175),
.B(n_987),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1195),
.B(n_945),
.Y(n_1559)
);

A2O1A1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1191),
.C(n_1233),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1183),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1153),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1153),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1308),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1308),
.Y(n_1565)
);

AO31x2_ASAP7_75t_L g1566 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1566)
);

AOI21xp33_ASAP7_75t_L g1567 ( 
.A1(n_1159),
.A2(n_1063),
.B(n_1045),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1174),
.Y(n_1568)
);

AOI21xp33_ASAP7_75t_L g1569 ( 
.A1(n_1159),
.A2(n_1063),
.B(n_1045),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1179),
.B(n_1093),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1308),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1315),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1191),
.C(n_1233),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1161),
.B(n_970),
.Y(n_1574)
);

AO31x2_ASAP7_75t_L g1575 ( 
.A1(n_1275),
.A2(n_1183),
.A3(n_1218),
.B(n_1072),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1411),
.A2(n_1336),
.B(n_1537),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1500),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1340),
.A2(n_1469),
.B(n_1453),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1504),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1511),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1524),
.A2(n_1573),
.B(n_1560),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1338),
.B(n_1436),
.C(n_1466),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1351),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1520),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1525),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1334),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1507),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1334),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1528),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1436),
.B(n_1419),
.C(n_1345),
.Y(n_1591)
);

INVx3_ASAP7_75t_SL g1592 ( 
.A(n_1571),
.Y(n_1592)
);

BUFx2_ASAP7_75t_SL g1593 ( 
.A(n_1341),
.Y(n_1593)
);

NOR2xp67_ASAP7_75t_L g1594 ( 
.A(n_1536),
.B(n_1511),
.Y(n_1594)
);

BUFx4_ASAP7_75t_SL g1595 ( 
.A(n_1341),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1507),
.B(n_1571),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1357),
.B(n_1531),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1508),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1564),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1547),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1508),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1549),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1357),
.B(n_1550),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1352),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1518),
.B(n_1519),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1507),
.B(n_1571),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1553),
.Y(n_1607)
);

INVx5_ASAP7_75t_L g1608 ( 
.A(n_1415),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1493),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_SL g1610 ( 
.A(n_1415),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1493),
.Y(n_1611)
);

INVx4_ASAP7_75t_L g1612 ( 
.A(n_1493),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1336),
.A2(n_1523),
.B(n_1514),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1460),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1554),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1556),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1402),
.B(n_1423),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1330),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1565),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1530),
.B(n_1535),
.Y(n_1620)
);

BUFx2_ASAP7_75t_SL g1621 ( 
.A(n_1403),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1534),
.B(n_1526),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1526),
.B(n_1570),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1532),
.A2(n_1561),
.B(n_1545),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1540),
.B(n_1543),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1460),
.Y(n_1626)
);

INVx6_ASAP7_75t_L g1627 ( 
.A(n_1409),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1356),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1501),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1399),
.A2(n_1393),
.B1(n_1407),
.B2(n_1362),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_SL g1631 ( 
.A1(n_1332),
.A2(n_1495),
.B(n_1378),
.Y(n_1631)
);

BUFx4f_ASAP7_75t_SL g1632 ( 
.A(n_1506),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1345),
.B(n_1569),
.C(n_1567),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1502),
.Y(n_1634)
);

NAND2x1p5_ASAP7_75t_L g1635 ( 
.A(n_1499),
.B(n_1456),
.Y(n_1635)
);

BUFx2_ASAP7_75t_SL g1636 ( 
.A(n_1403),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1452),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1570),
.B(n_1410),
.Y(n_1638)
);

INVx4_ASAP7_75t_L g1639 ( 
.A(n_1456),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_SL g1640 ( 
.A1(n_1437),
.A2(n_1445),
.B(n_1367),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1473),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1346),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1524),
.A2(n_1573),
.B(n_1560),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1410),
.B(n_1463),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1473),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1516),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1488),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1462),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1450),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1521),
.A2(n_1522),
.B(n_1515),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1555),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1385),
.B(n_1348),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1376),
.A2(n_1477),
.B(n_1406),
.C(n_1407),
.Y(n_1653)
);

INVx6_ASAP7_75t_L g1654 ( 
.A(n_1409),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1505),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1505),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1546),
.A2(n_1344),
.B1(n_1544),
.B2(n_1574),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1387),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1394),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1396),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_SL g1661 ( 
.A1(n_1498),
.A2(n_1355),
.B(n_1430),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1387),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1377),
.B(n_1364),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1427),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1539),
.B(n_1559),
.Y(n_1665)
);

INVx3_ASAP7_75t_SL g1666 ( 
.A(n_1538),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1517),
.B(n_1558),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1471),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1375),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1539),
.B(n_1559),
.Y(n_1670)
);

INVx6_ASAP7_75t_L g1671 ( 
.A(n_1506),
.Y(n_1671)
);

CKINVDCx16_ASAP7_75t_R g1672 ( 
.A(n_1487),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1527),
.Y(n_1673)
);

AO21x2_ASAP7_75t_L g1674 ( 
.A1(n_1478),
.A2(n_1448),
.B(n_1490),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1375),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1389),
.B(n_1353),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1413),
.A2(n_1539),
.B1(n_1559),
.B2(n_1344),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1474),
.A2(n_1446),
.B1(n_1465),
.B2(n_1331),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1359),
.A2(n_1468),
.B(n_1424),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1360),
.B(n_1333),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1517),
.B(n_1558),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1372),
.B(n_1438),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1446),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1383),
.B(n_1384),
.Y(n_1684)
);

INVx4_ASAP7_75t_L g1685 ( 
.A(n_1529),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1413),
.A2(n_1452),
.B1(n_1416),
.B2(n_1424),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1404),
.B(n_1482),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1529),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1440),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1337),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1552),
.B(n_1461),
.Y(n_1691)
);

NOR2xp67_ASAP7_75t_SL g1692 ( 
.A(n_1512),
.B(n_1551),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1444),
.A2(n_1435),
.B(n_1475),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1479),
.B(n_1483),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1342),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1398),
.A2(n_1358),
.B(n_1329),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1440),
.B(n_1480),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1464),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1395),
.B(n_1366),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1418),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1339),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1433),
.A2(n_1443),
.B(n_1458),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1342),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1454),
.A2(n_1390),
.B1(n_1392),
.B2(n_1370),
.Y(n_1704)
);

INVx3_ASAP7_75t_SL g1705 ( 
.A(n_1568),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1562),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1439),
.B(n_1361),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1499),
.B(n_1542),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1485),
.B(n_1486),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1464),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1491),
.Y(n_1711)
);

AND2x4_ASAP7_75t_SL g1712 ( 
.A(n_1470),
.B(n_1496),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1339),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1408),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1381),
.A2(n_1354),
.B(n_1343),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_SL g1716 ( 
.A1(n_1491),
.A2(n_1432),
.B(n_1431),
.Y(n_1716)
);

AO31x2_ASAP7_75t_L g1717 ( 
.A1(n_1447),
.A2(n_1412),
.A3(n_1417),
.B(n_1455),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1380),
.B(n_1457),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1381),
.A2(n_1373),
.B(n_1420),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1335),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1414),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1369),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1421),
.Y(n_1723)
);

BUFx12f_ASAP7_75t_L g1724 ( 
.A(n_1426),
.Y(n_1724)
);

INVx11_ASAP7_75t_L g1725 ( 
.A(n_1328),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1451),
.A2(n_1429),
.B(n_1434),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_L g1727 ( 
.A(n_1390),
.B(n_1388),
.C(n_1347),
.Y(n_1727)
);

INVx6_ASAP7_75t_L g1728 ( 
.A(n_1489),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1489),
.B(n_1405),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1441),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1497),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1442),
.Y(n_1732)
);

OA21x2_ASAP7_75t_L g1733 ( 
.A1(n_1400),
.A2(n_1401),
.B(n_1449),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1371),
.A2(n_1422),
.B(n_1563),
.Y(n_1734)
);

AO21x2_ASAP7_75t_L g1735 ( 
.A1(n_1382),
.A2(n_1379),
.B(n_1386),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1397),
.A2(n_1425),
.B(n_1459),
.Y(n_1736)
);

O2A1O1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1391),
.A2(n_1374),
.B(n_1368),
.C(n_1481),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1428),
.A2(n_1575),
.B(n_1503),
.Y(n_1738)
);

AO21x2_ASAP7_75t_L g1739 ( 
.A1(n_1503),
.A2(n_1575),
.B(n_1513),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1503),
.A2(n_1541),
.B(n_1566),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1472),
.B(n_1481),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1513),
.A2(n_1548),
.B(n_1533),
.Y(n_1742)
);

AOI22x1_ASAP7_75t_L g1743 ( 
.A1(n_1484),
.A2(n_1572),
.B1(n_1557),
.B2(n_1472),
.Y(n_1743)
);

OAI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1513),
.A2(n_1566),
.B(n_1548),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1467),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1533),
.A2(n_1566),
.B(n_1548),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1533),
.A2(n_1566),
.B(n_1548),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1363),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1533),
.A2(n_1541),
.B(n_1557),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1492),
.A2(n_1349),
.B1(n_1494),
.B2(n_1365),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1541),
.A2(n_1350),
.B(n_1494),
.Y(n_1751)
);

OAI21x1_ASAP7_75t_L g1752 ( 
.A1(n_1541),
.A2(n_1350),
.B(n_1476),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1350),
.A2(n_1476),
.B(n_1492),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1476),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1365),
.B(n_1350),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1524),
.A2(n_1573),
.B(n_1560),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1334),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1500),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1518),
.B(n_852),
.Y(n_1759)
);

NAND2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1415),
.B(n_1182),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_SL g1761 ( 
.A(n_1415),
.B(n_1500),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1334),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1500),
.A2(n_945),
.B1(n_1135),
.B2(n_758),
.Y(n_1763)
);

NAND2x1p5_ASAP7_75t_L g1764 ( 
.A(n_1415),
.B(n_1182),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1500),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1500),
.B(n_1504),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1334),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1618),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1629),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1634),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1677),
.A2(n_1638),
.B1(n_1622),
.B2(n_1630),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1598),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1646),
.Y(n_1773)
);

BUFx8_ASAP7_75t_L g1774 ( 
.A(n_1589),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1584),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1608),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1598),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1759),
.B(n_1605),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1620),
.B(n_1625),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1642),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1584),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1651),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1612),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1686),
.A2(n_1597),
.B1(n_1603),
.B2(n_1637),
.Y(n_1784)
);

OAI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1644),
.A2(n_1638),
.B(n_1750),
.Y(n_1785)
);

INVxp33_ASAP7_75t_L g1786 ( 
.A(n_1581),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1659),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1597),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1612),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1604),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1660),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1597),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1664),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1668),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1614),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1587),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1684),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1727),
.A2(n_1583),
.B(n_1633),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1587),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1626),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1577),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1579),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1622),
.A2(n_1644),
.B1(n_1603),
.B2(n_1723),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1585),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1626),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1603),
.B(n_1766),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1641),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1608),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1586),
.Y(n_1809)
);

INVx4_ASAP7_75t_SL g1810 ( 
.A(n_1627),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1590),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1645),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1655),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1655),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1656),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1656),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1608),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1600),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1767),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1602),
.Y(n_1820)
);

BUFx2_ASAP7_75t_R g1821 ( 
.A(n_1757),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1619),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1639),
.B(n_1689),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1607),
.Y(n_1824)
);

AO21x2_ASAP7_75t_L g1825 ( 
.A1(n_1576),
.A2(n_1613),
.B(n_1661),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1713),
.A2(n_1748),
.B1(n_1637),
.B2(n_1678),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1615),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1616),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1623),
.A2(n_1657),
.B1(n_1763),
.B2(n_1704),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1758),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1767),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1765),
.B(n_1682),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1593),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1730),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1665),
.A2(n_1670),
.B1(n_1704),
.B2(n_1722),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1741),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1663),
.B(n_1697),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1706),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1706),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1649),
.B(n_1619),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1580),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1595),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1694),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1694),
.Y(n_1844)
);

INVx4_ASAP7_75t_L g1845 ( 
.A(n_1608),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1701),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1589),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1601),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1676),
.B(n_1687),
.Y(n_1849)
);

BUFx4f_ASAP7_75t_SL g1850 ( 
.A(n_1647),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1687),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1718),
.B(n_1599),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1639),
.B(n_1761),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1594),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1757),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1699),
.B(n_1680),
.Y(n_1856)
);

OR2x6_ASAP7_75t_L g1857 ( 
.A(n_1588),
.B(n_1596),
.Y(n_1857)
);

INVx6_ASAP7_75t_L g1858 ( 
.A(n_1639),
.Y(n_1858)
);

INVx6_ASAP7_75t_L g1859 ( 
.A(n_1627),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1669),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1675),
.Y(n_1861)
);

INVx6_ASAP7_75t_L g1862 ( 
.A(n_1627),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1731),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1697),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1712),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1709),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1665),
.A2(n_1670),
.B1(n_1720),
.B2(n_1640),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1714),
.A2(n_1591),
.B1(n_1754),
.B2(n_1696),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1695),
.B(n_1703),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1754),
.A2(n_1729),
.B1(n_1643),
.B2(n_1582),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1578),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1652),
.B(n_1681),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1700),
.A2(n_1617),
.B1(n_1693),
.B2(n_1653),
.Y(n_1873)
);

OAI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1672),
.A2(n_1606),
.B1(n_1596),
.B2(n_1685),
.Y(n_1874)
);

CKINVDCx8_ASAP7_75t_R g1875 ( 
.A(n_1762),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1729),
.A2(n_1756),
.B1(n_1732),
.B2(n_1679),
.Y(n_1876)
);

BUFx8_ASAP7_75t_L g1877 ( 
.A(n_1658),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1588),
.Y(n_1878)
);

CKINVDCx11_ASAP7_75t_R g1879 ( 
.A(n_1647),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1712),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1628),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1628),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1652),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1681),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1609),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1736),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1617),
.A2(n_1631),
.B1(n_1654),
.B2(n_1636),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1762),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1588),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1691),
.B(n_1690),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1596),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1592),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1609),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1606),
.Y(n_1894)
);

INVxp33_ASAP7_75t_L g1895 ( 
.A(n_1635),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1592),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1621),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1650),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1606),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1760),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1667),
.B(n_1745),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1708),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1654),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1708),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1650),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1711),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1755),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1632),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1611),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1745),
.B(n_1611),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1648),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1632),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1673),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1635),
.B(n_1673),
.Y(n_1914)
);

NOR2x1_ASAP7_75t_L g1915 ( 
.A(n_1892),
.B(n_1711),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1823),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1871),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1801),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1853),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1823),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1843),
.B(n_1653),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1907),
.B(n_1751),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1802),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1804),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1858),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1844),
.B(n_1737),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1838),
.B(n_1753),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1786),
.B(n_1753),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1809),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1853),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1853),
.B(n_1823),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1865),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1786),
.B(n_1717),
.Y(n_1933)
);

AND2x4_ASAP7_75t_SL g1934 ( 
.A(n_1857),
.B(n_1685),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1775),
.B(n_1752),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1811),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1882),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1851),
.B(n_1797),
.Y(n_1938)
);

NOR2x1_ASAP7_75t_L g1939 ( 
.A(n_1892),
.B(n_1896),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1865),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1818),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1781),
.B(n_1752),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1822),
.Y(n_1943)
);

BUFx2_ASAP7_75t_SL g1944 ( 
.A(n_1796),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1820),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1824),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1827),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1771),
.A2(n_1724),
.B1(n_1728),
.B2(n_1726),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1790),
.B(n_1738),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1790),
.B(n_1738),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1839),
.B(n_1738),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1906),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1795),
.B(n_1739),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1828),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1806),
.B(n_1739),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1874),
.B(n_1826),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1800),
.B(n_1740),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1805),
.B(n_1740),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1830),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1768),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1771),
.A2(n_1724),
.B1(n_1728),
.B2(n_1726),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1769),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1906),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1770),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1829),
.A2(n_1728),
.B1(n_1726),
.B2(n_1702),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1803),
.B(n_1740),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1807),
.B(n_1742),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1803),
.B(n_1742),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1856),
.B(n_1721),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_L g1970 ( 
.A1(n_1785),
.A2(n_1702),
.B1(n_1735),
.B2(n_1716),
.Y(n_1970)
);

INVx6_ASAP7_75t_L g1971 ( 
.A(n_1774),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1881),
.Y(n_1972)
);

OR2x6_ASAP7_75t_L g1973 ( 
.A(n_1857),
.B(n_1880),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1773),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1849),
.B(n_1717),
.Y(n_1975)
);

NAND2x1p5_ASAP7_75t_L g1976 ( 
.A(n_1880),
.B(n_1698),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1812),
.B(n_1744),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1780),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1813),
.B(n_1746),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1856),
.B(n_1717),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1782),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1885),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1787),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1858),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1791),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1814),
.B(n_1746),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1793),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1778),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1834),
.B(n_1883),
.Y(n_1989)
);

INVx5_ASAP7_75t_L g1990 ( 
.A(n_1776),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1815),
.B(n_1747),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1870),
.B(n_1788),
.Y(n_1992)
);

INVx3_ASAP7_75t_L g1993 ( 
.A(n_1776),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1879),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_L g1995 ( 
.A(n_1817),
.B(n_1760),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1874),
.B(n_1743),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1816),
.B(n_1747),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1850),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1776),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1887),
.A2(n_1725),
.B1(n_1764),
.B2(n_1710),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1784),
.A2(n_1764),
.B1(n_1710),
.B2(n_1698),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1845),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1893),
.Y(n_2003)
);

BUFx3_ASAP7_75t_L g2004 ( 
.A(n_1858),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1896),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1835),
.A2(n_1702),
.B1(n_1735),
.B2(n_1654),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1835),
.A2(n_1733),
.B1(n_1674),
.B2(n_1734),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1794),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1870),
.B(n_1624),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1832),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1846),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1860),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1909),
.Y(n_2013)
);

BUFx12f_ASAP7_75t_L g2014 ( 
.A(n_1879),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1861),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_1848),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1863),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_SL g2018 ( 
.A1(n_1841),
.A2(n_1721),
.B1(n_1719),
.B2(n_1671),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1956),
.A2(n_1867),
.B1(n_1779),
.B2(n_1876),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1917),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1982),
.Y(n_2021)
);

AND2x4_ASAP7_75t_SL g2022 ( 
.A(n_1931),
.B(n_1857),
.Y(n_2022)
);

AOI222xp33_ASAP7_75t_L g2023 ( 
.A1(n_1956),
.A2(n_1798),
.B1(n_1876),
.B2(n_1836),
.C1(n_1810),
.C2(n_1872),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1931),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2010),
.B(n_1886),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1918),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2003),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1951),
.Y(n_2028)
);

NOR2xp67_ASAP7_75t_L g2029 ( 
.A(n_1990),
.B(n_1897),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1980),
.A2(n_1867),
.B1(n_1792),
.B2(n_1873),
.Y(n_2030)
);

NAND4xp25_ASAP7_75t_L g2031 ( 
.A(n_1948),
.B(n_1868),
.C(n_1852),
.D(n_1890),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1923),
.B(n_1772),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1924),
.B(n_1777),
.Y(n_2033)
);

NOR2x1p5_ASAP7_75t_L g2034 ( 
.A(n_2014),
.B(n_1847),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1951),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1927),
.Y(n_2036)
);

NOR2xp67_ASAP7_75t_L g2037 ( 
.A(n_1990),
.B(n_1842),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1953),
.B(n_1967),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1961),
.A2(n_1884),
.B1(n_1837),
.B2(n_1866),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1927),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_2013),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1922),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1922),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1919),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1957),
.Y(n_2045)
);

INVxp67_ASAP7_75t_L g2046 ( 
.A(n_1943),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1957),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1929),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1931),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_1937),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_1944),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1977),
.B(n_1825),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1958),
.Y(n_2053)
);

NOR2xp67_ASAP7_75t_L g2054 ( 
.A(n_1990),
.B(n_1854),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1916),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1958),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1949),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1975),
.A2(n_1933),
.B1(n_1921),
.B2(n_1992),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1949),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1936),
.Y(n_2060)
);

OAI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2018),
.A2(n_1868),
.B1(n_1903),
.B2(n_1901),
.C(n_1840),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1977),
.B(n_1825),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1979),
.B(n_1898),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1971),
.A2(n_1895),
.B1(n_1900),
.B2(n_1878),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_2005),
.Y(n_2065)
);

BUFx3_ASAP7_75t_L g2066 ( 
.A(n_2005),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1941),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1950),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1979),
.B(n_1905),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1950),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_1952),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1945),
.B(n_1911),
.Y(n_2072)
);

INVxp67_ASAP7_75t_SL g2073 ( 
.A(n_1963),
.Y(n_2073)
);

AOI222xp33_ASAP7_75t_L g2074 ( 
.A1(n_2014),
.A2(n_1988),
.B1(n_1926),
.B2(n_2000),
.C1(n_1810),
.C2(n_2017),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1994),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1990),
.B(n_1783),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1986),
.B(n_1749),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1986),
.B(n_1991),
.Y(n_2078)
);

NAND2x1p5_ASAP7_75t_L g2079 ( 
.A(n_1990),
.B(n_1845),
.Y(n_2079)
);

INVxp67_ASAP7_75t_L g2080 ( 
.A(n_1972),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1978),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1946),
.B(n_1864),
.Y(n_2082)
);

INVxp67_ASAP7_75t_SL g2083 ( 
.A(n_1916),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1955),
.B(n_1624),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_2051),
.B(n_1998),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2078),
.B(n_1968),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2020),
.Y(n_2087)
);

INVxp67_ASAP7_75t_L g2088 ( 
.A(n_2071),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2020),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2057),
.B(n_1955),
.Y(n_2090)
);

NAND3xp33_ASAP7_75t_L g2091 ( 
.A(n_2023),
.B(n_2006),
.C(n_2016),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2078),
.B(n_1968),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_2075),
.Y(n_2093)
);

INVxp67_ASAP7_75t_L g2094 ( 
.A(n_2073),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2026),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2057),
.B(n_2059),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2048),
.Y(n_2097)
);

NAND2x1_ASAP7_75t_L g2098 ( 
.A(n_2055),
.B(n_1971),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2038),
.B(n_1966),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2060),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2059),
.B(n_2009),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2067),
.Y(n_2102)
);

INVx4_ASAP7_75t_L g2103 ( 
.A(n_2079),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2021),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2041),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_2054),
.B(n_2065),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2044),
.B(n_2036),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2081),
.B(n_2050),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2038),
.B(n_1966),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2027),
.B(n_1989),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_2065),
.B(n_1919),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2052),
.B(n_2009),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2052),
.B(n_1997),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2058),
.B(n_1989),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2062),
.B(n_1997),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2072),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2032),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2068),
.B(n_1928),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2033),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2068),
.B(n_1992),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2062),
.B(n_1935),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_2066),
.Y(n_2122)
);

CKINVDCx16_ASAP7_75t_R g2123 ( 
.A(n_2075),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2045),
.B(n_1935),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2045),
.B(n_1942),
.Y(n_2125)
);

AND2x4_ASAP7_75t_SL g2126 ( 
.A(n_2024),
.B(n_1973),
.Y(n_2126)
);

AND2x4_ASAP7_75t_SL g2127 ( 
.A(n_2024),
.B(n_1973),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2025),
.B(n_1947),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2028),
.B(n_1954),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2047),
.B(n_1942),
.Y(n_2130)
);

INVx2_ASAP7_75t_SL g2131 ( 
.A(n_2066),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2101),
.B(n_2047),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2101),
.B(n_2053),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2087),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2086),
.B(n_2077),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2086),
.B(n_2077),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2096),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2092),
.B(n_2053),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2092),
.B(n_2056),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2096),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2099),
.B(n_2056),
.Y(n_2141)
);

NAND2x1_ASAP7_75t_L g2142 ( 
.A(n_2103),
.B(n_1971),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2099),
.B(n_2109),
.Y(n_2143)
);

NOR3xp33_ASAP7_75t_L g2144 ( 
.A(n_2091),
.B(n_2061),
.C(n_1969),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2094),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_2123),
.B(n_2093),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2095),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2097),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2109),
.B(n_2070),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2087),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2120),
.B(n_2070),
.Y(n_2151)
);

NOR2xp67_ASAP7_75t_R g2152 ( 
.A(n_2103),
.B(n_1971),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2089),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2113),
.B(n_2063),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2100),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2114),
.B(n_2036),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2102),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2113),
.B(n_2063),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2124),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_2122),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2120),
.B(n_2084),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2124),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2125),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2116),
.B(n_2040),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2107),
.B(n_2040),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2129),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2125),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2117),
.B(n_2028),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2115),
.B(n_2069),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2115),
.B(n_2069),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2144),
.A2(n_2074),
.B1(n_2019),
.B2(n_2112),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2137),
.B(n_2112),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2147),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2143),
.B(n_2121),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2142),
.A2(n_2037),
.B(n_2029),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2147),
.Y(n_2176)
);

INVx4_ASAP7_75t_L g2177 ( 
.A(n_2152),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2148),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2137),
.B(n_2104),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2161),
.B(n_2110),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2148),
.Y(n_2181)
);

AO21x1_ASAP7_75t_L g2182 ( 
.A1(n_2142),
.A2(n_2103),
.B(n_2106),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2134),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2134),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2155),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2140),
.B(n_2105),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2161),
.B(n_2121),
.Y(n_2187)
);

AOI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_2156),
.A2(n_2119),
.B1(n_2085),
.B2(n_2031),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2150),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2155),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2140),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2151),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2159),
.B(n_2088),
.Y(n_2193)
);

AOI32xp33_ASAP7_75t_L g2194 ( 
.A1(n_2160),
.A2(n_1939),
.A3(n_2131),
.B1(n_2022),
.B2(n_2127),
.Y(n_2194)
);

AOI21xp33_ASAP7_75t_L g2195 ( 
.A1(n_2145),
.A2(n_2108),
.B(n_2080),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_2146),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2159),
.A2(n_2106),
.B1(n_2098),
.B2(n_2049),
.Y(n_2197)
);

AOI32xp33_ASAP7_75t_L g2198 ( 
.A1(n_2143),
.A2(n_2131),
.A3(n_2127),
.B1(n_2126),
.B2(n_2064),
.Y(n_2198)
);

INVxp67_ASAP7_75t_SL g2199 ( 
.A(n_2150),
.Y(n_2199)
);

INVx2_ASAP7_75t_SL g2200 ( 
.A(n_2154),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2162),
.A2(n_2049),
.B1(n_2055),
.B2(n_1920),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2151),
.Y(n_2202)
);

INVx1_ASAP7_75t_SL g2203 ( 
.A(n_2165),
.Y(n_2203)
);

OAI21xp33_ASAP7_75t_L g2204 ( 
.A1(n_2165),
.A2(n_2107),
.B(n_2118),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2132),
.Y(n_2205)
);

OAI221xp5_ASAP7_75t_SL g2206 ( 
.A1(n_2198),
.A2(n_2039),
.B1(n_2030),
.B2(n_2133),
.C(n_2132),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_SL g2207 ( 
.A1(n_2177),
.A2(n_2197),
.B1(n_2196),
.B2(n_1994),
.Y(n_2207)
);

OAI31xp33_ASAP7_75t_L g2208 ( 
.A1(n_2197),
.A2(n_2034),
.A3(n_2111),
.B(n_2165),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2173),
.Y(n_2209)
);

AOI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_2182),
.A2(n_2111),
.B(n_2076),
.Y(n_2210)
);

OAI21xp33_ASAP7_75t_SL g2211 ( 
.A1(n_2194),
.A2(n_2158),
.B(n_2154),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2200),
.Y(n_2212)
);

OAI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2177),
.A2(n_1920),
.B1(n_1973),
.B2(n_1930),
.Y(n_2213)
);

NOR4xp25_ASAP7_75t_SL g2214 ( 
.A(n_2195),
.B(n_1996),
.C(n_1869),
.D(n_1912),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2176),
.Y(n_2215)
);

OAI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2171),
.A2(n_1973),
.B1(n_1930),
.B2(n_2046),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2203),
.A2(n_2188),
.B1(n_2204),
.B2(n_2196),
.Y(n_2217)
);

OAI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2175),
.A2(n_1996),
.B(n_2079),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2203),
.B(n_2135),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2178),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2201),
.A2(n_2166),
.B1(n_2164),
.B2(n_2168),
.C(n_2157),
.Y(n_2221)
);

AOI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2201),
.A2(n_2163),
.B1(n_2167),
.B2(n_2162),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2181),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2185),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2190),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_2179),
.B(n_2163),
.Y(n_2226)
);

OAI322xp33_ASAP7_75t_L g2227 ( 
.A1(n_2180),
.A2(n_2133),
.A3(n_2167),
.B1(n_2128),
.B2(n_2118),
.C1(n_2090),
.C2(n_2035),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2209),
.Y(n_2228)
);

OAI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2208),
.A2(n_2175),
.B1(n_2186),
.B2(n_2193),
.C(n_2191),
.Y(n_2229)
);

AOI33xp33_ASAP7_75t_L g2230 ( 
.A1(n_2216),
.A2(n_2205),
.A3(n_2202),
.B1(n_2192),
.B2(n_1833),
.B3(n_1903),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2217),
.A2(n_2172),
.B1(n_2107),
.B2(n_2199),
.Y(n_2231)
);

AOI211xp5_ASAP7_75t_L g2232 ( 
.A1(n_2206),
.A2(n_1912),
.B(n_1908),
.C(n_1666),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2207),
.A2(n_2187),
.B1(n_2174),
.B2(n_2169),
.Y(n_2233)
);

AOI222xp33_ASAP7_75t_L g2234 ( 
.A1(n_2211),
.A2(n_1831),
.B1(n_1819),
.B2(n_1799),
.C1(n_1850),
.C2(n_1938),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2221),
.B(n_2138),
.Y(n_2235)
);

AOI211xp5_ASAP7_75t_SL g2236 ( 
.A1(n_2216),
.A2(n_1995),
.B(n_2001),
.C(n_1999),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2222),
.A2(n_2138),
.B1(n_2139),
.B2(n_2141),
.Y(n_2237)
);

BUFx2_ASAP7_75t_SL g2238 ( 
.A(n_2210),
.Y(n_2238)
);

OAI32xp33_ASAP7_75t_L g2239 ( 
.A1(n_2218),
.A2(n_2079),
.A3(n_1932),
.B1(n_1940),
.B2(n_1796),
.Y(n_2239)
);

AOI221xp5_ASAP7_75t_L g2240 ( 
.A1(n_2227),
.A2(n_2139),
.B1(n_2149),
.B2(n_2141),
.C(n_2183),
.Y(n_2240)
);

AO22x2_ASAP7_75t_L g2241 ( 
.A1(n_2212),
.A2(n_1960),
.B1(n_1964),
.B2(n_1962),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2215),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2213),
.A2(n_2226),
.B1(n_2219),
.B2(n_2223),
.Y(n_2243)
);

OA22x2_ASAP7_75t_L g2244 ( 
.A1(n_2220),
.A2(n_2126),
.B1(n_2149),
.B2(n_2136),
.Y(n_2244)
);

NOR3xp33_ASAP7_75t_SL g2245 ( 
.A(n_2213),
.B(n_1908),
.C(n_1869),
.Y(n_2245)
);

INVx1_ASAP7_75t_SL g2246 ( 
.A(n_2224),
.Y(n_2246)
);

OAI222xp33_ASAP7_75t_L g2247 ( 
.A1(n_2226),
.A2(n_2135),
.B1(n_2136),
.B2(n_2090),
.C1(n_2169),
.C2(n_2170),
.Y(n_2247)
);

AOI221xp5_ASAP7_75t_L g2248 ( 
.A1(n_2225),
.A2(n_2184),
.B1(n_2189),
.B2(n_2170),
.C(n_2158),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2214),
.A2(n_2130),
.B1(n_2035),
.B2(n_2083),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2207),
.A2(n_1930),
.B1(n_1965),
.B2(n_1993),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2217),
.A2(n_2130),
.B1(n_1910),
.B2(n_2043),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2207),
.A2(n_1995),
.B(n_1915),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_SL g2253 ( 
.A(n_2252),
.B(n_1821),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2229),
.B(n_2233),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2246),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_SL g2256 ( 
.A(n_2245),
.B(n_1666),
.Y(n_2256)
);

OAI21xp33_ASAP7_75t_L g2257 ( 
.A1(n_2234),
.A2(n_1819),
.B(n_1799),
.Y(n_2257)
);

NAND4xp25_ASAP7_75t_L g2258 ( 
.A(n_2232),
.B(n_1831),
.C(n_1847),
.D(n_1932),
.Y(n_2258)
);

NOR3xp33_ASAP7_75t_L g2259 ( 
.A(n_2239),
.B(n_1888),
.C(n_1855),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2235),
.B(n_2153),
.Y(n_2260)
);

NAND4xp25_ASAP7_75t_L g2261 ( 
.A(n_2236),
.B(n_1940),
.C(n_1683),
.D(n_1662),
.Y(n_2261)
);

OAI321xp33_ASAP7_75t_L g2262 ( 
.A1(n_2243),
.A2(n_1976),
.A3(n_1970),
.B1(n_1925),
.B2(n_2082),
.C(n_2007),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_L g2263 ( 
.A(n_2238),
.B(n_2251),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2241),
.Y(n_2264)
);

NAND3xp33_ASAP7_75t_SL g2265 ( 
.A(n_2230),
.B(n_1875),
.C(n_1845),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_2231),
.B(n_2247),
.Y(n_2266)
);

NOR3xp33_ASAP7_75t_L g2267 ( 
.A(n_2250),
.B(n_1707),
.C(n_1719),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2237),
.B(n_1671),
.Y(n_2268)
);

OAI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2244),
.A2(n_1999),
.B1(n_2002),
.B2(n_1993),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2241),
.B(n_2153),
.Y(n_2270)
);

NAND2x1_ASAP7_75t_L g2271 ( 
.A(n_2228),
.B(n_1993),
.Y(n_2271)
);

NOR2x1_ASAP7_75t_L g2272 ( 
.A(n_2261),
.B(n_2242),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_L g2273 ( 
.A(n_2255),
.B(n_2263),
.C(n_2254),
.Y(n_2273)
);

OAI211xp5_ASAP7_75t_L g2274 ( 
.A1(n_2256),
.A2(n_1875),
.B(n_2240),
.C(n_2249),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2264),
.B(n_2248),
.Y(n_2275)
);

NOR2xp67_ASAP7_75t_L g2276 ( 
.A(n_2262),
.B(n_1999),
.Y(n_2276)
);

NAND3xp33_ASAP7_75t_L g2277 ( 
.A(n_2266),
.B(n_1774),
.C(n_1692),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2253),
.B(n_2268),
.Y(n_2278)
);

OAI211xp5_ASAP7_75t_L g2279 ( 
.A1(n_2257),
.A2(n_2259),
.B(n_2267),
.C(n_2258),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2270),
.Y(n_2280)
);

NAND3x1_ASAP7_75t_SL g2281 ( 
.A(n_2265),
.B(n_1774),
.C(n_1671),
.Y(n_2281)
);

NOR3x1_ASAP7_75t_L g2282 ( 
.A(n_2260),
.B(n_1705),
.C(n_1891),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2269),
.B(n_1974),
.Y(n_2283)
);

NOR3xp33_ASAP7_75t_L g2284 ( 
.A(n_2271),
.B(n_1808),
.C(n_1900),
.Y(n_2284)
);

AOI322xp5_ASAP7_75t_L g2285 ( 
.A1(n_2254),
.A2(n_1985),
.A3(n_2008),
.B1(n_1981),
.B2(n_1983),
.C1(n_1987),
.C2(n_1959),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2255),
.Y(n_2286)
);

NOR3xp33_ASAP7_75t_L g2287 ( 
.A(n_2261),
.B(n_1808),
.C(n_1900),
.Y(n_2287)
);

NOR2x1_ASAP7_75t_L g2288 ( 
.A(n_2261),
.B(n_1810),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2286),
.B(n_2011),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2280),
.B(n_2042),
.Y(n_2290)
);

NAND3xp33_ASAP7_75t_SL g2291 ( 
.A(n_2279),
.B(n_1705),
.C(n_1976),
.Y(n_2291)
);

NAND4xp75_ASAP7_75t_L g2292 ( 
.A(n_2272),
.B(n_1877),
.C(n_1862),
.D(n_1859),
.Y(n_2292)
);

NOR3xp33_ASAP7_75t_L g2293 ( 
.A(n_2273),
.B(n_1808),
.C(n_1878),
.Y(n_2293)
);

NOR3xp33_ASAP7_75t_L g2294 ( 
.A(n_2277),
.B(n_1889),
.C(n_1878),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2278),
.B(n_1859),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2283),
.Y(n_2296)
);

NOR2x1_ASAP7_75t_L g2297 ( 
.A(n_2288),
.B(n_1889),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2282),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2285),
.B(n_2012),
.Y(n_2299)
);

AOI211x1_ASAP7_75t_L g2300 ( 
.A1(n_2274),
.A2(n_2015),
.B(n_1877),
.C(n_1904),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_2275),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2281),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2289),
.Y(n_2303)
);

XOR2xp5_ASAP7_75t_L g2304 ( 
.A(n_2291),
.B(n_1895),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2292),
.A2(n_2276),
.B1(n_2287),
.B2(n_2284),
.Y(n_2305)
);

XOR2xp5_ASAP7_75t_L g2306 ( 
.A(n_2302),
.B(n_1877),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2301),
.B(n_2042),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2289),
.Y(n_2308)
);

NAND2x1p5_ASAP7_75t_L g2309 ( 
.A(n_2295),
.B(n_1889),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_2298),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2296),
.B(n_1859),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2290),
.B(n_2043),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2311),
.Y(n_2313)
);

OR2x6_ASAP7_75t_L g2314 ( 
.A(n_2303),
.B(n_2300),
.Y(n_2314)
);

AND4x1_ASAP7_75t_L g2315 ( 
.A(n_2306),
.B(n_2293),
.C(n_2297),
.D(n_2294),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2310),
.B(n_2299),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2308),
.Y(n_2317)
);

AOI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_2304),
.A2(n_1862),
.B1(n_1925),
.B2(n_1894),
.Y(n_2318)
);

OR3x2_ASAP7_75t_L g2319 ( 
.A(n_2305),
.B(n_1862),
.C(n_1902),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2307),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2312),
.B(n_1984),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2319),
.A2(n_2305),
.B1(n_2309),
.B2(n_2004),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2316),
.B(n_2044),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2313),
.Y(n_2324)
);

OAI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2317),
.A2(n_1715),
.B(n_1817),
.Y(n_2325)
);

XOR2x2_ASAP7_75t_L g2326 ( 
.A(n_2322),
.B(n_2315),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2324),
.A2(n_2314),
.B(n_2320),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2323),
.A2(n_2314),
.B1(n_2321),
.B2(n_2318),
.Y(n_2328)
);

NOR2x1p5_ASAP7_75t_L g2329 ( 
.A(n_2325),
.B(n_1984),
.Y(n_2329)
);

XOR2xp5_ASAP7_75t_L g2330 ( 
.A(n_2324),
.B(n_1891),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2329),
.Y(n_2331)
);

NOR2x1_ASAP7_75t_L g2332 ( 
.A(n_2327),
.B(n_2004),
.Y(n_2332)
);

OAI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2328),
.A2(n_1899),
.B1(n_1894),
.B2(n_2002),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2332),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2331),
.A2(n_2330),
.B1(n_2326),
.B2(n_1899),
.Y(n_2335)
);

AOI31xp33_ASAP7_75t_L g2336 ( 
.A1(n_2333),
.A2(n_1914),
.A3(n_1610),
.B(n_1913),
.Y(n_2336)
);

AOI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2335),
.A2(n_1934),
.B1(n_2002),
.B2(n_1789),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2337),
.B(n_2334),
.Y(n_2338)
);

BUFx24_ASAP7_75t_SL g2339 ( 
.A(n_2338),
.Y(n_2339)
);

AOI21xp33_ASAP7_75t_L g2340 ( 
.A1(n_2339),
.A2(n_2336),
.B(n_1688),
.Y(n_2340)
);


endmodule