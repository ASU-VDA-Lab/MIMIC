module real_jpeg_7185_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_173;
wire n_40;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_178;
wire n_67;
wire n_76;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_110;
wire n_61;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_0),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_0),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_0),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_0),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_0),
.B(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_3),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_3),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_4),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_4),
.B(n_193),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_14),
.Y(n_61)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_9),
.A2(n_29),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_9),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_9),
.B(n_50),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_9),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_12),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_12),
.B(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_13),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_13),
.Y(n_193)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_14),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_15),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_15),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_15),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_178),
.B1(n_283),
.B2(n_284),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_176),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_134),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_20),
.B(n_134),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.C(n_110),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_21),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_23),
.B(n_35),
.C(n_51),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_33),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_25),
.B(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_28),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_33),
.B(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_47),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_42),
.B2(n_46),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_37),
.B(n_42),
.C(n_47),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_39),
.Y(n_220)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_39),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_60),
.C(n_62),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_52),
.A2(n_53),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_54),
.A2(n_57),
.B1(n_146),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_54),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_55),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_56),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_57),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_57),
.Y(n_146)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_69),
.B(n_110),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_84),
.C(n_99),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_70),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_80),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_77),
.C(n_80),
.Y(n_133)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_83),
.Y(n_190)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_83),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_84),
.A2(n_99),
.B1(n_100),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_84),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_95),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_85),
.A2(n_86),
.B1(n_95),
.B2(n_96),
.Y(n_262)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_90),
.B(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_91),
.B(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_129),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_130),
.C(n_133),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_120),
.C(n_128),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_128),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_141),
.Y(n_140)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_158),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_149),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_175),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_178),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_278),
.B(n_282),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_264),
.B(n_277),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_250),
.B(n_263),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_226),
.B(n_249),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_216),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_216),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_197),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_198),
.C(n_206),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_185),
.B(n_192),
.C(n_194),
.Y(n_260)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_202),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_212),
.B(n_214),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.C(n_221),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_243),
.B(n_248),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_236),
.B(n_242),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_235),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_233),
.Y(n_244)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_260),
.C(n_261),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_253),
.Y(n_285)
);

FAx1_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.CI(n_258),
.CON(n_253),
.SN(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_256),
.C(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_276),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_276),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_270),
.C(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);


endmodule