module real_jpeg_31447_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_595, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_595;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_0),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_0),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_2),
.A2(n_178),
.B1(n_254),
.B2(n_258),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_2),
.A2(n_178),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_2),
.A2(n_178),
.B1(n_408),
.B2(n_411),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_3),
.A2(n_110),
.B1(n_115),
.B2(n_116),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_3),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_3),
.A2(n_115),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_3),
.A2(n_115),
.B1(n_375),
.B2(n_378),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_3),
.A2(n_115),
.B1(n_462),
.B2(n_465),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_4),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_4),
.A2(n_75),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_4),
.A2(n_75),
.B1(n_275),
.B2(n_281),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_5),
.A2(n_146),
.B1(n_342),
.B2(n_346),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_5),
.A2(n_146),
.B1(n_433),
.B2(n_436),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_5),
.A2(n_146),
.B1(n_533),
.B2(n_535),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_6),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_6),
.A2(n_100),
.B1(n_266),
.B2(n_270),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_7),
.B(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_7),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_7),
.B(n_119),
.Y(n_413)
);

OAI32xp33_ASAP7_75t_L g440 ( 
.A1(n_7),
.A2(n_441),
.A3(n_444),
.B1(n_446),
.B2(n_451),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_7),
.A2(n_371),
.B1(n_483),
.B2(n_486),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g514 ( 
.A1(n_7),
.A2(n_89),
.B(n_515),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_9),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_10),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_11),
.A2(n_60),
.B1(n_187),
.B2(n_190),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_11),
.A2(n_60),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B(n_592),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_13),
.B(n_593),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_14),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_16),
.A2(n_233),
.B1(n_234),
.B2(n_240),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_16),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_16),
.A2(n_233),
.B1(n_386),
.B2(n_392),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_16),
.A2(n_233),
.B1(n_489),
.B2(n_491),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_16),
.A2(n_233),
.B1(n_503),
.B2(n_507),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_17),
.Y(n_168)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_17),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_18),
.A2(n_81),
.B1(n_85),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_296),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_295),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_259),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_24),
.B(n_259),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_193),
.C(n_215),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_25),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_106),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_26),
.B(n_153),
.C(n_192),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_79),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_27),
.B(n_79),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_55),
.B1(n_67),
.B2(n_69),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_28),
.A2(n_67),
.B1(n_69),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_28),
.A2(n_55),
.B1(n_67),
.B2(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g431 ( 
.A1(n_28),
.A2(n_432),
.B(n_438),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_28),
.A2(n_67),
.B1(n_432),
.B2(n_488),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_43),
.Y(n_28)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

OAI22x1_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_31),
.Y(n_509)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_36),
.Y(n_550)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_38),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_40),
.Y(n_466)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_42),
.Y(n_464)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_42),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_43)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_44),
.Y(n_445)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_45),
.Y(n_379)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_47),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_47),
.Y(n_163)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_51),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_51),
.Y(n_437)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_58),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_59),
.Y(n_435)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_65),
.Y(n_209)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_65),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_66),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g556 ( 
.A(n_66),
.Y(n_556)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_67),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_68),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_68),
.B(n_371),
.Y(n_500)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_89),
.B1(n_96),
.B2(n_104),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_80),
.A2(n_89),
.B1(n_244),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_83),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_84),
.Y(n_247)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_84),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_88),
.A2(n_202),
.B(n_206),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_88),
.B(n_207),
.Y(n_206)
);

OAI22x1_ASAP7_75t_L g402 ( 
.A1(n_89),
.A2(n_329),
.B1(n_403),
.B2(n_407),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_89),
.A2(n_515),
.B(n_532),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_90),
.A2(n_97),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_90),
.A2(n_97),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_90),
.A2(n_105),
.B1(n_245),
.B2(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_90),
.B(n_461),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_90),
.A2(n_250),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_95),
.Y(n_512)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_102),
.Y(n_248)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_102),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_103),
.Y(n_332)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_103),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_103),
.Y(n_412)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_153),
.B1(n_191),
.B2(n_192),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_107),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_133),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_108),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

NAND2x1_ASAP7_75t_SL g293 ( 
.A(n_109),
.B(n_134),
.Y(n_293)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_111),
.Y(n_291)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_135)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_114),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_114),
.Y(n_319)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_119),
.A2(n_134),
.B1(n_145),
.B2(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_119),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_119),
.B(n_232),
.Y(n_338)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_130),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_123),
.Y(n_325)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_125),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_130),
.Y(n_322)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_132),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_132),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_145),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_134),
.B(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_136),
.Y(n_292)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_140),
.Y(n_312)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_152),
.Y(n_241)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_174),
.B1(n_183),
.B2(n_185),
.Y(n_153)
);

OAI22x1_ASAP7_75t_L g218 ( 
.A1(n_154),
.A2(n_174),
.B1(n_219),
.B2(n_229),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_154),
.A2(n_341),
.B(n_347),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_154),
.A2(n_347),
.B(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_155),
.A2(n_184),
.B1(n_186),
.B2(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_155),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_155),
.B(n_419),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_157),
.Y(n_271)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_160),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_165),
.B1(n_169),
.B2(n_173),
.Y(n_164)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_165),
.Y(n_346)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_168),
.Y(n_282)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_177),
.Y(n_190)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_177),
.Y(n_345)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_184),
.B(n_220),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_184),
.B(n_385),
.Y(n_416)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

BUFx4f_ASAP7_75t_L g310 ( 
.A(n_190),
.Y(n_310)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_194),
.B(n_216),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B1(n_210),
.B2(n_211),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_196),
.B(n_200),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_197),
.Y(n_459)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g490 ( 
.A(n_205),
.Y(n_490)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_211),
.A2(n_212),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_214),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_214),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_230),
.C(n_242),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_218),
.B(n_231),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_219),
.Y(n_419)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_224),
.Y(n_453)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_228),
.Y(n_391)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_229),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_229),
.B(n_371),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_242),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_252),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_243),
.B(n_252),
.Y(n_361)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_251),
.Y(n_523)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_253),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_294),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_284),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_273),
.B(n_283),
.Y(n_261)
);

NAND2x1_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_273),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_272),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_263),
.A2(n_374),
.B1(n_380),
.B2(n_381),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_263),
.B(n_565),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_263),
.A2(n_272),
.B1(n_374),
.B2(n_575),
.Y(n_574)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_272),
.B(n_374),
.Y(n_438)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_280),
.Y(n_393)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_338),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_348),
.B(n_590),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_299),
.B(n_301),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.C(n_306),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_336),
.C(n_339),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_SL g357 ( 
.A(n_307),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_326),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_308),
.A2(n_309),
.B1(n_326),
.B2(n_327),
.Y(n_420)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI32xp33_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.A3(n_313),
.B1(n_317),
.B2(n_320),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_334),
.Y(n_537)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_421),
.B(n_587),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_355),
.B(n_394),
.Y(n_350)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_351),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g587 ( 
.A(n_356),
.B(n_588),
.C(n_589),
.Y(n_587)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.C(n_362),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_363),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_373),
.C(n_382),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_364),
.B(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_371),
.B(n_372),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_371),
.B(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_371),
.B(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_371),
.B(n_553),
.Y(n_552)
);

OAI21xp33_ASAP7_75t_SL g565 ( 
.A1(n_371),
.A2(n_552),
.B(n_566),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_382),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_377),
.Y(n_495)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_395),
.B(n_397),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.C(n_420),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_401),
.A2(n_420),
.B1(n_469),
.B2(n_470),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_413),
.B1(n_414),
.B2(n_417),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_413),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_413),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_402),
.A2(n_413),
.B1(n_414),
.B2(n_417),
.Y(n_471)
);

INVx3_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_407),
.A2(n_459),
.B(n_460),
.Y(n_458)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_418),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_420),
.Y(n_469)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_472),
.B(n_585),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_467),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_425),
.B(n_586),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_430),
.C(n_439),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_430),
.A2(n_431),
.B1(n_439),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_435),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_438),
.B(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_458),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_458),
.Y(n_479)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_460),
.A2(n_502),
.B(n_510),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_461),
.B(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_467),
.Y(n_586)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_496),
.B(n_584),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_474),
.B(n_477),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.C(n_487),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_479),
.B(n_570),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_481),
.B(n_487),
.Y(n_570)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_488),
.Y(n_575)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

OAI321xp33_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_568),
.A3(n_577),
.B1(n_582),
.B2(n_583),
.C(n_595),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_528),
.B(n_567),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_499),
.A2(n_513),
.B(n_527),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_500),
.B(n_501),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g530 ( 
.A(n_502),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx2_ASAP7_75t_SL g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_521),
.Y(n_513)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_522),
.B(n_524),
.Y(n_521)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_538),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_529),
.B(n_538),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_563),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_539),
.B(n_563),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_551),
.B1(n_557),
.B2(n_562),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_541),
.B(n_545),
.Y(n_540)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_541),
.Y(n_562)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_560),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_559),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_569),
.B(n_571),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_571),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_573),
.C(n_576),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_572),
.B(n_580),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_573),
.A2(n_574),
.B1(n_576),
.B2(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_576),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_579),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_578),
.B(n_579),
.Y(n_582)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);


endmodule