module real_aes_6703_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_1034;
wire n_549;
wire n_571;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_1078;
wire n_384;
wire n_938;
wire n_744;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_951;
wire n_875;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_369;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_973;
wire n_1081;
wire n_1084;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_598;
wire n_404;
wire n_735;
wire n_1073;
wire n_713;
wire n_728;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_1014;
wire n_1083;
wire n_727;
wire n_649;
wire n_749;
wire n_385;
wire n_397;
wire n_663;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_1045;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g663 ( .A(n_0), .B(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g1080 ( .A1(n_1), .A2(n_230), .B1(n_523), .B2(n_1081), .Y(n_1080) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_2), .A2(n_170), .B1(n_317), .B2(n_449), .C1(n_451), .C2(n_455), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_3), .A2(n_245), .B1(n_488), .B2(n_610), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_4), .A2(n_100), .B1(n_752), .B2(n_753), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_5), .A2(n_152), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_6), .A2(n_78), .B1(n_455), .B2(n_919), .Y(n_918) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_7), .B(n_474), .Y(n_473) );
AO22x2_ASAP7_75t_L g398 ( .A1(n_8), .A2(n_216), .B1(n_390), .B2(n_395), .Y(n_398) );
INVx1_ASAP7_75t_L g1059 ( .A(n_8), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_9), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_10), .A2(n_161), .B1(n_419), .B2(n_422), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_11), .A2(n_342), .B1(n_440), .B2(n_468), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_12), .A2(n_148), .B1(n_490), .B2(n_555), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_13), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_14), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_15), .A2(n_186), .B1(n_471), .B2(n_645), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_16), .A2(n_241), .B1(n_555), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_17), .A2(n_103), .B1(n_752), .B2(n_760), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_18), .A2(n_305), .B1(n_759), .B2(n_760), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_19), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_20), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_21), .A2(n_291), .B1(n_614), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_22), .A2(n_221), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_23), .A2(n_292), .B1(n_425), .B2(n_776), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_24), .Y(n_536) );
AOI22xp5_ASAP7_75t_SL g630 ( .A1(n_25), .A2(n_238), .B1(n_490), .B2(n_631), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_26), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_27), .A2(n_289), .B1(n_614), .B2(n_753), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_28), .A2(n_244), .B1(n_419), .B2(n_610), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_29), .A2(n_349), .B1(n_483), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_30), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_31), .A2(n_235), .B1(n_422), .B2(n_486), .Y(n_945) );
AO22x2_ASAP7_75t_L g400 ( .A1(n_32), .A2(n_117), .B1(n_390), .B2(n_391), .Y(n_400) );
INVx1_ASAP7_75t_L g863 ( .A(n_33), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_34), .A2(n_165), .B1(n_413), .B2(n_426), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_35), .A2(n_56), .B1(n_486), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g948 ( .A1(n_36), .A2(n_59), .B1(n_407), .B2(n_419), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_37), .A2(n_64), .B1(n_482), .B2(n_622), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_38), .A2(n_278), .B1(n_455), .B2(n_668), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_39), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_40), .A2(n_60), .B1(n_384), .B2(n_421), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_41), .A2(n_155), .B1(n_422), .B2(n_619), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_42), .B(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_43), .A2(n_120), .B1(n_529), .B2(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_44), .B(n_471), .Y(n_792) );
INVx1_ASAP7_75t_L g1011 ( .A(n_45), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_46), .A2(n_351), .B1(n_444), .B2(n_666), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_47), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_48), .A2(n_306), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp5_ASAP7_75t_SL g629 ( .A1(n_49), .A2(n_299), .B1(n_488), .B2(n_556), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g766 ( .A1(n_50), .A2(n_284), .B1(n_304), .B2(n_504), .C1(n_598), .C2(n_714), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_51), .A2(n_283), .B1(n_436), .B2(n_1007), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_52), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_53), .Y(n_458) );
AOI22xp5_ASAP7_75t_SL g554 ( .A1(n_54), .A2(n_214), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_55), .A2(n_72), .B1(n_506), .B2(n_594), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_57), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g711 ( .A(n_58), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_61), .B(n_598), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_62), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g847 ( .A1(n_63), .A2(n_237), .B1(n_526), .B2(n_733), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g1012 ( .A1(n_65), .A2(n_91), .B1(n_455), .B2(n_476), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_66), .Y(n_534) );
INVx1_ASAP7_75t_L g868 ( .A(n_67), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_68), .A2(n_124), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_69), .A2(n_333), .B1(n_419), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_70), .A2(n_143), .B1(n_425), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_71), .A2(n_196), .B1(n_526), .B2(n_1037), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_73), .A2(n_90), .B1(n_655), .B2(n_658), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_74), .A2(n_210), .B1(n_472), .B2(n_645), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_75), .Y(n_812) );
AOI211xp5_ASAP7_75t_SL g367 ( .A1(n_76), .A2(n_368), .B(n_376), .C(n_1061), .Y(n_367) );
INVx1_ASAP7_75t_L g1070 ( .A(n_77), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_79), .A2(n_94), .B1(n_610), .B2(n_612), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_80), .A2(n_218), .B1(n_560), .B2(n_850), .Y(n_849) );
AOI22xp5_ASAP7_75t_SL g559 ( .A1(n_81), .A2(n_95), .B1(n_486), .B2(n_560), .Y(n_559) );
AO22x2_ASAP7_75t_L g394 ( .A1(n_82), .A2(n_249), .B1(n_390), .B2(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g1056 ( .A(n_82), .Y(n_1056) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_83), .A2(n_84), .B1(n_655), .B2(n_658), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_85), .A2(n_337), .B1(n_726), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_86), .A2(n_334), .B1(n_428), .B2(n_619), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_87), .A2(n_355), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_88), .A2(n_361), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_89), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_92), .A2(n_295), .B1(n_384), .B2(n_480), .Y(n_817) );
OA22x2_ASAP7_75t_L g747 ( .A1(n_93), .A2(n_748), .B1(n_749), .B2(n_767), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_93), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_96), .A2(n_197), .B1(n_523), .B2(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_97), .A2(n_110), .B1(n_479), .B2(n_486), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_98), .A2(n_106), .B1(n_440), .B2(n_504), .Y(n_941) );
INVx1_ASAP7_75t_L g551 ( .A(n_99), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_101), .A2(n_227), .B1(n_969), .B2(n_992), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_102), .A2(n_328), .B1(n_444), .B2(n_690), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_104), .A2(n_150), .B1(n_690), .B2(n_719), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_105), .A2(n_204), .B1(n_692), .B2(n_693), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_107), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_108), .B(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_109), .A2(n_135), .B1(n_759), .B2(n_882), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_111), .A2(n_267), .B1(n_556), .B2(n_850), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_112), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_113), .A2(n_266), .B1(n_523), .B2(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_114), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_115), .Y(n_706) );
INVx1_ASAP7_75t_L g964 ( .A(n_116), .Y(n_964) );
INVx1_ASAP7_75t_L g1060 ( .A(n_117), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_118), .A2(n_140), .B1(n_756), .B2(n_885), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_119), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_121), .A2(n_194), .B1(n_441), .B2(n_684), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_122), .A2(n_126), .B1(n_523), .B2(n_969), .Y(n_1019) );
INVx1_ASAP7_75t_L g1092 ( .A(n_123), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_123), .A2(n_1063), .B1(n_1084), .B2(n_1092), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_125), .Y(n_567) );
XNOR2x2_ASAP7_75t_L g648 ( .A(n_127), .B(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_128), .A2(n_714), .B(n_715), .C(n_721), .Y(n_713) );
INVx1_ASAP7_75t_L g972 ( .A(n_129), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_130), .A2(n_187), .B1(n_631), .B2(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1020 ( .A(n_131), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_132), .A2(n_185), .B1(n_526), .B2(n_1037), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_133), .A2(n_319), .B1(n_521), .B2(n_731), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_134), .A2(n_164), .B1(n_401), .B2(n_479), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_136), .A2(n_247), .B1(n_444), .B2(n_506), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_137), .A2(n_232), .B1(n_606), .B2(n_776), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_138), .A2(n_213), .B1(n_428), .B2(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_139), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g700 ( .A1(n_141), .A2(n_538), .B(n_701), .C(n_707), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_142), .A2(n_345), .B1(n_440), .B2(n_468), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_144), .A2(n_176), .B1(n_407), .B2(n_413), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_145), .A2(n_344), .B1(n_690), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_146), .A2(n_262), .B1(n_445), .B2(n_690), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_147), .Y(n_498) );
AND2x6_ASAP7_75t_L g370 ( .A(n_149), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_149), .Y(n_1053) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_151), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_153), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_154), .A2(n_248), .B1(n_683), .B2(n_870), .Y(n_982) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_156), .A2(n_339), .B1(n_407), .B2(n_614), .Y(n_1018) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_157), .A2(n_229), .B1(n_445), .B2(n_455), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_158), .A2(n_357), .B1(n_422), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_159), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g1041 ( .A1(n_160), .A2(n_179), .B1(n_200), .B2(n_451), .C1(n_506), .C2(n_670), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_162), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_163), .A2(n_256), .B1(n_529), .B2(n_756), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_166), .A2(n_363), .B1(n_871), .B2(n_919), .Y(n_965) );
INVx1_ASAP7_75t_L g978 ( .A(n_167), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_168), .Y(n_539) );
INVx1_ASAP7_75t_L g1074 ( .A(n_169), .Y(n_1074) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_171), .A2(n_177), .B1(n_425), .B2(n_969), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_172), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_173), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_174), .A2(n_254), .B1(n_533), .B2(n_759), .Y(n_902) );
AO22x2_ASAP7_75t_L g389 ( .A1(n_175), .A2(n_239), .B1(n_390), .B2(n_391), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_175), .B(n_1058), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_178), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_180), .A2(n_253), .B1(n_488), .B2(n_490), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_181), .A2(n_242), .B1(n_384), .B2(n_401), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_182), .A2(n_290), .B1(n_506), .B2(n_837), .Y(n_836) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_183), .A2(n_215), .B1(n_277), .B2(n_468), .C1(n_506), .C2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g970 ( .A1(n_184), .A2(n_330), .B1(n_401), .B2(n_555), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_188), .A2(n_366), .B1(n_468), .B2(n_506), .Y(n_1071) );
INVx1_ASAP7_75t_L g1066 ( .A(n_189), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_190), .Y(n_687) );
INVx1_ASAP7_75t_L g1073 ( .A(n_191), .Y(n_1073) );
AOI22xp5_ASAP7_75t_SL g633 ( .A1(n_192), .A2(n_264), .B1(n_562), .B2(n_634), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_193), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_195), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_198), .A2(n_325), .B1(n_413), .B2(n_521), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_199), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_201), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_202), .B(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_203), .A2(n_336), .B1(n_476), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_205), .A2(n_240), .B1(n_690), .B2(n_719), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_206), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g930 ( .A1(n_207), .A2(n_358), .B1(n_556), .B2(n_752), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_208), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_209), .A2(n_1063), .B1(n_1083), .B2(n_1084), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g1083 ( .A(n_209), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_211), .Y(n_805) );
INVx1_ASAP7_75t_L g867 ( .A(n_212), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_217), .A2(n_340), .B1(n_521), .B2(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_219), .B(n_471), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_220), .A2(n_353), .B1(n_425), .B2(n_428), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_222), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_223), .A2(n_281), .B1(n_521), .B2(n_524), .Y(n_520) );
XNOR2xp5_ASAP7_75t_L g889 ( .A(n_224), .B(n_890), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_225), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_226), .A2(n_258), .B1(n_634), .B2(n_845), .Y(n_844) );
AOI22xp5_ASAP7_75t_SL g858 ( .A1(n_228), .A2(n_859), .B1(n_886), .B2(n_887), .Y(n_858) );
INVx1_ASAP7_75t_L g887 ( .A(n_228), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_231), .A2(n_362), .B1(n_526), .B2(n_529), .Y(n_525) );
AND2x2_ASAP7_75t_L g374 ( .A(n_233), .B(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g467 ( .A1(n_234), .A2(n_313), .B1(n_456), .B2(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_236), .Y(n_681) );
INVx1_ASAP7_75t_L g862 ( .A(n_243), .Y(n_862) );
INVx1_ASAP7_75t_L g874 ( .A(n_246), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_250), .A2(n_297), .B1(n_482), .B2(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_251), .A2(n_346), .B1(n_658), .B2(n_996), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_252), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_255), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_257), .A2(n_332), .B1(n_845), .B2(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_259), .A2(n_293), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_260), .A2(n_303), .B1(n_692), .B2(n_764), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_261), .A2(n_279), .B1(n_480), .B2(n_524), .Y(n_1031) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_263), .B(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_265), .A2(n_302), .B1(n_775), .B2(n_776), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_268), .A2(n_365), .B1(n_610), .B2(n_658), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_269), .Y(n_568) );
INVx1_ASAP7_75t_L g390 ( .A(n_270), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_270), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_271), .A2(n_276), .B1(n_692), .B2(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1067 ( .A(n_272), .Y(n_1067) );
INVx1_ASAP7_75t_L g915 ( .A(n_273), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_274), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_275), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_280), .A2(n_322), .B1(n_479), .B2(n_731), .Y(n_971) );
INVx1_ASAP7_75t_L g913 ( .A(n_282), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_285), .Y(n_576) );
INVx1_ASAP7_75t_L g979 ( .A(n_286), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_287), .A2(n_331), .B1(n_441), .B2(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_288), .B(n_870), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_294), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_296), .A2(n_323), .B1(n_440), .B2(n_444), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g897 ( .A(n_298), .B(n_645), .Y(n_897) );
AO22x2_ASAP7_75t_L g797 ( .A1(n_300), .A2(n_798), .B1(n_819), .B2(n_820), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_300), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_301), .A2(n_326), .B1(n_505), .B2(n_594), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_307), .Y(n_830) );
INVx1_ASAP7_75t_L g375 ( .A(n_308), .Y(n_375) );
AOI22xp5_ASAP7_75t_SL g974 ( .A1(n_309), .A2(n_975), .B1(n_998), .B2(n_999), .Y(n_974) );
INVx1_ASAP7_75t_L g999 ( .A(n_309), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_310), .A2(n_318), .B1(n_611), .B2(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_311), .Y(n_781) );
INVx1_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
XOR2x2_ASAP7_75t_L g1023 ( .A(n_314), .B(n_1024), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_315), .B(n_436), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_316), .B(n_693), .Y(n_896) );
AOI22xp5_ASAP7_75t_SL g492 ( .A1(n_320), .A2(n_493), .B1(n_543), .B2(n_544), .Y(n_492) );
INVx1_ASAP7_75t_L g544 ( .A(n_320), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_321), .B(n_664), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_324), .A2(n_341), .B1(n_666), .B2(n_668), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_327), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_329), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_335), .Y(n_923) );
INVx1_ASAP7_75t_L g741 ( .A(n_338), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_343), .B(n_436), .Y(n_960) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_347), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_348), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_350), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_352), .A2(n_770), .B1(n_771), .B2(n_796), .Y(n_769) );
INVx1_ASAP7_75t_L g796 ( .A(n_352), .Y(n_796) );
INVx1_ASAP7_75t_L g873 ( .A(n_354), .Y(n_873) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_356), .B(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_359), .Y(n_917) );
OA22x2_ASAP7_75t_L g579 ( .A1(n_360), .A2(n_580), .B1(n_581), .B2(n_623), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_360), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g938 ( .A(n_364), .Y(n_938) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_371), .Y(n_1052) );
OAI21xp5_ASAP7_75t_L g1090 ( .A1(n_372), .A2(n_1051), .B(n_1091), .Y(n_1090) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_825), .B1(n_1046), .B2(n_1047), .C(n_1048), .Y(n_376) );
INVx1_ASAP7_75t_L g1046 ( .A(n_377), .Y(n_1046) );
AOI22xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_675), .B1(n_823), .B2(n_824), .Y(n_377) );
INVx1_ASAP7_75t_L g823 ( .A(n_378), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_548), .B1(n_673), .B2(n_674), .Y(n_378) );
INVx1_ASAP7_75t_L g673 ( .A(n_379), .Y(n_673) );
AO22x1_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_459), .B1(n_460), .B2(n_547), .Y(n_379) );
INVx2_ASAP7_75t_SL g547 ( .A(n_380), .Y(n_547) );
XOR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_458), .Y(n_380) );
NAND4xp75_ASAP7_75t_L g381 ( .A(n_382), .B(n_417), .C(n_431), .D(n_448), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_406), .Y(n_382) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g479 ( .A(n_385), .Y(n_479) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_SL g538 ( .A(n_386), .Y(n_538) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_386), .Y(n_611) );
BUFx2_ASAP7_75t_SL g631 ( .A(n_386), .Y(n_631) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_396), .Y(n_386) );
AND2x6_ASAP7_75t_L g403 ( .A(n_387), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g421 ( .A(n_387), .B(n_412), .Y(n_421) );
AND2x6_ASAP7_75t_L g450 ( .A(n_387), .B(n_447), .Y(n_450) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_393), .Y(n_387) );
AND2x2_ASAP7_75t_L g427 ( .A(n_388), .B(n_394), .Y(n_427) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g410 ( .A(n_389), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_389), .B(n_394), .Y(n_416) );
AND2x2_ASAP7_75t_L g443 ( .A(n_389), .B(n_398), .Y(n_443) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_392), .Y(n_395) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g411 ( .A(n_394), .Y(n_411) );
INVx1_ASAP7_75t_L g454 ( .A(n_394), .Y(n_454) );
AND2x2_ASAP7_75t_L g423 ( .A(n_396), .B(n_410), .Y(n_423) );
AND2x4_ASAP7_75t_L g426 ( .A(n_396), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g429 ( .A(n_396), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_396), .B(n_410), .Y(n_542) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
OR2x2_ASAP7_75t_L g405 ( .A(n_397), .B(n_400), .Y(n_405) );
AND2x2_ASAP7_75t_L g412 ( .A(n_397), .B(n_400), .Y(n_412) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_400), .Y(n_447) );
AND2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g511 ( .A(n_399), .Y(n_511) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g415 ( .A(n_400), .Y(n_415) );
INVx1_ASAP7_75t_L g782 ( .A(n_401), .Y(n_782) );
INVx5_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx4_ASAP7_75t_L g533 ( .A(n_402), .Y(n_533) );
INVx2_ASAP7_75t_SL g619 ( .A(n_402), .Y(n_619) );
INVx1_ASAP7_75t_L g652 ( .A(n_402), .Y(n_652) );
INVx2_ASAP7_75t_L g879 ( .A(n_402), .Y(n_879) );
INVx11_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx11_ASAP7_75t_L g489 ( .A(n_403), .Y(n_489) );
AND2x4_ASAP7_75t_L g438 ( .A(n_404), .B(n_427), .Y(n_438) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g496 ( .A(n_405), .B(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g621 ( .A(n_407), .Y(n_621) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_407), .Y(n_884) );
INVx5_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g482 ( .A(n_408), .Y(n_482) );
INVx4_ASAP7_75t_L g528 ( .A(n_408), .Y(n_528) );
INVx3_ASAP7_75t_L g556 ( .A(n_408), .Y(n_556) );
INVx2_ASAP7_75t_L g816 ( .A(n_408), .Y(n_816) );
BUFx3_ASAP7_75t_L g993 ( .A(n_408), .Y(n_993) );
INVx8_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_410), .B(n_412), .Y(n_703) );
INVx1_ASAP7_75t_L g446 ( .A(n_411), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_412), .B(n_427), .Y(n_434) );
AND2x6_ASAP7_75t_L g472 ( .A(n_412), .B(n_427), .Y(n_472) );
BUFx2_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
BUFx2_ASAP7_75t_L g529 ( .A(n_413), .Y(n_529) );
BUFx4f_ASAP7_75t_SL g885 ( .A(n_413), .Y(n_885) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_413), .Y(n_1037) );
INVx6_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g622 ( .A(n_414), .Y(n_622) );
INVx1_ASAP7_75t_SL g733 ( .A(n_414), .Y(n_733) );
INVx1_ASAP7_75t_SL g969 ( .A(n_414), .Y(n_969) );
OR2x6_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g442 ( .A(n_415), .Y(n_442) );
INVx1_ASAP7_75t_L g430 ( .A(n_416), .Y(n_430) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_424), .Y(n_417) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_420), .A2(n_531), .B1(n_532), .B2(n_534), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_420), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g752 ( .A(n_420), .Y(n_752) );
INVx2_ASAP7_75t_L g850 ( .A(n_420), .Y(n_850) );
INVx6_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g490 ( .A(n_421), .Y(n_490) );
BUFx3_ASAP7_75t_L g614 ( .A(n_421), .Y(n_614) );
BUFx3_ASAP7_75t_L g653 ( .A(n_421), .Y(n_653) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g555 ( .A(n_423), .Y(n_555) );
BUFx3_ASAP7_75t_L g608 ( .A(n_423), .Y(n_608) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_423), .Y(n_1030) );
BUFx2_ASAP7_75t_L g882 ( .A(n_425), .Y(n_882) );
BUFx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_426), .Y(n_523) );
BUFx3_ASAP7_75t_L g636 ( .A(n_426), .Y(n_636) );
INVx2_ASAP7_75t_L g846 ( .A(n_426), .Y(n_846) );
INVx1_ASAP7_75t_L g497 ( .A(n_427), .Y(n_497) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g486 ( .A(n_429), .Y(n_486) );
BUFx3_ASAP7_75t_L g524 ( .A(n_429), .Y(n_524) );
BUFx3_ASAP7_75t_L g634 ( .A(n_429), .Y(n_634) );
BUFx2_ASAP7_75t_SL g655 ( .A(n_429), .Y(n_655) );
BUFx2_ASAP7_75t_L g731 ( .A(n_429), .Y(n_731) );
BUFx2_ASAP7_75t_SL g990 ( .A(n_429), .Y(n_990) );
AND2x2_ASAP7_75t_L g562 ( .A(n_430), .B(n_511), .Y(n_562) );
OA211x2_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_435), .C(n_439), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_433), .A2(n_496), .B1(n_498), .B2(n_499), .Y(n_495) );
INVx2_ASAP7_75t_L g589 ( .A(n_433), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_433), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_433), .A2(n_585), .B1(n_978), .B2(n_979), .Y(n_977) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_433), .Y(n_1068) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g566 ( .A(n_434), .Y(n_566) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
INVx5_ASAP7_75t_L g645 ( .A(n_437), .Y(n_645) );
INVx2_ASAP7_75t_L g664 ( .A(n_437), .Y(n_664) );
INVx4_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g667 ( .A(n_441), .Y(n_667) );
BUFx2_ASAP7_75t_L g690 ( .A(n_441), .Y(n_690) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AND2x4_ASAP7_75t_L g452 ( .A(n_443), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g456 ( .A(n_443), .B(n_457), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_443), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_SL g720 ( .A(n_444), .Y(n_720) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g476 ( .A(n_445), .Y(n_476) );
BUFx2_ASAP7_75t_SL g668 ( .A(n_445), .Y(n_668) );
BUFx2_ASAP7_75t_SL g919 ( .A(n_445), .Y(n_919) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g516 ( .A(n_446), .Y(n_516) );
INVx1_ASAP7_75t_L g515 ( .A(n_447), .Y(n_515) );
INVx2_ASAP7_75t_L g834 ( .A(n_449), .Y(n_834) );
INVx2_ASAP7_75t_SL g866 ( .A(n_449), .Y(n_866) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g465 ( .A(n_450), .Y(n_465) );
INVx4_ASAP7_75t_L g501 ( .A(n_450), .Y(n_501) );
INVx2_ASAP7_75t_L g640 ( .A(n_450), .Y(n_640) );
BUFx3_ASAP7_75t_L g714 ( .A(n_450), .Y(n_714) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_452), .Y(n_468) );
BUFx4f_ASAP7_75t_SL g504 ( .A(n_452), .Y(n_504) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_452), .Y(n_684) );
BUFx2_ASAP7_75t_L g808 ( .A(n_452), .Y(n_808) );
INVx1_ASAP7_75t_L g457 ( .A(n_454), .Y(n_457) );
BUFx4f_ASAP7_75t_SL g598 ( .A(n_455), .Y(n_598) );
INVx2_ASAP7_75t_L g727 ( .A(n_455), .Y(n_727) );
BUFx12f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_456), .Y(n_506) );
BUFx6f_ASAP7_75t_L g871 ( .A(n_456), .Y(n_871) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AO22x2_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_492), .B1(n_545), .B2(n_546), .Y(n_460) );
INVx4_ASAP7_75t_SL g545 ( .A(n_461), .Y(n_545) );
XOR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_491), .Y(n_461) );
NAND3x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .C(n_484), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_469), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_466), .B(n_467), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_465), .A2(n_938), .B(n_939), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g963 ( .A1(n_465), .A2(n_964), .B(n_965), .Y(n_963) );
OAI21xp5_ASAP7_75t_SL g1010 ( .A1(n_465), .A2(n_1011), .B(n_1012), .Y(n_1010) );
INVx2_ASAP7_75t_L g575 ( .A(n_468), .Y(n_575) );
INVx4_ASAP7_75t_L g595 ( .A(n_468), .Y(n_595) );
BUFx2_ASAP7_75t_L g837 ( .A(n_468), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .C(n_475), .Y(n_469) );
INVx1_ASAP7_75t_L g694 ( .A(n_471), .Y(n_694) );
BUFx4f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g764 ( .A(n_472), .Y(n_764) );
INVx1_ASAP7_75t_SL g842 ( .A(n_472), .Y(n_842) );
BUFx2_ASAP7_75t_L g1007 ( .A(n_472), .Y(n_1007) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_481), .Y(n_477) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g736 ( .A(n_488), .Y(n_736) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
INVx2_ASAP7_75t_SL g760 ( .A(n_489), .Y(n_760) );
INVx4_ASAP7_75t_L g1027 ( .A(n_489), .Y(n_1027) );
INVx1_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
INVx1_ASAP7_75t_L g543 ( .A(n_493), .Y(n_543) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_518), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .C(n_507), .Y(n_494) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx2_ASAP7_75t_L g586 ( .A(n_496), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g500 ( .A1(n_501), .A2(n_502), .B(n_503), .Y(n_500) );
OAI22xp5_ASAP7_75t_SL g573 ( .A1(n_501), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_573) );
BUFx2_ASAP7_75t_L g591 ( .A(n_501), .Y(n_591) );
INVx4_ASAP7_75t_L g670 ( .A(n_501), .Y(n_670) );
OAI21xp5_ASAP7_75t_SL g788 ( .A1(n_501), .A2(n_789), .B(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g922 ( .A(n_504), .Y(n_922) );
BUFx4f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g686 ( .A(n_506), .Y(n_686) );
OAI22xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_512), .B1(n_513), .B2(n_517), .Y(n_507) );
OAI22xp5_ASAP7_75t_SL g564 ( .A1(n_508), .A2(n_565), .B1(n_567), .B2(n_568), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_508), .A2(n_513), .B1(n_873), .B2(n_874), .Y(n_872) );
INVx3_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g811 ( .A(n_509), .Y(n_811) );
INVx4_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx3_ASAP7_75t_L g601 ( .A(n_510), .Y(n_601) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_510), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_510), .A2(n_513), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_513), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_599) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_514), .A2(n_810), .B1(n_811), .B2(n_812), .Y(n_809) );
CKINVDCx16_ASAP7_75t_R g987 ( .A(n_514), .Y(n_987) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .C(n_535), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g775 ( .A(n_522), .Y(n_775) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g777 ( .A(n_524), .Y(n_777) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g756 ( .A(n_528), .Y(n_756) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_528), .Y(n_779) );
INVx1_ASAP7_75t_L g705 ( .A(n_529), .Y(n_705) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B1(n_539), .B2(n_540), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_537), .A2(n_540), .B1(n_785), .B2(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_540), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g674 ( .A(n_548), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_577), .B1(n_671), .B2(n_672), .Y(n_548) );
INVx1_ASAP7_75t_SL g671 ( .A(n_549), .Y(n_671) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
XNOR2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND3x1_ASAP7_75t_SL g552 ( .A(n_553), .B(n_558), .C(n_563), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
BUFx2_ASAP7_75t_L g697 ( .A(n_555), .Y(n_697) );
INVx1_ASAP7_75t_L g754 ( .A(n_555), .Y(n_754) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g709 ( .A(n_560), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .C(n_573), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_565), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g662 ( .A(n_566), .Y(n_662) );
INVx1_ASAP7_75t_SL g864 ( .A(n_566), .Y(n_864) );
OAI21xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_571), .B(n_572), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_570), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
INVx1_ASAP7_75t_L g672 ( .A(n_577), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_624), .B2(n_625), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_603), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .C(n_599), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_587), .B2(n_588), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_585), .A2(n_1066), .B1(n_1067), .B2(n_1068), .Y(n_1065) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g802 ( .A(n_586), .Y(n_802) );
INVx1_ASAP7_75t_SL g914 ( .A(n_586), .Y(n_914) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_588), .A2(n_716), .B(n_717), .C(n_718), .Y(n_715) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_593), .B2(n_596), .C(n_597), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g865 ( .A1(n_593), .A2(n_866), .B1(n_867), .B2(n_868), .C(n_869), .Y(n_865) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_601), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
NOR2xp67_ASAP7_75t_L g603 ( .A(n_604), .B(n_615), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx4f_ASAP7_75t_SL g658 ( .A(n_608), .Y(n_658) );
INVx1_ASAP7_75t_SL g740 ( .A(n_610), .Y(n_740) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx3_ASAP7_75t_L g759 ( .A(n_611), .Y(n_759) );
INVx3_ASAP7_75t_L g997 ( .A(n_611), .Y(n_997) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_613), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_647), .B2(n_648), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
XOR2x2_ASAP7_75t_L g828 ( .A(n_627), .B(n_829), .Y(n_828) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_646), .Y(n_627) );
NAND4xp75_ASAP7_75t_SL g628 ( .A(n_629), .B(n_630), .C(n_632), .D(n_637), .Y(n_628) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_636), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_641), .Y(n_638) );
OAI222xp33_ASAP7_75t_L g680 ( .A1(n_640), .A2(n_681), .B1(n_682), .B2(n_685), .C1(n_686), .C2(n_687), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_645), .Y(n_692) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_645), .Y(n_794) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_650), .B(n_656), .C(n_660), .D(n_669), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx3_ASAP7_75t_L g1035 ( .A(n_653), .Y(n_1035) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
OA211x2_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_663), .C(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g824 ( .A(n_675), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_744), .B1(n_745), .B2(n_822), .Y(n_675) );
INVx1_ASAP7_75t_L g822 ( .A(n_676), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_710), .B1(n_742), .B2(n_743), .Y(n_676) );
INVx1_ASAP7_75t_L g743 ( .A(n_677), .Y(n_743) );
NAND3x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_695), .C(n_700), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_688), .Y(n_679) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g723 ( .A(n_684), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
OAI22xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_701) );
BUFx2_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx2_ASAP7_75t_L g742 ( .A(n_710), .Y(n_742) );
XNOR2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_728), .Y(n_712) );
INVx3_ASAP7_75t_L g806 ( .A(n_714), .Y(n_806) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_734), .C(n_738), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AO22x1_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_768), .B2(n_821), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g767 ( .A(n_749), .Y(n_767) );
NAND4xp75_ASAP7_75t_L g749 ( .A(n_750), .B(n_757), .C(n_762), .D(n_766), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_755), .Y(n_750) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .Y(n_757) );
AND2x2_ASAP7_75t_SL g762 ( .A(n_763), .B(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g821 ( .A(n_768), .Y(n_821) );
XNOR2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_797), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_SL g771 ( .A(n_772), .B(n_787), .Y(n_771) );
NOR3xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_780), .C(n_784), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g1081 ( .A(n_782), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .C(n_795), .Y(n_791) );
INVx1_ASAP7_75t_SL g819 ( .A(n_798), .Y(n_819) );
AND2x2_ASAP7_75t_SL g798 ( .A(n_799), .B(n_813), .Y(n_798) );
NOR3xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_804), .C(n_809), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B(n_807), .Y(n_804) );
OAI21xp33_ASAP7_75t_L g980 ( .A1(n_806), .A2(n_981), .B(n_982), .Y(n_980) );
AND4x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .C(n_817), .D(n_818), .Y(n_813) );
INVx1_ASAP7_75t_L g1047 ( .A(n_825), .Y(n_1047) );
XNOR2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_952), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_828), .B1(n_852), .B2(n_853), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_843), .C(n_848), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_838), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g833 ( .A1(n_834), .A2(n_835), .B(n_836), .Y(n_833) );
OAI21xp5_ASAP7_75t_SL g892 ( .A1(n_834), .A2(n_893), .B(n_894), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx1_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_847), .Y(n_843) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AND2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
OAI22xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_904), .B1(n_905), .B2(n_951), .Y(n_853) );
INVx1_ASAP7_75t_L g951 ( .A(n_854), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B1(n_888), .B2(n_889), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_SL g886 ( .A(n_859), .Y(n_886) );
AND2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_875), .Y(n_859) );
NOR3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_865), .C(n_872), .Y(n_860) );
OAI21xp33_ASAP7_75t_L g916 ( .A1(n_866), .A2(n_917), .B(n_918), .Y(n_916) );
OAI21xp33_ASAP7_75t_SL g1069 ( .A1(n_866), .A2(n_1070), .B(n_1071), .Y(n_1069) );
BUFx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_880), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_883), .Y(n_880) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NAND4xp75_ASAP7_75t_SL g890 ( .A(n_891), .B(n_899), .C(n_902), .D(n_903), .Y(n_890) );
NOR2xp67_ASAP7_75t_L g891 ( .A(n_892), .B(n_895), .Y(n_891) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .C(n_898), .Y(n_895) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .B1(n_933), .B2(n_934), .Y(n_907) );
INVx1_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_932), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_925), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_916), .C(n_920), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_922), .B1(n_923), .B2(n_924), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_929), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
AO22x1_ASAP7_75t_SL g1022 ( .A1(n_933), .A2(n_934), .B1(n_1023), .B2(n_1042), .Y(n_1022) );
INVx3_ASAP7_75t_SL g933 ( .A(n_934), .Y(n_933) );
XOR2x2_ASAP7_75t_L g934 ( .A(n_935), .B(n_950), .Y(n_934) );
NAND2xp5_ASAP7_75t_SL g935 ( .A(n_936), .B(n_943), .Y(n_935) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_937), .B(n_940), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_947), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_1000), .B1(n_1044), .B2(n_1045), .Y(n_952) );
INVx1_ASAP7_75t_L g1044 ( .A(n_953), .Y(n_1044) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
OAI22xp5_ASAP7_75t_SL g954 ( .A1(n_955), .A2(n_956), .B1(n_973), .B2(n_974), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
XOR2x2_ASAP7_75t_L g956 ( .A(n_957), .B(n_972), .Y(n_956) );
NAND4xp75_ASAP7_75t_SL g957 ( .A(n_958), .B(n_966), .C(n_970), .D(n_971), .Y(n_957) );
NOR2xp67_ASAP7_75t_SL g958 ( .A(n_959), .B(n_963), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .C(n_962), .Y(n_959) );
AND2x2_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx2_ASAP7_75t_SL g998 ( .A(n_975), .Y(n_998) );
AND2x2_ASAP7_75t_SL g975 ( .A(n_976), .B(n_988), .Y(n_975) );
NOR3xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_980), .C(n_983), .Y(n_976) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
AND4x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_991), .C(n_994), .D(n_995), .Y(n_988) );
INVx3_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1000), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1021), .B1(n_1022), .B2(n_1043), .Y(n_1000) );
INVx1_ASAP7_75t_SL g1043 ( .A(n_1001), .Y(n_1043) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
XOR2x2_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1020), .Y(n_1002) );
NAND2x1p5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1013), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1010), .Y(n_1004) );
NAND3xp33_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1008), .C(n_1009), .Y(n_1005) );
NOR2x1_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1023), .Y(n_1042) );
NAND4xp75_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1032), .C(n_1038), .D(n_1041), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1031), .Y(n_1025) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1036), .Y(n_1032) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
AND2x2_ASAP7_75t_SL g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_SL g1048 ( .A(n_1049), .Y(n_1048) );
NOR2x1_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1054), .Y(n_1049) );
OR2x2_ASAP7_75t_SL g1098 ( .A(n_1050), .B(n_1055), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1053), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
OAI322xp33_ASAP7_75t_L g1061 ( .A1(n_1052), .A2(n_1062), .A3(n_1085), .B1(n_1089), .B2(n_1092), .C1(n_1093), .C2(n_1096), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1052), .B(n_1088), .Y(n_1091) );
CKINVDCx16_ASAP7_75t_R g1088 ( .A(n_1053), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_1055), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_1063), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1075), .Y(n_1063) );
NOR3xp33_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1069), .C(n_1072), .Y(n_1064) );
NOR2xp33_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1079), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1082), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
CKINVDCx16_ASAP7_75t_R g1089 ( .A(n_1090), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_1097), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_1098), .Y(n_1097) );
endmodule