module fake_jpeg_12081_n_120 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_29),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_1),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_9),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_18),
.B1(n_15),
.B2(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_15),
.B1(n_23),
.B2(n_17),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_23),
.B1(n_11),
.B2(n_13),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_13),
.B1(n_21),
.B2(n_16),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_16),
.B1(n_21),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_23),
.B1(n_4),
.B2(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_65),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_62),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_28),
.A2(n_3),
.B(n_4),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_32),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_3),
.A3(n_6),
.B1(n_10),
.B2(n_35),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_47),
.B(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_74),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_54),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_47),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_63),
.B1(n_51),
.B2(n_53),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_79),
.B1(n_77),
.B2(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_78),
.B1(n_73),
.B2(n_81),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_71),
.B1(n_80),
.B2(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_70),
.Y(n_96)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_74),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_82),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_80),
.B1(n_63),
.B2(n_51),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_88),
.C(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_104),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_99),
.B(n_86),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_98),
.B(n_94),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_85),
.C(n_89),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_R g108 ( 
.A1(n_106),
.A2(n_107),
.B1(n_93),
.B2(n_103),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.Y(n_112)
);

AO221x1_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_87),
.B1(n_101),
.B2(n_90),
.C(n_91),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_91),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_83),
.C(n_87),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_115),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_111),
.B1(n_92),
.B2(n_55),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_55),
.B(n_82),
.Y(n_120)
);


endmodule