module fake_jpeg_31682_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_5),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_1),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_60),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_51),
.B1(n_52),
.B2(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_49),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_49),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_54),
.B1(n_61),
.B2(n_48),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_4),
.C(n_6),
.Y(n_107)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_96),
.C(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_64),
.B(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_52),
.B1(n_65),
.B2(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_106),
.B1(n_107),
.B2(n_17),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_89),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_8),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_96),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_11),
.C(n_12),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_129),
.B(n_46),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_127),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_47),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_141)
);

NOR4xp25_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_123),
.C(n_114),
.D(n_125),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_117),
.C(n_39),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_36),
.B(n_37),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_23),
.C(n_25),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_141),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_35),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_149),
.B1(n_38),
.B2(n_45),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_147),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_119),
.B(n_41),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_144),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_135),
.C(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_143),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_152),
.CI(n_134),
.CON(n_159),
.SN(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_155),
.B(n_148),
.C(n_151),
.D(n_134),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_160),
.Y(n_161)
);


endmodule