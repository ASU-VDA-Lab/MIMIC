module fake_jpeg_30825_n_449 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_449);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_449;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_56),
.B(n_72),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_60),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_65),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_33),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_1),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_82),
.Y(n_145)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_30),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_84),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_2),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_31),
.B1(n_20),
.B2(n_41),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_93),
.A2(n_110),
.B1(n_124),
.B2(n_126),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_41),
.B1(n_34),
.B2(n_44),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_120),
.B1(n_72),
.B2(n_59),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_48),
.A2(n_20),
.B1(n_31),
.B2(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_114),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_113),
.B(n_12),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_45),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_54),
.A2(n_44),
.B1(n_45),
.B2(n_33),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_62),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_52),
.A2(n_31),
.B1(n_20),
.B2(n_24),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_57),
.A2(n_31),
.B1(n_18),
.B2(n_24),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_64),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_138),
.B1(n_8),
.B2(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_91),
.Y(n_158)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_90),
.C(n_88),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_11),
.Y(n_187)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_46),
.Y(n_137)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_68),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_83),
.B(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_62),
.Y(n_160)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_147),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_82),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_150),
.B(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_151),
.A2(n_153),
.B1(n_167),
.B2(n_168),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_71),
.B1(n_87),
.B2(n_79),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_159),
.B1(n_173),
.B2(n_138),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_100),
.A2(n_70),
.B1(n_78),
.B2(n_77),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_105),
.A2(n_89),
.B1(n_69),
.B2(n_49),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_155),
.A2(n_171),
.B1(n_179),
.B2(n_13),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_158),
.B(n_160),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_92),
.A2(n_91),
.B1(n_67),
.B2(n_25),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_162),
.B(n_176),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_163),
.A2(n_184),
.B1(n_13),
.B2(n_14),
.Y(n_234)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_165),
.Y(n_242)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_60),
.B1(n_25),
.B2(n_5),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_60),
.B1(n_25),
.B2(n_5),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_169),
.Y(n_239)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_171)
);

NAND2x1_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_25),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_172),
.B(n_177),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_99),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_7),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_101),
.B(n_7),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_115),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_112),
.B(n_8),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_191),
.B1(n_118),
.B2(n_136),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_108),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_109),
.B(n_118),
.Y(n_222)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_119),
.B(n_11),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_193),
.Y(n_232)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_14),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_134),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_132),
.C(n_122),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_202),
.B(n_217),
.C(n_226),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_140),
.B1(n_115),
.B2(n_117),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_206),
.A2(n_241),
.B1(n_194),
.B2(n_166),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_209),
.B(n_234),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_128),
.C(n_109),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_140),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_228),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_229),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_159),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_117),
.C(n_123),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_143),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_143),
.C(n_141),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_124),
.B(n_141),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_231),
.B(n_172),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_177),
.A2(n_13),
.B(n_14),
.C(n_157),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_147),
.B1(n_192),
.B2(n_154),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_164),
.B(n_175),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_181),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_152),
.A2(n_157),
.B1(n_184),
.B2(n_173),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_245),
.A2(n_259),
.B1(n_265),
.B2(n_284),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_172),
.B(n_196),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_246),
.A2(n_258),
.B(n_271),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_247),
.A2(n_255),
.B1(n_252),
.B2(n_261),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_248),
.A2(n_283),
.B1(n_264),
.B2(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_252),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_253),
.A2(n_237),
.B(n_205),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_223),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_161),
.B1(n_189),
.B2(n_195),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_174),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_260),
.Y(n_293)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

AO21x2_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_193),
.B(n_190),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_161),
.B1(n_174),
.B2(n_188),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_214),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_262),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_263),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_212),
.B(n_148),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_268),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_209),
.A2(n_208),
.B1(n_230),
.B2(n_212),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_148),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_273),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_169),
.B(n_170),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_238),
.B(n_221),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_165),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_208),
.A2(n_149),
.B1(n_165),
.B2(n_216),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_220),
.A2(n_149),
.B(n_217),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_207),
.B(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_214),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_232),
.Y(n_303)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_278),
.Y(n_286)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_234),
.A3(n_222),
.B1(n_235),
.B2(n_227),
.Y(n_280)
);

OAI32xp33_ASAP7_75t_L g319 ( 
.A1(n_280),
.A2(n_272),
.A3(n_284),
.B1(n_258),
.B2(n_266),
.Y(n_319)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_282),
.Y(n_310)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_234),
.A2(n_229),
.B1(n_204),
.B2(n_205),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_234),
.B1(n_243),
.B2(n_218),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_316),
.B1(n_257),
.B2(n_269),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_287),
.B(n_295),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_258),
.A2(n_238),
.B(n_219),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_292),
.B(n_299),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_237),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_301),
.C(n_305),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_219),
.B(n_201),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_294),
.B(n_258),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_242),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_243),
.C(n_200),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_311),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_258),
.A2(n_239),
.B(n_201),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_200),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_303),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_265),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_210),
.B1(n_232),
.B2(n_224),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_306),
.A2(n_258),
.B1(n_259),
.B2(n_249),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_279),
.A2(n_210),
.B(n_267),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_246),
.B(n_210),
.C(n_272),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_283),
.C(n_263),
.Y(n_344)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_255),
.B1(n_247),
.B2(n_268),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_321),
.A2(n_343),
.B1(n_346),
.B2(n_306),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_322),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_316),
.B1(n_285),
.B2(n_299),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_303),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_326),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_328),
.A2(n_342),
.B(n_345),
.Y(n_352)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_275),
.Y(n_331)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_335),
.Y(n_349)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_317),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_303),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_337),
.B(n_341),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_315),
.A2(n_245),
.B1(n_280),
.B2(n_282),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_340),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_276),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_309),
.B(n_278),
.Y(n_341)
);

XOR2x2_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_277),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_348),
.C(n_294),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_263),
.B(n_307),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_295),
.C(n_301),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_360),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_327),
.A2(n_290),
.B1(n_300),
.B2(n_289),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_355),
.A2(n_356),
.B1(n_359),
.B2(n_362),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_334),
.A2(n_289),
.B(n_311),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_348),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_361),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_327),
.A2(n_319),
.B1(n_292),
.B2(n_313),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_308),
.B1(n_307),
.B2(n_298),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_336),
.B(n_298),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_320),
.A2(n_308),
.B1(n_310),
.B2(n_286),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_325),
.A2(n_286),
.B1(n_310),
.B2(n_297),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_363),
.A2(n_370),
.B1(n_337),
.B2(n_326),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_333),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_367),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_324),
.B(n_287),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_344),
.C(n_347),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_297),
.B1(n_302),
.B2(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_349),
.Y(n_373)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_388),
.Y(n_400)
);

A2O1A1O1Ixp25_ASAP7_75t_L g375 ( 
.A1(n_357),
.A2(n_324),
.B(n_340),
.C(n_342),
.D(n_330),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_383),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_346),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_369),
.B(n_314),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_378),
.B(n_389),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_381),
.A2(n_386),
.B1(n_351),
.B2(n_370),
.Y(n_397)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_334),
.B(n_323),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_367),
.Y(n_402)
);

A2O1A1O1Ixp25_ASAP7_75t_L g383 ( 
.A1(n_359),
.A2(n_331),
.B(n_338),
.C(n_329),
.D(n_332),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_355),
.A2(n_343),
.B1(n_339),
.B2(n_335),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_390),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_312),
.C(n_322),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_322),
.C(n_304),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_369),
.C(n_352),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_371),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_391),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_354),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_354),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_384),
.A2(n_364),
.B(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_401),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_364),
.B(n_363),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_396),
.A2(n_398),
.B(n_402),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_397),
.A2(n_404),
.B1(n_366),
.B2(n_353),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_377),
.A2(n_364),
.B(n_371),
.Y(n_398)
);

A2O1A1O1Ixp25_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_380),
.B(n_390),
.C(n_382),
.D(n_361),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_403),
.B(n_407),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_377),
.A2(n_353),
.B1(n_366),
.B2(n_358),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_382),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_396),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_395),
.A2(n_386),
.B1(n_380),
.B2(n_383),
.Y(n_410)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_397),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_387),
.C(n_389),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_402),
.C(n_393),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_394),
.A2(n_379),
.B1(n_385),
.B2(n_399),
.Y(n_413)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_413),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_400),
.A2(n_379),
.B1(n_385),
.B2(n_409),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_418),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_404),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_407),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_419),
.B(n_398),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_420),
.A2(n_419),
.B(n_409),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_405),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_414),
.B(n_408),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_424),
.B(n_428),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_410),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_429),
.A2(n_430),
.B(n_431),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_414),
.A2(n_394),
.B(n_403),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_431),
.B(n_416),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_428),
.A2(n_421),
.B(n_416),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_436),
.B(n_422),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_441),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_SL g440 ( 
.A(n_437),
.B(n_425),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_440),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_427),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_442),
.A2(n_439),
.B(n_434),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_445),
.B(n_415),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_426),
.C(n_423),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_434),
.C(n_412),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_411),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_415),
.Y(n_449)
);


endmodule