module fake_ariane_3244_n_966 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_966);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_966;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_731;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_872;
wire n_933;
wire n_774;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_137),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_55),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_49),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_77),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_11),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_67),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_108),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_18),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_79),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_144),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_24),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_26),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_38),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_88),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_44),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_60),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_13),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_106),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_89),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_158),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_124),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_78),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_63),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_123),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_51),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_56),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_82),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_148),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_91),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_100),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_92),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_41),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_66),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_160),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_87),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_81),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_71),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_135),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_211),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

BUFx6f_ASAP7_75t_SL g278 ( 
.A(n_193),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_212),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_194),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_212),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_193),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_199),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_200),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_257),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_201),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_193),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_197),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_197),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_244),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_250),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_203),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_204),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_190),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_195),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_206),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_196),
.B(n_0),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_207),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_202),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_218),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_225),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_210),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_268),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_R g325 ( 
.A(n_276),
.B(n_281),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_286),
.B(n_243),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_254),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_269),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_284),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_285),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_270),
.B(n_264),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_246),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_277),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_288),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_304),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_R g344 ( 
.A(n_302),
.B(n_305),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_256),
.B(n_253),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_307),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_301),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_318),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_286),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_283),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_318),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_287),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_287),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_279),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_279),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_282),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_278),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_282),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_314),
.B(n_259),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_278),
.Y(n_376)
);

NAND3xp33_ASAP7_75t_L g377 ( 
.A(n_329),
.B(n_306),
.C(n_272),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_296),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_363),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_345),
.B1(n_354),
.B2(n_336),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_296),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_299),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_325),
.B(n_260),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_375),
.A2(n_299),
.B1(n_192),
.B2(n_215),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_213),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_214),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_363),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_219),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_349),
.B(n_371),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_363),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

BUFx4f_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_372),
.A2(n_263),
.B1(n_262),
.B2(n_261),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_217),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_325),
.B(n_219),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_362),
.B(n_221),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_223),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_344),
.B(n_219),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_321),
.B(n_1),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_354),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_L g418 ( 
.A(n_336),
.B(n_226),
.C(n_224),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_319),
.B(n_228),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_360),
.B(n_1),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_343),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_258),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_230),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_233),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_341),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_334),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_352),
.B(n_235),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_353),
.B(n_236),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_344),
.B(n_219),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_338),
.B(n_252),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_335),
.B(n_232),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_355),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_327),
.A2(n_232),
.B1(n_249),
.B2(n_248),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_237),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_337),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_337),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_342),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_350),
.B(n_240),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_356),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_378),
.B(n_2),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_405),
.B(n_232),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_2),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_369),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_370),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_247),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_423),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

NOR2x1p5_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_374),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_3),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_381),
.B(n_368),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_388),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_419),
.A2(n_391),
.B(n_396),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_446),
.B(n_405),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_445),
.B(n_251),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_409),
.B(n_232),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_411),
.A2(n_98),
.B(n_187),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_432),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_445),
.B(n_3),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_383),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_425),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_392),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_410),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_387),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_424),
.B(n_5),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_403),
.B(n_7),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_445),
.B(n_8),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_9),
.Y(n_490)
);

OAI221xp5_ASAP7_75t_L g491 ( 
.A1(n_390),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_377),
.B(n_10),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_427),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_416),
.Y(n_495)
);

BUFx6f_ASAP7_75t_SL g496 ( 
.A(n_451),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_12),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_420),
.B(n_14),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_410),
.A2(n_414),
.B1(n_435),
.B2(n_418),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_399),
.B(n_14),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_426),
.B(n_15),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_436),
.B(n_15),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_436),
.B(n_16),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_16),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_399),
.B(n_17),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_380),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_380),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_420),
.B(n_17),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_420),
.B(n_18),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_19),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_438),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_414),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_415),
.B(n_22),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_23),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_442),
.B(n_23),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_398),
.B(n_24),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_380),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_404),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_25),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_443),
.B(n_25),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_404),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_413),
.B(n_188),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_394),
.B(n_27),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_437),
.B(n_29),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_386),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_447),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_431),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_386),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_37),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_382),
.B(n_186),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_443),
.B(n_444),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_468),
.A2(n_433),
.B(n_434),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_486),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_483),
.A2(n_415),
.B(n_450),
.C(n_431),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_471),
.A2(n_438),
.B(n_439),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_478),
.A2(n_438),
.B(n_439),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_452),
.B(n_397),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_452),
.B(n_415),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_524),
.A2(n_397),
.B(n_393),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_461),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_460),
.A2(n_407),
.B(n_395),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_507),
.A2(n_407),
.B(n_395),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_508),
.A2(n_393),
.B(n_430),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_518),
.A2(n_430),
.B(n_444),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_474),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_455),
.B(n_441),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_519),
.A2(n_523),
.B(n_522),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_464),
.A2(n_406),
.B(n_400),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_529),
.A2(n_417),
.B(n_428),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_455),
.B(n_400),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_400),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_464),
.A2(n_400),
.B(n_428),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_477),
.B(n_428),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_465),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_481),
.B(n_484),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_453),
.A2(n_400),
.B(n_428),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_505),
.B(n_40),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_482),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_477),
.B(n_185),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_489),
.B(n_43),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_503),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_498),
.B(n_48),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_532),
.A2(n_52),
.B(n_53),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_492),
.A2(n_54),
.B(n_57),
.C(n_59),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_517),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_498),
.B(n_61),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_474),
.A2(n_62),
.B(n_64),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_68),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_459),
.A2(n_70),
.B(n_72),
.Y(n_576)
);

A2O1A1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_492),
.A2(n_73),
.B(n_74),
.C(n_76),
.Y(n_577)
);

AO21x1_ASAP7_75t_L g578 ( 
.A1(n_497),
.A2(n_182),
.B(n_84),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_462),
.A2(n_83),
.B(n_85),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_521),
.B(n_86),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_504),
.A2(n_90),
.B1(n_93),
.B2(n_95),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_467),
.A2(n_96),
.B(n_97),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_511),
.B(n_99),
.C(n_101),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_487),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_102),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_528),
.B(n_104),
.Y(n_586)
);

BUFx12f_ASAP7_75t_L g587 ( 
.A(n_463),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_469),
.B(n_181),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_502),
.A2(n_105),
.B(n_107),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_509),
.B(n_109),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_516),
.B(n_110),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_509),
.B(n_111),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_495),
.A2(n_112),
.B(n_113),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_517),
.B(n_114),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_512),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_473),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_540),
.A2(n_542),
.B(n_535),
.Y(n_597)
);

O2A1O1Ixp5_ASAP7_75t_L g598 ( 
.A1(n_585),
.A2(n_540),
.B(n_550),
.C(n_552),
.Y(n_598)
);

OAI21xp33_ASAP7_75t_L g599 ( 
.A1(n_584),
.A2(n_512),
.B(n_564),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_539),
.A2(n_533),
.B(n_470),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_544),
.B(n_534),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_563),
.B(n_515),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_511),
.C(n_491),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_543),
.A2(n_454),
.B(n_514),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_541),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_538),
.A2(n_472),
.B(n_485),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_559),
.A2(n_510),
.B1(n_499),
.B2(n_500),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_563),
.B(n_496),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_551),
.A2(n_490),
.B(n_520),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_558),
.B(n_458),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_557),
.B(n_510),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_562),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

A2O1A1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_526),
.B(n_506),
.C(n_501),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_596),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_536),
.B(n_525),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_545),
.A2(n_494),
.B(n_454),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_553),
.A2(n_526),
.B(n_475),
.Y(n_618)
);

CKINVDCx11_ASAP7_75t_R g619 ( 
.A(n_587),
.Y(n_619)
);

NAND2x1_ASAP7_75t_L g620 ( 
.A(n_549),
.B(n_531),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_537),
.A2(n_480),
.B1(n_513),
.B2(n_501),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_574),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_574),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_537),
.A2(n_488),
.B(n_506),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_546),
.A2(n_530),
.B(n_527),
.Y(n_625)
);

AOI21x1_ASAP7_75t_L g626 ( 
.A1(n_554),
.A2(n_547),
.B(n_556),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_558),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_560),
.A2(n_118),
.B(n_119),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_565),
.A2(n_575),
.B(n_561),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_548),
.A2(n_555),
.B(n_591),
.Y(n_631)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_578),
.A2(n_120),
.B(n_122),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_549),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_590),
.A2(n_496),
.B(n_126),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_576),
.A2(n_125),
.B(n_128),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_570),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_571),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_567),
.B(n_133),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_579),
.A2(n_134),
.B(n_139),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_593),
.A2(n_140),
.B(n_142),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_580),
.A2(n_149),
.B(n_150),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_592),
.A2(n_151),
.B(n_152),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_568),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_588),
.B(n_153),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_595),
.A2(n_154),
.B(n_155),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_573),
.A2(n_157),
.B(n_162),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_567),
.B(n_163),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_594),
.B(n_164),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_628),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_614),
.A2(n_589),
.B1(n_577),
.B2(n_583),
.Y(n_651)
);

AOI21xp33_ASAP7_75t_L g652 ( 
.A1(n_603),
.A2(n_581),
.B(n_566),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_605),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_601),
.B(n_569),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_627),
.B(n_582),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_602),
.B(n_179),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_603),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_612),
.Y(n_658)
);

BUFx2_ASAP7_75t_SL g659 ( 
.A(n_601),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_619),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_597),
.A2(n_168),
.B(n_169),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_637),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_615),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_599),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_610),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_176),
.Y(n_667)
);

AO21x1_ASAP7_75t_L g668 ( 
.A1(n_621),
.A2(n_178),
.B(n_634),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_628),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_622),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_613),
.B(n_633),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_637),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_599),
.A2(n_607),
.B1(n_645),
.B2(n_634),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_637),
.B(n_616),
.Y(n_674)
);

NOR2x1_ASAP7_75t_L g675 ( 
.A(n_611),
.B(n_646),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_608),
.B(n_616),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_613),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_644),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_648),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_644),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_613),
.B(n_620),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_624),
.A2(n_625),
.B1(n_636),
.B2(n_638),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_623),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_644),
.B(n_649),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_642),
.B(n_644),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_629),
.B(n_618),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_609),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_604),
.B(n_642),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_640),
.A2(n_639),
.B1(n_635),
.B2(n_631),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_598),
.B(n_630),
.C(n_600),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

INVx3_ASAP7_75t_SL g692 ( 
.A(n_641),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_617),
.B(n_647),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_606),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_632),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_599),
.B(n_603),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_627),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_605),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_599),
.A2(n_603),
.B(n_452),
.C(n_614),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_678),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_679),
.A2(n_696),
.B1(n_668),
.B2(n_666),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_678),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_691),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_691),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_670),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_699),
.A2(n_673),
.B1(n_651),
.B2(n_697),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_687),
.Y(n_707)
);

BUFx8_ASAP7_75t_SL g708 ( 
.A(n_660),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_686),
.A2(n_682),
.B(n_693),
.Y(n_709)
);

BUFx4f_ASAP7_75t_SL g710 ( 
.A(n_662),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_685),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_658),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_678),
.A2(n_680),
.B1(n_675),
.B2(n_652),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_683),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_SL g715 ( 
.A1(n_657),
.A2(n_675),
.B(n_665),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_666),
.B(n_698),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_694),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_659),
.B(n_654),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_672),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_680),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_677),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_653),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_680),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_671),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_696),
.B(n_676),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_663),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_695),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_674),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_654),
.B(n_684),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_695),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_664),
.B(n_671),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_688),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_671),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_690),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_689),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_690),
.A2(n_689),
.B(n_661),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_681),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_665),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_650),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_656),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_667),
.Y(n_745)
);

BUFx8_ASAP7_75t_SL g746 ( 
.A(n_650),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_657),
.A2(n_603),
.B1(n_357),
.B2(n_368),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_669),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_664),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_669),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_664),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_678),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_691),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_678),
.B(n_680),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_678),
.B(n_680),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_691),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_691),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_686),
.A2(n_626),
.B(n_606),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_738),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_717),
.Y(n_760)
);

AOI21x1_ASAP7_75t_L g761 ( 
.A1(n_713),
.A2(n_738),
.B(n_706),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_733),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_735),
.Y(n_763)
);

AO21x1_ASAP7_75t_L g764 ( 
.A1(n_715),
.A2(n_742),
.B(n_701),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_711),
.B(n_716),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_708),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_733),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_729),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_722),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_740),
.A2(n_758),
.B(n_709),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_722),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_729),
.B(n_718),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_705),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_724),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_724),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_740),
.A2(n_758),
.B(n_709),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_721),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_707),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_721),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_735),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_714),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_754),
.B(n_718),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_724),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_707),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_704),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_716),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_739),
.A2(n_727),
.B(n_730),
.Y(n_787)
);

OA21x2_ASAP7_75t_L g788 ( 
.A1(n_742),
.A2(n_739),
.B(n_703),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_729),
.B(n_718),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_737),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_729),
.B(n_718),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_703),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_725),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_753),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_711),
.B(n_725),
.Y(n_795)
);

AO21x2_ASAP7_75t_L g796 ( 
.A1(n_727),
.A2(n_730),
.B(n_756),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_753),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_756),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_704),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_757),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_757),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_726),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_760),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_766),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_759),
.B(n_790),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_777),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_765),
.A2(n_747),
.B1(n_712),
.B2(n_745),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_795),
.B(n_793),
.Y(n_808)
);

OA21x2_ASAP7_75t_L g809 ( 
.A1(n_770),
.A2(n_744),
.B(n_748),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_769),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_769),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_778),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_783),
.Y(n_813)
);

NOR4xp25_ASAP7_75t_SL g814 ( 
.A(n_766),
.B(n_712),
.C(n_736),
.D(n_734),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_771),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_780),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_795),
.B(n_744),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_780),
.B(n_750),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_L g819 ( 
.A1(n_764),
.A2(n_732),
.B1(n_719),
.B2(n_728),
.C(n_748),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_770),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_771),
.Y(n_821)
);

INVxp67_ASAP7_75t_SL g822 ( 
.A(n_800),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_792),
.Y(n_823)
);

AND2x4_ASAP7_75t_SL g824 ( 
.A(n_782),
.B(n_755),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_759),
.B(n_750),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_792),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_784),
.B(n_719),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_765),
.B(n_743),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_773),
.Y(n_829)
);

OAI221xp5_ASAP7_75t_L g830 ( 
.A1(n_761),
.A2(n_741),
.B1(n_754),
.B2(n_751),
.C(n_700),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_773),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_781),
.Y(n_832)
);

AOI211xp5_ASAP7_75t_SL g833 ( 
.A1(n_764),
.A2(n_700),
.B(n_752),
.C(n_755),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_786),
.B(n_743),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_785),
.B(n_743),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_776),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_805),
.B(n_763),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_805),
.B(n_763),
.Y(n_838)
);

AOI221xp5_ASAP7_75t_L g839 ( 
.A1(n_807),
.A2(n_819),
.B1(n_802),
.B2(n_832),
.C(n_831),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_812),
.B(n_822),
.Y(n_840)
);

AOI211xp5_ASAP7_75t_L g841 ( 
.A1(n_807),
.A2(n_802),
.B(n_777),
.C(n_779),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_SL g842 ( 
.A1(n_833),
.A2(n_761),
.B(n_785),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_808),
.B(n_779),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_817),
.B(n_786),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_817),
.B(n_816),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_804),
.B(n_708),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_816),
.B(n_801),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_830),
.A2(n_791),
.B1(n_772),
.B2(n_789),
.Y(n_848)
);

NAND4xp25_ASAP7_75t_L g849 ( 
.A(n_835),
.B(n_799),
.C(n_801),
.D(n_797),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_833),
.B(n_799),
.C(n_794),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_828),
.B(n_798),
.Y(n_851)
);

OA21x2_ASAP7_75t_L g852 ( 
.A1(n_823),
.A2(n_776),
.B(n_787),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_828),
.B(n_827),
.Y(n_853)
);

AND2x2_ASAP7_75t_SL g854 ( 
.A(n_824),
.B(n_791),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_803),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_808),
.B(n_772),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_818),
.B(n_798),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_806),
.B(n_789),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_L g859 ( 
.A(n_834),
.B(n_797),
.C(n_794),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_818),
.B(n_825),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_825),
.B(n_788),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_SL g862 ( 
.A1(n_835),
.A2(n_772),
.B(n_791),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_806),
.B(n_788),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_823),
.B(n_788),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_864),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_843),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_837),
.B(n_821),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_856),
.B(n_860),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_845),
.B(n_806),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_852),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_862),
.B(n_823),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_837),
.B(n_821),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_838),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_861),
.B(n_826),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_838),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_858),
.B(n_850),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_853),
.B(n_826),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_852),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_857),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_851),
.B(n_826),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_844),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_855),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_881),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_874),
.B(n_849),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_881),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_877),
.A2(n_841),
.B1(n_839),
.B2(n_842),
.Y(n_887)
);

NOR2x1_ASAP7_75t_L g888 ( 
.A(n_877),
.B(n_846),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_867),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_873),
.Y(n_890)
);

AND3x2_ASAP7_75t_L g891 ( 
.A(n_877),
.B(n_755),
.C(n_731),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_876),
.B(n_847),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_880),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_868),
.B(n_859),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_890),
.B(n_865),
.Y(n_895)
);

OAI33xp33_ASAP7_75t_L g896 ( 
.A1(n_887),
.A2(n_865),
.A3(n_875),
.B1(n_879),
.B2(n_871),
.B3(n_863),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_885),
.B(n_882),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_894),
.B(n_875),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_893),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_884),
.B(n_878),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_889),
.B(n_872),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_888),
.B(n_869),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_889),
.B(n_872),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_886),
.B(n_869),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_892),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_902),
.B(n_878),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_905),
.B(n_891),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_899),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_897),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_904),
.B(n_870),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_908),
.B(n_901),
.C(n_903),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_909),
.B(n_898),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_907),
.Y(n_913)
);

AOI21xp33_ASAP7_75t_L g914 ( 
.A1(n_906),
.A2(n_895),
.B(n_879),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_912),
.B(n_910),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_911),
.B(n_910),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_913),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_914),
.A2(n_896),
.B1(n_871),
.B2(n_895),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_913),
.A2(n_848),
.B1(n_900),
.B2(n_789),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_915),
.B(n_866),
.Y(n_920)
);

NAND4xp25_ASAP7_75t_L g921 ( 
.A(n_916),
.B(n_870),
.C(n_820),
.D(n_836),
.Y(n_921)
);

AOI211xp5_ASAP7_75t_L g922 ( 
.A1(n_917),
.A2(n_918),
.B(n_919),
.C(n_813),
.Y(n_922)
);

AOI322xp5_ASAP7_75t_L g923 ( 
.A1(n_918),
.A2(n_864),
.A3(n_883),
.B1(n_854),
.B2(n_810),
.C1(n_815),
.C2(n_811),
.Y(n_923)
);

AOI221x1_ASAP7_75t_L g924 ( 
.A1(n_917),
.A2(n_820),
.B1(n_836),
.B2(n_815),
.C(n_810),
.Y(n_924)
);

AOI211x1_ASAP7_75t_L g925 ( 
.A1(n_916),
.A2(n_811),
.B(n_829),
.C(n_831),
.Y(n_925)
);

NAND5xp2_ASAP7_75t_L g926 ( 
.A(n_916),
.B(n_746),
.C(n_754),
.D(n_814),
.E(n_710),
.Y(n_926)
);

NAND4xp25_ASAP7_75t_L g927 ( 
.A(n_916),
.B(n_836),
.C(n_820),
.D(n_746),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_925),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_922),
.B(n_883),
.C(n_749),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_927),
.B(n_702),
.C(n_720),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_920),
.B(n_883),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_L g932 ( 
.A(n_926),
.B(n_702),
.C(n_720),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_923),
.B(n_883),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_928),
.B(n_924),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_931),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_929),
.B(n_921),
.C(n_702),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_933),
.B(n_883),
.C(n_820),
.Y(n_937)
);

NAND5xp2_ASAP7_75t_L g938 ( 
.A(n_932),
.B(n_814),
.C(n_832),
.D(n_829),
.E(n_813),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_930),
.B(n_836),
.C(n_809),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_934),
.A2(n_809),
.B1(n_813),
.B2(n_723),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_935),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_937),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_938),
.B(n_939),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_936),
.Y(n_944)
);

NOR2x1_ASAP7_75t_L g945 ( 
.A(n_941),
.B(n_720),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_943),
.A2(n_809),
.B1(n_813),
.B2(n_723),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_942),
.B(n_940),
.Y(n_947)
);

NOR4xp75_ASAP7_75t_SL g948 ( 
.A(n_944),
.B(n_813),
.C(n_723),
.D(n_775),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_945),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_947),
.Y(n_950)
);

XOR2xp5_ASAP7_75t_L g951 ( 
.A(n_946),
.B(n_731),
.Y(n_951)
);

AO22x2_ASAP7_75t_L g952 ( 
.A1(n_950),
.A2(n_948),
.B1(n_751),
.B2(n_741),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_951),
.A2(n_809),
.B1(n_813),
.B2(n_731),
.Y(n_953)
);

NAND4xp25_ASAP7_75t_L g954 ( 
.A(n_953),
.B(n_949),
.C(n_775),
.D(n_774),
.Y(n_954)
);

NAND4xp25_ASAP7_75t_L g955 ( 
.A(n_952),
.B(n_775),
.C(n_774),
.D(n_752),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_954),
.A2(n_700),
.B1(n_752),
.B2(n_774),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_956),
.B(n_955),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_783),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_957),
.A2(n_783),
.B1(n_724),
.B2(n_789),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_958),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_960),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_959),
.A2(n_724),
.B1(n_783),
.B2(n_782),
.Y(n_962)
);

AOI222xp33_ASAP7_75t_L g963 ( 
.A1(n_961),
.A2(n_791),
.B1(n_772),
.B2(n_824),
.C1(n_762),
.C2(n_767),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_962),
.A2(n_762),
.B1(n_767),
.B2(n_796),
.Y(n_964)
);

OAI221xp5_ASAP7_75t_R g965 ( 
.A1(n_964),
.A2(n_824),
.B1(n_783),
.B2(n_782),
.C(n_768),
.Y(n_965)
);

AOI211xp5_ASAP7_75t_L g966 ( 
.A1(n_965),
.A2(n_963),
.B(n_768),
.C(n_781),
.Y(n_966)
);


endmodule