module fake_jpeg_18363_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_7),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_71),
.Y(n_81)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_2),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_45),
.B1(n_51),
.B2(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_79),
.B1(n_82),
.B2(n_58),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_59),
.C(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_45),
.B1(n_66),
.B2(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_62),
.B1(n_59),
.B2(n_54),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_56),
.B1(n_29),
.B2(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_58),
.B1(n_60),
.B2(n_50),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_84),
.B1(n_44),
.B2(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_75),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_3),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_15),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_23),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_96),
.A2(n_63),
.B1(n_52),
.B2(n_48),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_19),
.B1(n_42),
.B2(n_8),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_4),
.B(n_5),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_111),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_115),
.B(n_117),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_17),
.C(n_18),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_114),
.C(n_115),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_123),
.B(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_109),
.C(n_98),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_110),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_107),
.C(n_106),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_109),
.A3(n_119),
.B1(n_35),
.B2(n_36),
.C1(n_32),
.C2(n_41),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_33),
.C(n_38),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_43),
.Y(n_132)
);


endmodule