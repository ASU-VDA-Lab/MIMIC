module fake_jpeg_9977_n_37 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_14),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_3),
.Y(n_21)
);

NAND2xp33_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_13),
.B1(n_5),
.B2(n_10),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_1),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_R g27 ( 
.A(n_19),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_28),
.CI(n_30),
.CON(n_32),
.SN(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_23),
.C(n_21),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_32),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_16),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_12),
.B(n_20),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_15),
.B(n_16),
.Y(n_37)
);


endmodule