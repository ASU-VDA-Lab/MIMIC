module fake_aes_4381_n_7 (n_1, n_0, n_7);
input n_1;
input n_0;
output n_7;
wire n_2;
wire n_6;
wire n_4;
wire n_3;
wire n_5;
INVx2_ASAP7_75t_L g2 ( .A(n_0), .Y(n_2) );
OR2x6_ASAP7_75t_L g3 ( .A(n_1), .B(n_0), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
OAI22xp5_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_1), .B1(n_3), .B2(n_2), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_5), .B(n_3), .Y(n_6) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_6), .Y(n_7) );
endmodule