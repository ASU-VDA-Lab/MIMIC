module fake_ibex_198_n_998 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_998);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_998;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_510;
wire n_947;
wire n_972;
wire n_845;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_357;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_375;
wire n_280;
wire n_317;
wire n_340;
wire n_698;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_506;
wire n_444;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_955;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_885;
wire n_588;
wire n_212;
wire n_513;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_921;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_179),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_22),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_56),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_17),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_152),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_160),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_47),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_138),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_49),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_78),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_96),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_21),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_117),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_85),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_66),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_38),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_113),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_60),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_94),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_91),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_146),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_172),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_30),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_42),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_95),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_126),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_136),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_144),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_163),
.B(n_2),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_102),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_176),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_40),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_67),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_86),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_70),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_38),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_116),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_89),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_120),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_174),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_26),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_157),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_88),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_59),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_158),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_13),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_99),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_159),
.B(n_101),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_105),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_173),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_162),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_98),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_43),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_73),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_77),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_178),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_48),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_10),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_177),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_124),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_186),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_169),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_58),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_16),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_30),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_92),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_155),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_151),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_74),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_188),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_93),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_183),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_65),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_53),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_129),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_80),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_182),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_79),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_32),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_20),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_3),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_32),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_197),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_197),
.B(n_0),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_238),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_197),
.Y(n_321)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_212),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_211),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_252),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_274),
.A2(n_97),
.B(n_194),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_197),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_260),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_237),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_246),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_274),
.A2(n_100),
.B(n_193),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_234),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_338)
);

OAI22x1_ASAP7_75t_L g339 ( 
.A1(n_260),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_9),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_273),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_286),
.A2(n_104),
.B(n_192),
.Y(n_343)
);

BUFx8_ASAP7_75t_L g344 ( 
.A(n_197),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_265),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

OAI22x1_ASAP7_75t_R g347 ( 
.A1(n_290),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_197),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_275),
.Y(n_349)
);

BUFx8_ASAP7_75t_L g350 ( 
.A(n_255),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_200),
.B(n_12),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_14),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_214),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_198),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_360)
);

OAI21x1_ASAP7_75t_L g361 ( 
.A1(n_286),
.A2(n_107),
.B(n_185),
.Y(n_361)
);

CKINVDCx11_ASAP7_75t_R g362 ( 
.A(n_313),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_300),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_201),
.Y(n_364)
);

BUFx12f_ASAP7_75t_L g365 ( 
.A(n_196),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_198),
.A2(n_270),
.B1(n_249),
.B2(n_232),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_212),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_226),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_245),
.B(n_15),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_200),
.B(n_19),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_218),
.B(n_19),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_199),
.B(n_20),
.Y(n_374)
);

BUFx8_ASAP7_75t_L g375 ( 
.A(n_255),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_235),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_245),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_248),
.Y(n_379)
);

OAI22x1_ASAP7_75t_L g380 ( 
.A1(n_259),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_218),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_255),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_304),
.A2(n_109),
.B(n_180),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_304),
.A2(n_108),
.B(n_175),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_209),
.A2(n_106),
.B(n_171),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_255),
.Y(n_386)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_301),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_301),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_261),
.B(n_23),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_257),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_344),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_388),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_381),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_388),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_250),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

BUFx6f_ASAP7_75t_SL g398 ( 
.A(n_370),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_277),
.B1(n_312),
.B2(n_298),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_250),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_352),
.B(n_371),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_388),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_316),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_350),
.B(n_255),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_360),
.A2(n_249),
.B1(n_270),
.B2(n_284),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_326),
.A2(n_203),
.B1(n_206),
.B2(n_208),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_324),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_266),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_324),
.Y(n_424)
);

OR2x6_ASAP7_75t_L g425 ( 
.A(n_338),
.B(n_288),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_L g426 ( 
.A(n_352),
.B(n_255),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_324),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_378),
.B(n_315),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_217),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_322),
.A2(n_297),
.B1(n_267),
.B2(n_276),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_375),
.B(n_370),
.Y(n_435)
);

AND3x2_ASAP7_75t_L g436 ( 
.A(n_347),
.B(n_221),
.C(n_219),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_375),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_375),
.B(n_348),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_223),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_377),
.B(n_224),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_325),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_325),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_367),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_336),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_387),
.B(n_227),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_371),
.B(n_254),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_322),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_318),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_387),
.B(n_233),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_387),
.B(n_239),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_387),
.B(n_241),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_336),
.B(n_244),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_318),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_345),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_318),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_387),
.B(n_251),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_349),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_323),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_323),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_323),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_323),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_355),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_372),
.B(n_202),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_365),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_365),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_328),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_342),
.B(n_351),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_351),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_328),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_351),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_358),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_328),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_328),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_358),
.B(n_204),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_328),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_319),
.A2(n_283),
.B1(n_302),
.B2(n_280),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_317),
.B(n_264),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_337),
.B(n_305),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_329),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_329),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_337),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_329),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_329),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_343),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_329),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_331),
.Y(n_500)
);

AND3x2_ASAP7_75t_L g501 ( 
.A(n_339),
.B(n_307),
.C(n_306),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_343),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_361),
.B(n_279),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_331),
.B(n_205),
.Y(n_504)
);

AND3x2_ASAP7_75t_L g505 ( 
.A(n_339),
.B(n_24),
.C(n_25),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_362),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_361),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_402),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_403),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_407),
.A2(n_334),
.B1(n_380),
.B2(n_207),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_403),
.B(n_220),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_383),
.C(n_330),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_411),
.A2(n_222),
.B(n_242),
.C(n_213),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_460),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_391),
.B(n_216),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_407),
.A2(n_380),
.B1(n_225),
.B2(n_285),
.Y(n_522)
);

OAI221xp5_ASAP7_75t_L g523 ( 
.A1(n_400),
.A2(n_393),
.B1(n_457),
.B2(n_488),
.C(n_419),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_391),
.B(n_228),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_457),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_398),
.A2(n_384),
.B1(n_383),
.B2(n_330),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_437),
.B(n_229),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_230),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_477),
.B(n_362),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_460),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_431),
.B(n_331),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_398),
.A2(n_384),
.B1(n_383),
.B2(n_330),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_477),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_425),
.A2(n_385),
.B1(n_384),
.B2(n_311),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_437),
.B(n_231),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_460),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_464),
.B(n_236),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_431),
.B(n_240),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_456),
.B(n_243),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_423),
.B(n_253),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_480),
.Y(n_543)
);

AO22x2_ASAP7_75t_L g544 ( 
.A1(n_420),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_428),
.B(n_256),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_422),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_506),
.A2(n_414),
.B1(n_397),
.B2(n_404),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_478),
.B(n_376),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_430),
.B(n_262),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_425),
.A2(n_293),
.B1(n_268),
.B2(n_269),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_441),
.B(n_263),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_445),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_449),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_454),
.B(n_27),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_434),
.B(n_272),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_435),
.B(n_278),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_503),
.A2(n_376),
.B(n_373),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_465),
.B(n_281),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_435),
.B(n_282),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_447),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_491),
.B(n_287),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_398),
.B(n_289),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_456),
.B(n_291),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_454),
.B(n_292),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_484),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_396),
.B(n_294),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_406),
.B(n_295),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_303),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_410),
.A2(n_503),
.B1(n_425),
.B2(n_507),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_492),
.B(n_335),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_467),
.B(n_308),
.Y(n_576)
);

OAI22x1_ASAP7_75t_SL g577 ( 
.A1(n_436),
.A2(n_309),
.B1(n_310),
.B2(n_31),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_335),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_490),
.A2(n_376),
.B1(n_373),
.B2(n_363),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_335),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_426),
.A2(n_376),
.B1(n_373),
.B2(n_363),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_456),
.B(n_44),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_426),
.A2(n_376),
.B1(n_373),
.B2(n_363),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_409),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_456),
.B(n_28),
.Y(n_586)
);

OAI221xp5_ASAP7_75t_L g587 ( 
.A1(n_483),
.A2(n_373),
.B1(n_363),
.B2(n_357),
.C(n_346),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_492),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_425),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_498),
.B(n_340),
.Y(n_590)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_440),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_439),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_440),
.B(n_340),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_498),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_412),
.B(n_346),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_412),
.B(n_346),
.Y(n_596)
);

O2A1O1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_413),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_440),
.B(n_346),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_440),
.B(n_498),
.Y(n_599)
);

OAI221xp5_ASAP7_75t_L g600 ( 
.A1(n_413),
.A2(n_363),
.B1(n_357),
.B2(n_346),
.C(n_37),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_415),
.B(n_416),
.Y(n_601)
);

AND2x6_ASAP7_75t_SL g602 ( 
.A(n_505),
.B(n_34),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_501),
.B(n_35),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_502),
.A2(n_357),
.B(n_118),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_502),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_590),
.A2(n_469),
.B(n_463),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_455),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_523),
.A2(n_446),
.B1(n_453),
.B2(n_451),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_590),
.A2(n_469),
.B(n_463),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_525),
.B(n_417),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_588),
.A2(n_462),
.B(n_461),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_599),
.A2(n_455),
.B(n_417),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_554),
.A2(n_438),
.B1(n_451),
.B2(n_450),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_591),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_516),
.A2(n_444),
.B(n_418),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_515),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_564),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_585),
.A2(n_433),
.B1(n_450),
.B2(n_448),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_541),
.B(n_433),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_534),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_564),
.A2(n_592),
.B1(n_514),
.B2(n_512),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_516),
.A2(n_438),
.B(n_444),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_526),
.A2(n_533),
.B(n_558),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_541),
.A2(n_446),
.B1(n_504),
.B2(n_392),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_529),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_522),
.B(n_36),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_508),
.A2(n_509),
.B(n_562),
.C(n_553),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_567),
.B(n_36),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_565),
.B(n_392),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_566),
.A2(n_394),
.B1(n_395),
.B2(n_405),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_594),
.A2(n_394),
.B(n_395),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_511),
.A2(n_405),
.B(n_408),
.C(n_500),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_559),
.B(n_43),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_512),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_517),
.B(n_408),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_566),
.B(n_551),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_591),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_551),
.B(n_45),
.Y(n_643)
);

OR2x6_ASAP7_75t_SL g644 ( 
.A(n_530),
.B(n_51),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_513),
.A2(n_474),
.B(n_497),
.C(n_496),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_532),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_605),
.A2(n_535),
.B(n_601),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_549),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_548),
.B(n_52),
.Y(n_649)
);

O2A1O1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_573),
.A2(n_497),
.B(n_496),
.C(n_494),
.Y(n_650)
);

BUFx12f_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_521),
.B(n_54),
.Y(n_652)
);

OAI21xp33_ASAP7_75t_L g653 ( 
.A1(n_548),
.A2(n_473),
.B(n_459),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_573),
.B(n_399),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_597),
.A2(n_489),
.B(n_486),
.C(n_485),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_518),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_550),
.B(n_55),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_569),
.A2(n_479),
.B(n_468),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_586),
.B(n_57),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_549),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_570),
.A2(n_482),
.B(n_471),
.Y(n_662)
);

AO21x1_ASAP7_75t_L g663 ( 
.A1(n_604),
.A2(n_489),
.B(n_486),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_572),
.B(n_61),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_532),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_552),
.B(n_62),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_528),
.B(n_63),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_530),
.B(n_64),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_542),
.A2(n_472),
.B(n_493),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_545),
.A2(n_539),
.B(n_576),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_68),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_561),
.B(n_72),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_583),
.A2(n_499),
.B1(n_493),
.B2(n_466),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_532),
.Y(n_675)
);

NOR2x1_ASAP7_75t_L g676 ( 
.A(n_555),
.B(n_499),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_563),
.B(n_76),
.Y(n_677)
);

NAND2x1p5_ASAP7_75t_L g678 ( 
.A(n_524),
.B(n_466),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_580),
.B(n_399),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_527),
.B(n_81),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_536),
.B(n_83),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_520),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_556),
.A2(n_84),
.B1(n_87),
.B2(n_90),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_540),
.B(n_195),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_531),
.B(n_538),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_568),
.B(n_110),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_589),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_571),
.A2(n_115),
.B(n_119),
.C(n_122),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_575),
.A2(n_125),
.B(n_128),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_575),
.B(n_168),
.Y(n_690)
);

OAI21xp33_ASAP7_75t_L g691 ( 
.A1(n_579),
.A2(n_131),
.B(n_133),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_639),
.B(n_603),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_656),
.B(n_544),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_646),
.B(n_544),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_641),
.B(n_577),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_639),
.B(n_602),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_618),
.A2(n_595),
.B(n_596),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_612),
.B(n_581),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_608),
.B(n_633),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_619),
.B(n_593),
.Y(n_700)
);

AO21x1_ASAP7_75t_L g701 ( 
.A1(n_654),
.A2(n_598),
.B(n_600),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_652),
.A2(n_584),
.B1(n_582),
.B2(n_587),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_627),
.A2(n_134),
.B(n_135),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_620),
.B(n_137),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_651),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_644),
.B(n_139),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_623),
.B(n_632),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_660),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_671),
.B(n_147),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_627),
.A2(n_148),
.B(n_149),
.Y(n_710)
);

NAND2x1p5_ASAP7_75t_L g711 ( 
.A(n_660),
.B(n_150),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_675),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_R g713 ( 
.A(n_624),
.B(n_153),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_617),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_648),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_626),
.B(n_154),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_669),
.B(n_164),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_638),
.B(n_167),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_609),
.B(n_165),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_609),
.B(n_166),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_631),
.B(n_630),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_648),
.Y(n_722)
);

AOI21xp33_ASAP7_75t_L g723 ( 
.A1(n_655),
.A2(n_653),
.B(n_643),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_642),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_606),
.B(n_642),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_647),
.A2(n_614),
.B(n_610),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_684),
.B(n_659),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_682),
.Y(n_728)
);

OAI21x1_ASAP7_75t_SL g729 ( 
.A1(n_689),
.A2(n_675),
.B(n_680),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_615),
.A2(n_687),
.B1(n_649),
.B2(n_640),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_684),
.A2(n_673),
.B1(n_681),
.B2(n_635),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_622),
.A2(n_670),
.B(n_650),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_616),
.B(n_625),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_646),
.B(n_665),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_637),
.A2(n_607),
.B(n_611),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_665),
.Y(n_736)
);

NOR2x1_ASAP7_75t_SL g737 ( 
.A(n_672),
.B(n_621),
.Y(n_737)
);

OA22x2_ASAP7_75t_L g738 ( 
.A1(n_689),
.A2(n_629),
.B1(n_634),
.B2(n_683),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_616),
.B(n_685),
.Y(n_739)
);

NOR2x1_ASAP7_75t_SL g740 ( 
.A(n_690),
.B(n_664),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_678),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_657),
.B(n_667),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_678),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_676),
.B(n_661),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_663),
.A2(n_636),
.B(n_686),
.Y(n_745)
);

OA21x2_ASAP7_75t_L g746 ( 
.A1(n_691),
.A2(n_645),
.B(n_679),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_661),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_SL g748 ( 
.A1(n_677),
.A2(n_668),
.B(n_688),
.C(n_674),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_613),
.A2(n_662),
.B(n_658),
.Y(n_749)
);

CKINVDCx11_ASAP7_75t_R g750 ( 
.A(n_651),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_639),
.B(n_391),
.Y(n_751)
);

CKINVDCx11_ASAP7_75t_R g752 ( 
.A(n_651),
.Y(n_752)
);

OA21x2_ASAP7_75t_L g753 ( 
.A1(n_628),
.A2(n_516),
.B(n_503),
.Y(n_753)
);

OAI21x1_ASAP7_75t_SL g754 ( 
.A1(n_689),
.A2(n_675),
.B(n_671),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_671),
.A2(n_632),
.B(n_655),
.C(n_657),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_652),
.A2(n_641),
.B1(n_612),
.B2(n_643),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_628),
.A2(n_654),
.B(n_653),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_628),
.A2(n_627),
.B(n_618),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_SL g759 ( 
.A1(n_675),
.A2(n_689),
.B(n_588),
.Y(n_759)
);

AO32x2_ASAP7_75t_L g760 ( 
.A1(n_626),
.A2(n_535),
.A3(n_610),
.B1(n_674),
.B2(n_615),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_608),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_671),
.A2(n_632),
.B(n_655),
.C(n_657),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_639),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_671),
.A2(n_590),
.B(n_588),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_656),
.B(n_666),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_656),
.B(n_666),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_608),
.B(n_543),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_671),
.A2(n_632),
.B(n_655),
.C(n_657),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_628),
.A2(n_627),
.B(n_618),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_660),
.B(n_639),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_641),
.B(n_578),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_656),
.B(n_666),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_639),
.B(n_543),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_543),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_619),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_775),
.Y(n_776)
);

AOI221xp5_ASAP7_75t_L g777 ( 
.A1(n_771),
.A2(n_756),
.B1(n_693),
.B2(n_699),
.C(n_695),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_727),
.B(n_763),
.Y(n_778)
);

AO21x2_ASAP7_75t_L g779 ( 
.A1(n_758),
.A2(n_769),
.B(n_729),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_767),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_763),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_750),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_752),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_705),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_761),
.B(n_774),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_694),
.A2(n_706),
.B1(n_713),
.B2(n_693),
.Y(n_786)
);

AO21x2_ASAP7_75t_L g787 ( 
.A1(n_723),
.A2(n_726),
.B(n_754),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_765),
.B(n_766),
.Y(n_788)
);

INVx6_ASAP7_75t_L g789 ( 
.A(n_700),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_766),
.B(n_772),
.Y(n_790)
);

AO22x2_ASAP7_75t_L g791 ( 
.A1(n_730),
.A2(n_694),
.B1(n_724),
.B2(n_773),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_772),
.B(n_714),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_728),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_696),
.B(n_692),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_721),
.A2(n_716),
.B1(n_707),
.B2(n_731),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_770),
.Y(n_796)
);

OA21x2_ASAP7_75t_L g797 ( 
.A1(n_745),
.A2(n_732),
.B(n_735),
.Y(n_797)
);

AO31x2_ASAP7_75t_L g798 ( 
.A1(n_701),
.A2(n_740),
.A3(n_709),
.B(n_764),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_725),
.A2(n_751),
.B(n_742),
.C(n_722),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_736),
.B(n_712),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_715),
.A2(n_719),
.B1(n_720),
.B2(n_704),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_747),
.A2(n_724),
.B1(n_717),
.B2(n_708),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_770),
.Y(n_803)
);

AO32x2_ASAP7_75t_L g804 ( 
.A1(n_757),
.A2(n_702),
.A3(n_760),
.B1(n_736),
.B2(n_753),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_738),
.A2(n_753),
.B(n_697),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_698),
.Y(n_806)
);

AO32x2_ASAP7_75t_L g807 ( 
.A1(n_757),
.A2(n_702),
.A3(n_760),
.B1(n_738),
.B2(n_759),
.Y(n_807)
);

AO32x2_ASAP7_75t_L g808 ( 
.A1(n_760),
.A2(n_746),
.A3(n_703),
.B1(n_710),
.B2(n_711),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_708),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_712),
.B(n_743),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_711),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_741),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_739),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_746),
.A2(n_734),
.B(n_744),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_733),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_718),
.B(n_737),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_761),
.B(n_510),
.Y(n_817)
);

AO31x2_ASAP7_75t_L g818 ( 
.A1(n_755),
.A2(n_762),
.A3(n_768),
.B(n_701),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_771),
.B(n_578),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_705),
.B(n_651),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_761),
.B(n_510),
.Y(n_821)
);

BUFx12f_ASAP7_75t_L g822 ( 
.A(n_750),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_771),
.A2(n_641),
.B1(n_554),
.B2(n_420),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_727),
.B(n_763),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_765),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_765),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_756),
.A2(n_366),
.B1(n_530),
.B2(n_420),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_767),
.B(n_771),
.Y(n_828)
);

AO31x2_ASAP7_75t_L g829 ( 
.A1(n_755),
.A2(n_762),
.A3(n_768),
.B(n_701),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_771),
.B(n_641),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_750),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_767),
.B(n_771),
.Y(n_832)
);

AOI22x1_ASAP7_75t_L g833 ( 
.A1(n_754),
.A2(n_729),
.B1(n_711),
.B2(n_749),
.Y(n_833)
);

CKINVDCx6p67_ASAP7_75t_R g834 ( 
.A(n_775),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_748),
.A2(n_762),
.B(n_755),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_750),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_771),
.A2(n_554),
.B(n_565),
.Y(n_837)
);

AO21x2_ASAP7_75t_L g838 ( 
.A1(n_758),
.A2(n_769),
.B(n_729),
.Y(n_838)
);

BUFx8_ASAP7_75t_L g839 ( 
.A(n_705),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_694),
.A2(n_771),
.B1(n_641),
.B2(n_756),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_761),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_771),
.B(n_641),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_727),
.B(n_763),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_771),
.B(n_578),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_705),
.B(n_651),
.Y(n_845)
);

CKINVDCx11_ASAP7_75t_R g846 ( 
.A(n_822),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_SL g847 ( 
.A1(n_811),
.A2(n_803),
.B(n_827),
.C(n_826),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_784),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_788),
.B(n_790),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_841),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_839),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_777),
.B(n_835),
.C(n_833),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_825),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_790),
.B(n_826),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_806),
.B(n_793),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_792),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_L g858 ( 
.A1(n_819),
.A2(n_844),
.B1(n_830),
.B2(n_842),
.C(n_840),
.Y(n_858)
);

CKINVDCx6p67_ASAP7_75t_R g859 ( 
.A(n_834),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_780),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_839),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_828),
.B(n_832),
.Y(n_862)
);

AO31x2_ASAP7_75t_L g863 ( 
.A1(n_816),
.A2(n_812),
.A3(n_818),
.B(n_829),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_810),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_809),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_815),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_814),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_785),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_817),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_795),
.B(n_843),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_800),
.B(n_810),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_791),
.B(n_778),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_786),
.A2(n_823),
.B1(n_801),
.B2(n_837),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_831),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_824),
.A2(n_789),
.B1(n_794),
.B2(n_821),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_813),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_804),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_779),
.B(n_838),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_779),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_838),
.B(n_807),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_820),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_807),
.B(n_829),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_818),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_883),
.B(n_797),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_872),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_855),
.B(n_807),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_883),
.B(n_787),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_868),
.B(n_857),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_805),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_863),
.B(n_884),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_855),
.B(n_856),
.Y(n_892)
);

BUFx8_ASAP7_75t_L g893 ( 
.A(n_851),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_SL g894 ( 
.A1(n_874),
.A2(n_870),
.B1(n_864),
.B2(n_850),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_SL g895 ( 
.A1(n_870),
.A2(n_789),
.B1(n_783),
.B2(n_776),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_856),
.B(n_818),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_863),
.B(n_829),
.Y(n_897)
);

NOR2x1_ASAP7_75t_R g898 ( 
.A(n_851),
.B(n_782),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_879),
.B(n_808),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_873),
.B(n_800),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_849),
.A2(n_876),
.B1(n_854),
.B2(n_872),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_863),
.B(n_802),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_871),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_881),
.B(n_798),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_852),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_901),
.B(n_853),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_905),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_889),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_905),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_889),
.B(n_863),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_896),
.B(n_881),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_891),
.B(n_873),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_901),
.B(n_853),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_891),
.B(n_873),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_892),
.B(n_873),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_887),
.B(n_880),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_887),
.B(n_880),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_891),
.B(n_867),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_893),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_900),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_890),
.B(n_878),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_866),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_911),
.B(n_888),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_919),
.B(n_898),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_921),
.B(n_885),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_918),
.B(n_912),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_907),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_907),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_916),
.B(n_885),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_908),
.B(n_897),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_916),
.B(n_899),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_922),
.B(n_910),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_917),
.B(n_904),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_909),
.B(n_886),
.Y(n_934)
);

OR2x2_ASAP7_75t_SL g935 ( 
.A(n_915),
.B(n_902),
.Y(n_935)
);

AND2x4_ASAP7_75t_SL g936 ( 
.A(n_912),
.B(n_900),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_926),
.B(n_912),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_932),
.B(n_922),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_923),
.B(n_903),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_930),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_924),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_926),
.B(n_912),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_923),
.B(n_903),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_925),
.B(n_914),
.Y(n_944)
);

INVxp33_ASAP7_75t_L g945 ( 
.A(n_934),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_932),
.B(n_910),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_930),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_946),
.B(n_931),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_937),
.B(n_926),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_944),
.B(n_929),
.Y(n_950)
);

INVxp33_ASAP7_75t_L g951 ( 
.A(n_945),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_SL g952 ( 
.A1(n_945),
.A2(n_927),
.B(n_913),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_940),
.B(n_933),
.Y(n_953)
);

NAND4xp25_ASAP7_75t_L g954 ( 
.A(n_941),
.B(n_906),
.C(n_913),
.D(n_895),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_938),
.Y(n_955)
);

NOR4xp25_ASAP7_75t_L g956 ( 
.A(n_939),
.B(n_882),
.C(n_847),
.D(n_848),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_946),
.A2(n_906),
.B(n_900),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_SL g958 ( 
.A1(n_957),
.A2(n_898),
.B(n_861),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_947),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_956),
.A2(n_954),
.B(n_957),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_949),
.B(n_820),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_953),
.Y(n_962)
);

AOI222xp33_ASAP7_75t_L g963 ( 
.A1(n_952),
.A2(n_943),
.B1(n_928),
.B2(n_882),
.C1(n_860),
.C2(n_869),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_961),
.A2(n_951),
.B(n_895),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_SL g965 ( 
.A1(n_960),
.A2(n_861),
.B(n_894),
.Y(n_965)
);

AOI221xp5_ASAP7_75t_SL g966 ( 
.A1(n_962),
.A2(n_935),
.B1(n_953),
.B2(n_928),
.C(n_944),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_965),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_964),
.B(n_846),
.C(n_875),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_967),
.B(n_966),
.Y(n_969)
);

NOR2x1_ASAP7_75t_L g970 ( 
.A(n_968),
.B(n_958),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_970),
.B(n_875),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_969),
.A2(n_836),
.B(n_963),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_971),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_972),
.A2(n_959),
.B(n_859),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_973),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_974),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_974),
.Y(n_977)
);

OAI22x1_ASAP7_75t_L g978 ( 
.A1(n_975),
.A2(n_859),
.B1(n_865),
.B2(n_845),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_976),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_977),
.B(n_949),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_975),
.B(n_893),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_977),
.B(n_865),
.Y(n_982)
);

INVxp33_ASAP7_75t_SL g983 ( 
.A(n_978),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_980),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_981),
.A2(n_845),
.B1(n_894),
.B2(n_948),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_979),
.B(n_982),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_938),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_978),
.A2(n_799),
.B(n_862),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_981),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_989),
.A2(n_877),
.B1(n_858),
.B2(n_935),
.Y(n_990)
);

NAND3x2_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_893),
.C(n_920),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_983),
.A2(n_927),
.B1(n_934),
.B2(n_937),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_SL g993 ( 
.A1(n_986),
.A2(n_893),
.B(n_936),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_SL g994 ( 
.A1(n_990),
.A2(n_987),
.B1(n_985),
.B2(n_988),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_991),
.A2(n_950),
.B(n_942),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_994),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_996),
.B(n_993),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_997),
.A2(n_992),
.B1(n_995),
.B2(n_942),
.Y(n_998)
);


endmodule