module fake_jpeg_30712_n_502 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_54),
.Y(n_158)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_19),
.B(n_8),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_19),
.B(n_8),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_9),
.CON(n_61),
.SN(n_61)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_69),
.Y(n_117)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_24),
.B(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_77),
.B(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_7),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_83),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_97),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_91),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_99),
.Y(n_133)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_10),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

BUFx16f_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_108),
.B(n_91),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_28),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_33),
.B1(n_37),
.B2(n_54),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_113),
.A2(n_115),
.B1(n_130),
.B2(n_139),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_43),
.B1(n_41),
.B2(n_29),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_160),
.B1(n_30),
.B2(n_31),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_33),
.B1(n_37),
.B2(n_18),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_33),
.B1(n_41),
.B2(n_43),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_147),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_37),
.B1(n_18),
.B2(n_49),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_32),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_32),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_29),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_52),
.A2(n_30),
.B1(n_27),
.B2(n_38),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_155),
.B1(n_67),
.B2(n_65),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_81),
.A2(n_18),
.B1(n_44),
.B2(n_38),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_63),
.A2(n_28),
.B1(n_44),
.B2(n_25),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_162),
.B(n_173),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_63),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_163),
.B(n_164),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_110),
.A2(n_53),
.B1(n_55),
.B2(n_51),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_165),
.A2(n_182),
.B1(n_184),
.B2(n_188),
.Y(n_225)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_172),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_47),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_193),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_102),
.B1(n_96),
.B2(n_66),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_185),
.B1(n_206),
.B2(n_208),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_104),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_88),
.B1(n_86),
.B2(n_71),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_73),
.B1(n_22),
.B2(n_72),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_95),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_70),
.B1(n_79),
.B2(n_89),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_116),
.B(n_68),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_189),
.B(n_215),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_104),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_192),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_119),
.B(n_18),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_111),
.B(n_124),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_91),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_200),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_195),
.Y(n_260)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_107),
.B(n_60),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_151),
.A2(n_99),
.B1(n_47),
.B2(n_85),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_144),
.B1(n_173),
.B2(n_125),
.Y(n_234)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_106),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_203),
.A2(n_205),
.B1(n_108),
.B2(n_158),
.Y(n_219)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_124),
.A2(n_79),
.B1(n_94),
.B2(n_2),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_117),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_10),
.B1(n_16),
.B2(n_3),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_123),
.A2(n_6),
.B1(n_15),
.B2(n_3),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_161),
.B1(n_157),
.B2(n_142),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_0),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_122),
.Y(n_254)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_213),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_146),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_132),
.B(n_6),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_142),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_145),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_234),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_146),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_249),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_163),
.A2(n_141),
.B1(n_123),
.B2(n_154),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_232),
.A2(n_236),
.B1(n_245),
.B2(n_257),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_173),
.A2(n_144),
.B(n_143),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_216),
.C(n_195),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_168),
.A2(n_161),
.B1(n_157),
.B2(n_140),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_247),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_177),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g248 ( 
.A1(n_176),
.A2(n_109),
.A3(n_103),
.B1(n_112),
.B2(n_143),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_195),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_193),
.B(n_151),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_112),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_210),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_197),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_178),
.A2(n_103),
.B1(n_122),
.B2(n_138),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_194),
.A2(n_145),
.B(n_11),
.C(n_4),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_172),
.B(n_11),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_167),
.B(n_210),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_238),
.B(n_258),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_205),
.B1(n_191),
.B2(n_213),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_263),
.A2(n_278),
.B(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_272),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_167),
.B1(n_200),
.B2(n_201),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_266),
.A2(n_269),
.B1(n_284),
.B2(n_295),
.Y(n_308)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_182),
.A3(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_267)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_175),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_268),
.B(n_292),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_188),
.B1(n_187),
.B2(n_171),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_206),
.B1(n_214),
.B2(n_183),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_271),
.A2(n_282),
.B1(n_237),
.B2(n_253),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_204),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_273),
.B(n_288),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_220),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_202),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_289),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_235),
.B1(n_253),
.B2(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_203),
.B1(n_211),
.B2(n_198),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_283),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_224),
.A2(n_180),
.B1(n_169),
.B2(n_207),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_227),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_286),
.Y(n_319)
);

INVx3_ASAP7_75t_SL g287 ( 
.A(n_243),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_287),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_166),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_224),
.A2(n_172),
.B1(n_174),
.B2(n_196),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_250),
.A2(n_138),
.B1(n_212),
.B2(n_195),
.Y(n_295)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_234),
.A2(n_0),
.B1(n_1),
.B2(n_170),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_298),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_297),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_170),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_244),
.B1(n_236),
.B2(n_234),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_304),
.B1(n_306),
.B2(n_331),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_233),
.C(n_254),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_311),
.C(n_312),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_292),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_270),
.A2(n_234),
.B1(n_231),
.B2(n_248),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_226),
.C(n_232),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_238),
.C(n_257),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_231),
.B1(n_245),
.B2(n_223),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_316),
.A2(n_271),
.B1(n_274),
.B2(n_282),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_230),
.C(n_222),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_333),
.C(n_274),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_294),
.B(n_274),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_261),
.B(n_222),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_332),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_285),
.A2(n_251),
.B(n_241),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_274),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_270),
.A2(n_259),
.B1(n_230),
.B2(n_243),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_261),
.B(n_251),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_218),
.C(n_240),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_323),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_335),
.Y(n_373)
);

BUFx2_ASAP7_75t_SL g336 ( 
.A(n_328),
.Y(n_336)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_319),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_337),
.Y(n_382)
);

NAND2x1_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_278),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_338),
.A2(n_263),
.B(n_309),
.Y(n_391)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_346),
.Y(n_390)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_349),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_268),
.Y(n_345)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_314),
.B(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_354),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_277),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_350),
.C(n_362),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_272),
.C(n_264),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_351),
.B(n_312),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_314),
.B(n_326),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_353),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_298),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_356),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_283),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_305),
.B1(n_304),
.B2(n_331),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_266),
.B1(n_265),
.B2(n_267),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

CKINVDCx12_ASAP7_75t_R g360 ( 
.A(n_318),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_324),
.B(n_332),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_295),
.C(n_284),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_237),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_252),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_367),
.A2(n_381),
.B1(n_340),
.B2(n_308),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_317),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_371),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_349),
.C(n_348),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_378),
.C(n_383),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_350),
.B(n_302),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_385),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_315),
.B(n_324),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_376),
.A2(n_352),
.B(n_303),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_393),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_317),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_305),
.B1(n_313),
.B2(n_300),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_302),
.C(n_333),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_296),
.B(n_343),
.C(n_341),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_312),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_333),
.C(n_322),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_388),
.B(n_389),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_322),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_391),
.A2(n_290),
.B(n_296),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_321),
.C(n_300),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_321),
.C(n_315),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_346),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_361),
.Y(n_395)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_400),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_398),
.A2(n_399),
.B1(n_403),
.B2(n_415),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_373),
.A2(n_340),
.B1(n_335),
.B2(n_316),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_401),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_410),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_367),
.A2(n_308),
.B1(n_338),
.B2(n_352),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_392),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_404),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_374),
.A2(n_338),
.B1(n_337),
.B2(n_359),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_405),
.A2(n_418),
.B1(n_293),
.B2(n_252),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_407),
.A2(n_408),
.B(n_412),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_365),
.B(n_363),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_355),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_413),
.A2(n_387),
.B(n_388),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_414),
.A2(n_296),
.B(n_279),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_381),
.B1(n_394),
.B2(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

BUFx12_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_378),
.A2(n_347),
.B1(n_329),
.B2(n_330),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_330),
.Y(n_419)
);

OAI322xp33_ASAP7_75t_L g434 ( 
.A1(n_419),
.A2(n_366),
.A3(n_280),
.B1(n_276),
.B2(n_281),
.C1(n_299),
.C2(n_287),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_370),
.C(n_369),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_424),
.C(n_426),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_368),
.C(n_372),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_368),
.C(n_366),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_393),
.B1(n_383),
.B2(n_391),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_437),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_395),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_399),
.A2(n_385),
.B1(n_387),
.B2(n_371),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_431),
.A2(n_406),
.B1(n_397),
.B2(n_408),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_436),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_435),
.C(n_396),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_299),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_287),
.B1(n_259),
.B2(n_243),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_260),
.C(n_240),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_409),
.C(n_418),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_429),
.B1(n_439),
.B2(n_425),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_441),
.A2(n_428),
.B1(n_423),
.B2(n_435),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_404),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_446),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_445),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_421),
.B(n_401),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_449),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_SL g450 ( 
.A(n_420),
.B(n_412),
.C(n_414),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_452),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_419),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_454),
.Y(n_467)
);

HAxp5_ASAP7_75t_SL g452 ( 
.A(n_430),
.B(n_407),
.CON(n_452),
.SN(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_410),
.C(n_403),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_438),
.C(n_431),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_416),
.Y(n_454)
);

OAI21xp33_ASAP7_75t_L g455 ( 
.A1(n_425),
.A2(n_400),
.B(n_398),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_434),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_450),
.A2(n_420),
.B1(n_437),
.B2(n_422),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_457),
.A2(n_466),
.B1(n_423),
.B2(n_170),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_453),
.B(n_444),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_460),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_432),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_465),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_426),
.C(n_427),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_460),
.C(n_458),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_448),
.A2(n_428),
.B1(n_436),
.B2(n_433),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_448),
.A2(n_423),
.B1(n_291),
.B2(n_218),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_468),
.A2(n_423),
.B1(n_11),
.B2(n_4),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_SL g470 ( 
.A1(n_456),
.A2(n_452),
.B(n_451),
.C(n_447),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_469),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_456),
.A2(n_442),
.B(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_475),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_477),
.B(n_479),
.Y(n_484)
);

NOR5xp2_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_170),
.C(n_6),
.D(n_4),
.E(n_5),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_481),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_5),
.B(n_12),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_5),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_482),
.A2(n_470),
.B(n_480),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_467),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_485),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_471),
.B(n_457),
.Y(n_485)
);

OAI321xp33_ASAP7_75t_L g490 ( 
.A1(n_486),
.A2(n_470),
.A3(n_476),
.B1(n_480),
.B2(n_14),
.C(n_17),
.Y(n_490)
);

OAI21x1_ASAP7_75t_SL g497 ( 
.A1(n_490),
.A2(n_492),
.B(n_493),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_491),
.B(n_488),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_487),
.A2(n_470),
.B(n_12),
.C(n_14),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_484),
.Y(n_495)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_495),
.Y(n_499)
);

AOI321xp33_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_489),
.A3(n_14),
.B1(n_17),
.B2(n_1),
.C(n_0),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_498),
.B(n_17),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_497),
.C(n_499),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_0),
.Y(n_502)
);


endmodule