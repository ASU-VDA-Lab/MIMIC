module fake_netlist_1_12391_n_609 (n_117, n_44, n_133, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_16, n_13, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_122, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_132, n_51, n_96, n_39, n_609);
input n_117;
input n_44;
input n_133;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_122;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_51;
input n_96;
input n_39;
output n_609;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_19), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_58), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_2), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_73), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_22), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_53), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_110), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_57), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_52), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_76), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_68), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_44), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_88), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_96), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_51), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_29), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_75), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_54), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_13), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_50), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
INVx1_ASAP7_75t_SL g159 ( .A(n_131), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_84), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_43), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_124), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_10), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_122), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_69), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_78), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_85), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_101), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_11), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_10), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_11), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_82), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_103), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_104), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_28), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_70), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_91), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_24), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_31), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_21), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_128), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_115), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_126), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_120), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_17), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g187 ( .A(n_87), .B(n_40), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_86), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_65), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_63), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_127), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_92), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_46), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_121), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_72), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_98), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g197 ( .A(n_93), .B(n_108), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_14), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_105), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_59), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_35), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_55), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_118), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_99), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_117), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_125), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_153), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_170), .B(n_205), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_175), .B(n_0), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_140), .B(n_1), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_148), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_145), .B(n_3), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_137), .Y(n_215) );
AOI22x1_ASAP7_75t_SL g216 ( .A1(n_163), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_136), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_199), .B(n_6), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_138), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_138), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_139), .B(n_7), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
AOI22x1_ASAP7_75t_SL g224 ( .A1(n_172), .A2(n_8), .B1(n_9), .B2(n_12), .Y(n_224) );
INVx5_ASAP7_75t_L g225 ( .A(n_138), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_201), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_168), .Y(n_228) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_146), .A2(n_62), .B(n_130), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_147), .B(n_8), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_212), .Y(n_231) );
CKINVDCx6p67_ASAP7_75t_R g232 ( .A(n_226), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_227), .B(n_158), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_227), .B(n_150), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_212), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_225), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_214), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_215), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_225), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_209), .B(n_135), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_217), .B(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_214), .Y(n_243) );
INVx5_ASAP7_75t_L g244 ( .A(n_225), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_191), .B1(n_206), .B2(n_204), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_234), .B(n_226), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_234), .B(n_215), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_246), .B(n_219), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_238), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_247), .B(n_218), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_233), .B(n_210), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_231), .B(n_210), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_232), .B(n_228), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_235), .B(n_230), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_241), .B(n_230), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_238), .A2(n_208), .B1(n_213), .B2(n_194), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_248), .Y(n_260) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_242), .B(n_213), .Y(n_261) );
AO22x2_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_224), .B1(n_216), .B2(n_185), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g264 ( .A1(n_243), .A2(n_182), .B1(n_184), .B2(n_152), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_242), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_257), .A2(n_229), .B(n_245), .Y(n_266) );
OAI21xp33_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_141), .B(n_142), .Y(n_267) );
AO21x1_ASAP7_75t_L g268 ( .A1(n_265), .A2(n_188), .B(n_156), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_261), .A2(n_202), .B(n_154), .C(n_186), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_263), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_255), .A2(n_229), .B(n_239), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_252), .B(n_143), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_260), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_250), .B(n_149), .Y(n_274) );
AO21x1_ASAP7_75t_L g275 ( .A1(n_258), .A2(n_198), .B(n_166), .Y(n_275) );
AOI33xp33_ASAP7_75t_L g276 ( .A1(n_259), .A2(n_176), .A3(n_200), .B1(n_196), .B2(n_195), .B3(n_192), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_252), .B(n_169), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_254), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_256), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g280 ( .A1(n_251), .A2(n_159), .B(n_197), .C(n_187), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_264), .B(n_155), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_253), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_264), .B(n_157), .Y(n_283) );
OAI21x1_ASAP7_75t_SL g284 ( .A1(n_268), .A2(n_9), .B(n_262), .Y(n_284) );
AO22x2_ASAP7_75t_L g285 ( .A1(n_281), .A2(n_262), .B1(n_15), .B2(n_16), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_277), .A2(n_262), .B1(n_181), .B2(n_180), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_266), .A2(n_160), .B(n_161), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_278), .B(n_162), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_271), .A2(n_179), .B(n_167), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_279), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_270), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_269), .A2(n_183), .B(n_165), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_276), .B(n_164), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_282), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_272), .B(n_173), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_280), .A2(n_179), .B(n_18), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_281), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_283), .B(n_174), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_274), .A2(n_203), .B(n_178), .Y(n_301) );
AOI21xp33_ASAP7_75t_L g302 ( .A1(n_283), .A2(n_207), .B(n_189), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_270), .A2(n_177), .B1(n_190), .B2(n_193), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_267), .A2(n_244), .B(n_221), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g305 ( .A(n_275), .B(n_244), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_279), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_279), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_297), .A2(n_221), .B1(n_220), .B2(n_211), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_298), .Y(n_309) );
OR2x6_ASAP7_75t_L g310 ( .A(n_306), .B(n_220), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_307), .B(n_244), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_289), .A2(n_221), .B(n_220), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_285), .B(n_240), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_290), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_284), .A2(n_20), .B(n_23), .C(n_25), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_307), .B(n_244), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_285), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_296), .A2(n_27), .B(n_30), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_304), .A2(n_32), .B(n_33), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_304), .A2(n_240), .B(n_36), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
INVx5_ASAP7_75t_SL g323 ( .A(n_291), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_287), .A2(n_240), .B(n_37), .Y(n_324) );
AO32x2_ASAP7_75t_L g325 ( .A1(n_286), .A2(n_34), .A3(n_38), .B1(n_39), .B2(n_41), .Y(n_325) );
NAND3xp33_ASAP7_75t_L g326 ( .A(n_302), .B(n_42), .C(n_45), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
OAI21x1_ASAP7_75t_SL g328 ( .A1(n_292), .A2(n_47), .B(n_48), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_305), .A2(n_49), .B(n_56), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_291), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g331 ( .A1(n_293), .A2(n_60), .B1(n_61), .B2(n_64), .C1(n_66), .C2(n_67), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_300), .B(n_288), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_301), .A2(n_71), .B(n_74), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_298), .B(n_77), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_298), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_298), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_290), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_297), .A2(n_79), .B(n_80), .C(n_81), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_297), .A2(n_89), .B1(n_90), .B2(n_94), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_290), .B(n_95), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_290), .B(n_97), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_SL g347 ( .A1(n_297), .A2(n_102), .B(n_106), .C(n_107), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_298), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_298), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_289), .A2(n_109), .B(n_111), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_337), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_348), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_348), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_349), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_349), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_350), .B(n_112), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_350), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_338), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_309), .B(n_113), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_314), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
INVx5_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_346), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_322), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_322), .B(n_114), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_310), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_314), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_335), .Y(n_376) );
AO21x2_ASAP7_75t_L g377 ( .A1(n_318), .A2(n_116), .B(n_119), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_312), .A2(n_123), .B(n_132), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_314), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_332), .B(n_344), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_345), .B(n_341), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_311), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_336), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_317), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_330), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_334), .B(n_327), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_330), .B(n_325), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_325), .B(n_331), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_328), .A2(n_333), .B1(n_326), .B2(n_343), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_321), .Y(n_391) );
AOI21xp33_ASAP7_75t_SL g392 ( .A1(n_316), .A2(n_333), .B(n_329), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_320), .A2(n_319), .B(n_351), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_325), .Y(n_394) );
BUFx4f_ASAP7_75t_SL g395 ( .A(n_308), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_347), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_342), .B(n_324), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_337), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_332), .B(n_259), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_337), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_322), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_337), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_322), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_337), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_337), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_332), .B(n_259), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_337), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_337), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_309), .B(n_252), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_322), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_337), .B(n_348), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_337), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_374), .B(n_376), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_411), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_380), .B(n_413), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_401), .B(n_412), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_362), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_413), .B(n_382), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_401), .B(n_412), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_363), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_402), .B(n_404), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_399), .B(n_407), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_361), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_414), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_368), .B(n_370), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_352), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_410), .B(n_353), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_399), .B(n_407), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_409), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_355), .B(n_408), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_356), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_387), .B(n_406), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_371), .B(n_403), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_357), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_383), .Y(n_442) );
NAND2x1_ASAP7_75t_L g443 ( .A(n_373), .B(n_359), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_358), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_360), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_381), .B(n_384), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_372), .B(n_385), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_389), .B(n_383), .Y(n_448) );
AND2x4_ASAP7_75t_SL g449 ( .A(n_366), .B(n_373), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_365), .B(n_354), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_369), .Y(n_451) );
INVx5_ASAP7_75t_L g452 ( .A(n_369), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_369), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_388), .B(n_394), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_372), .B(n_359), .Y(n_455) );
AND2x4_ASAP7_75t_SL g456 ( .A(n_366), .B(n_359), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_364), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_379), .B(n_361), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_366), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_367), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_375), .B(n_367), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_367), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_375), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_375), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_395), .B(n_377), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_391), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_377), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_391), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_395), .B(n_396), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_396), .B(n_390), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_392), .B(n_397), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_390), .B(n_393), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_393), .B(n_378), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_369), .Y(n_475) );
INVx5_ASAP7_75t_L g476 ( .A(n_452), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_454), .B(n_417), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_425), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_442), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_418), .Y(n_481) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_424), .B(n_451), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_421), .B(n_437), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_454), .B(n_422), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_433), .B(n_427), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_452), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_422), .B(n_419), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_419), .B(n_473), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_475), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_418), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_429), .B(n_444), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_426), .B(n_423), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_452), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_429), .B(n_440), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_432), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_436), .B(n_444), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_436), .B(n_438), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_435), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_440), .B(n_472), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_472), .B(n_458), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_423), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_430), .B(n_416), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_469), .B(n_447), .Y(n_507) );
AND2x4_ASAP7_75t_SL g508 ( .A(n_455), .B(n_462), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_452), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_467), .B(n_474), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_420), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_445), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_448), .A2(n_471), .B1(n_470), .B2(n_457), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_479), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_498), .B(n_439), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_506), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_477), .B(n_428), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_492), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_501), .B(n_415), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_510), .B(n_456), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_493), .B(n_497), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_493), .B(n_466), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_495), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_477), .B(n_459), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_484), .B(n_464), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_507), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_484), .B(n_443), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_494), .B(n_446), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_488), .B(n_463), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_483), .B(n_465), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_480), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_507), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_481), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_488), .B(n_463), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_505), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_510), .B(n_456), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_503), .B(n_471), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_512), .B(n_461), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_504), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_491), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_512), .B(n_465), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_497), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_504), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_499), .B(n_468), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_499), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_508), .B(n_449), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_534), .B(n_513), .C(n_511), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_526), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_543), .B(n_502), .Y(n_551) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_547), .B(n_487), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_546), .B(n_502), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_531), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_515), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_518), .A2(n_486), .B1(n_487), .B2(n_476), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_525), .B(n_489), .Y(n_557) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_540), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_542), .B(n_489), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_519), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_527), .B(n_500), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_521), .B(n_503), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_524), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_530), .B(n_508), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_532), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_564), .B(n_541), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_552), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_549), .Y(n_570) );
XOR2x2_ASAP7_75t_L g571 ( .A(n_567), .B(n_536), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_555), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_551), .B(n_522), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_567), .A2(n_528), .B1(n_521), .B2(n_537), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_560), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g576 ( .A1(n_556), .A2(n_537), .B(n_538), .Y(n_576) );
OAI32xp33_ASAP7_75t_L g577 ( .A1(n_556), .A2(n_487), .A3(n_496), .B1(n_529), .B2(n_533), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_548), .A2(n_496), .B(n_424), .C(n_451), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_551), .B(n_522), .Y(n_579) );
AOI322xp5_ASAP7_75t_L g580 ( .A1(n_569), .A2(n_485), .A3(n_553), .B1(n_554), .B2(n_550), .C1(n_562), .C2(n_559), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_576), .A2(n_565), .B(n_553), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g582 ( .A1(n_578), .A2(n_558), .B1(n_516), .B2(n_520), .C(n_563), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_570), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_572), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_575), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_577), .A2(n_460), .B(n_482), .Y(n_586) );
OAI21xp33_ASAP7_75t_SL g587 ( .A1(n_580), .A2(n_571), .B(n_574), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_581), .A2(n_538), .B1(n_568), .B2(n_562), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_582), .B(n_544), .C(n_516), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_586), .A2(n_520), .B(n_460), .C(n_573), .Y(n_590) );
NAND3xp33_ASAP7_75t_SL g591 ( .A(n_590), .B(n_585), .C(n_583), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_589), .B(n_579), .Y(n_592) );
OAI21xp33_ASAP7_75t_L g593 ( .A1(n_587), .A2(n_584), .B(n_561), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_593), .B(n_588), .C(n_475), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_592), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_595), .B(n_591), .C(n_509), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_594), .B(n_449), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_596), .Y(n_598) );
NOR4xp75_ASAP7_75t_L g599 ( .A(n_597), .B(n_509), .C(n_561), .D(n_523), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_598), .B(n_539), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_599), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_600), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_601), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_603), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_604), .A2(n_602), .B(n_476), .C(n_490), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_605), .A2(n_490), .B1(n_476), .B2(n_566), .C(n_523), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_606), .A2(n_476), .B(n_490), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_607), .A2(n_476), .B(n_557), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_608), .A2(n_490), .B1(n_535), .B2(n_545), .Y(n_609) );
endmodule