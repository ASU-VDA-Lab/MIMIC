module fake_netlist_1_10166_n_641 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_641);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_641;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_60), .Y(n_73) );
HB1xp67_ASAP7_75t_L g74 ( .A(n_18), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_63), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_49), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_35), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_0), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_52), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_55), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_62), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_15), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_46), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_8), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_6), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_40), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_69), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_23), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_50), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_28), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_44), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_34), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_37), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_43), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_22), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_16), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_15), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_79), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_76), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_77), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_73), .B(n_1), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_79), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_91), .B(n_1), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_95), .B(n_2), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_75), .B(n_2), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_78), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_102), .B(n_74), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_92), .B(n_3), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_95), .B(n_3), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_78), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_82), .B(n_4), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
AND3x1_ASAP7_75t_L g145 ( .A(n_90), .B(n_4), .C(n_5), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
XOR2xp5_ASAP7_75t_L g148 ( .A(n_116), .B(n_5), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_96), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_113), .B(n_7), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_106), .B(n_9), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_78), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_143), .B(n_101), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g158 ( .A1(n_144), .A2(n_117), .B1(n_84), .B2(n_116), .Y(n_158) );
BUFx4f_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_143), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_143), .A2(n_110), .B1(n_109), .B2(n_108), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_136), .B(n_117), .Y(n_162) );
INVxp33_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_144), .B(n_88), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_144), .B(n_93), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_140), .B(n_78), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_118), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_140), .B(n_84), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_137), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_144), .B(n_86), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_130), .B(n_89), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_130), .B(n_114), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_122), .B(n_111), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_122), .B(n_112), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_123), .B(n_107), .Y(n_183) );
INVxp67_ASAP7_75t_SL g184 ( .A(n_130), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_152), .B(n_105), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_123), .B(n_104), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_124), .B(n_103), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_127), .B(n_100), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_118), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_150), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_127), .B(n_99), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_128), .B(n_96), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_128), .B(n_98), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_149), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_129), .B(n_97), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_129), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_118), .Y(n_207) );
NOR2xp33_ASAP7_75t_SL g208 ( .A(n_133), .B(n_41), .Y(n_208) );
NAND2xp33_ASAP7_75t_SL g209 ( .A(n_133), .B(n_10), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_118), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_138), .B(n_42), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_179), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_188), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_204), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_159), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_184), .B(n_145), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_190), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_178), .A2(n_145), .B1(n_125), .B2(n_134), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_163), .B(n_147), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_183), .B(n_189), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_195), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_183), .B(n_139), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_196), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_186), .B(n_153), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_159), .Y(n_228) );
OAI21xp33_ASAP7_75t_L g229 ( .A1(n_161), .A2(n_160), .B(n_167), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_206), .Y(n_232) );
AO22x1_ASAP7_75t_L g233 ( .A1(n_178), .A2(n_139), .B1(n_138), .B2(n_146), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_183), .B(n_146), .Y(n_234) );
NOR2xp33_ASAP7_75t_R g235 ( .A(n_204), .B(n_147), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_206), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_191), .B(n_153), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_171), .Y(n_238) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_158), .B(n_141), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_191), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_178), .A2(n_141), .B1(n_154), .B2(n_156), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_171), .Y(n_242) );
BUFx12f_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_185), .B(n_156), .Y(n_244) );
OR2x6_ASAP7_75t_SL g245 ( .A(n_177), .B(n_148), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_173), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_186), .B(n_154), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_202), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_203), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_178), .A2(n_156), .B1(n_154), .B2(n_151), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_185), .B(n_148), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_189), .B(n_192), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_191), .B(n_151), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_189), .B(n_151), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_192), .B(n_135), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_175), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_174), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_192), .B(n_10), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_163), .B(n_51), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_166), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_166), .Y(n_265) );
INVx5_ASAP7_75t_L g266 ( .A(n_198), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_178), .A2(n_126), .B1(n_120), .B2(n_142), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_180), .B(n_126), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_157), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_203), .A2(n_126), .B1(n_120), .B2(n_142), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_164), .B(n_132), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_231), .A2(n_162), .B1(n_170), .B2(n_177), .C(n_181), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_218), .A2(n_203), .B1(n_209), .B2(n_157), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_215), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_228), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_239), .A2(n_176), .B1(n_187), .B2(n_205), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_226), .B(n_176), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_250), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_226), .B(n_165), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_261), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_250), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_226), .B(n_201), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_243), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_228), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_243), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_249), .B(n_209), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_213), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_250), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_261), .A2(n_203), .B1(n_208), .B2(n_212), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_261), .A2(n_194), .B1(n_198), .B2(n_182), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_250), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_218), .A2(n_194), .B1(n_198), .B2(n_182), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_213), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_248), .B(n_200), .Y(n_295) );
BUFx12f_ASAP7_75t_L g296 ( .A(n_216), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_248), .B(n_200), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_235), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_215), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_222), .A2(n_120), .B1(n_132), .B2(n_142), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_232), .A2(n_210), .B(n_193), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_223), .Y(n_302) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_262), .A2(n_193), .B(n_12), .Y(n_303) );
OAI22x1_ASAP7_75t_L g304 ( .A1(n_218), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_304) );
NAND3xp33_ASAP7_75t_L g305 ( .A(n_220), .B(n_118), .C(n_119), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_258), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_248), .B(n_11), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_258), .Y(n_308) );
AND2x4_ASAP7_75t_SL g309 ( .A(n_258), .B(n_132), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_228), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_228), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_228), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_254), .B(n_16), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_223), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_282), .A2(n_229), .B1(n_256), .B2(n_221), .Y(n_317) );
OR2x6_ASAP7_75t_L g318 ( .A(n_280), .B(n_233), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
AOI222xp33_ASAP7_75t_L g320 ( .A1(n_272), .A2(n_216), .B1(n_244), .B2(n_245), .C1(n_265), .C2(n_234), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_307), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_298), .A2(n_245), .B1(n_252), .B2(n_241), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_287), .Y(n_323) );
CKINVDCx8_ASAP7_75t_R g324 ( .A(n_298), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_283), .B(n_214), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_277), .A2(n_244), .B1(n_252), .B2(n_265), .C(n_224), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_283), .B(n_214), .Y(n_327) );
NOR3xp33_ASAP7_75t_L g328 ( .A(n_276), .B(n_233), .C(n_237), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_277), .B(n_256), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_279), .B(n_256), .Y(n_331) );
CKINVDCx6p67_ASAP7_75t_R g332 ( .A(n_296), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_296), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_294), .B(n_219), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_295), .Y(n_338) );
NAND2x1_ASAP7_75t_L g339 ( .A(n_315), .B(n_219), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_274), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
AND2x6_ASAP7_75t_L g342 ( .A(n_291), .B(n_258), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_286), .A2(n_247), .B1(n_246), .B2(n_260), .C(n_230), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_320), .A2(n_296), .B1(n_280), .B2(n_273), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_322), .A2(n_304), .B1(n_230), .B2(n_264), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_326), .A2(n_293), .B1(n_290), .B2(n_291), .C(n_251), .Y(n_347) );
OAI211xp5_ASAP7_75t_SL g348 ( .A1(n_333), .A2(n_303), .B(n_271), .C(n_268), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_317), .A2(n_290), .B1(n_305), .B2(n_269), .C(n_264), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_344), .A2(n_340), .A3(n_323), .B(n_330), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_334), .B(n_329), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_334), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_318), .A2(n_299), .B1(n_274), .B2(n_314), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_342), .A2(n_285), .B1(n_283), .B2(n_314), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g356 ( .A1(n_317), .A2(n_305), .B1(n_269), .B2(n_214), .C(n_217), .Y(n_356) );
AND2x4_ASAP7_75t_SL g357 ( .A(n_318), .B(n_315), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_342), .A2(n_217), .B1(n_247), .B2(n_260), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_340), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_337), .B(n_283), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_338), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_342), .A2(n_217), .B1(n_246), .B2(n_285), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_342), .A2(n_285), .B1(n_274), .B2(n_314), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_318), .A2(n_302), .B(n_299), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_342), .A2(n_299), .B1(n_302), .B2(n_227), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_342), .A2(n_336), .B1(n_329), .B2(n_321), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g371 ( .A1(n_345), .A2(n_332), .B1(n_319), .B2(n_325), .Y(n_371) );
BUFx4f_ASAP7_75t_L g372 ( .A(n_357), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_352), .B(n_332), .Y(n_373) );
NOR2xp33_ASAP7_75t_R g374 ( .A(n_350), .B(n_315), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_346), .A2(n_328), .B1(n_343), .B2(n_331), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_352), .B(n_341), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_353), .A2(n_327), .B1(n_325), .B2(n_227), .C1(n_225), .C2(n_302), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g378 ( .A1(n_364), .A2(n_339), .B(n_331), .C(n_257), .Y(n_378) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_362), .A2(n_341), .B(n_255), .C(n_267), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_347), .A2(n_327), .B1(n_325), .B2(n_240), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_360), .A2(n_297), .B1(n_240), .B2(n_225), .C(n_300), .Y(n_381) );
NAND5xp2_ASAP7_75t_SL g382 ( .A(n_370), .B(n_17), .C(n_18), .D(n_19), .E(n_20), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_349), .A2(n_300), .B(n_301), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_361), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_361), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_353), .B(n_327), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_362), .A2(n_275), .B1(n_312), .B2(n_311), .C(n_310), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_284), .B1(n_312), .B2(n_311), .C(n_310), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_367), .A2(n_236), .B(n_232), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_275), .B1(n_312), .B2(n_311), .C(n_310), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_368), .A2(n_275), .B1(n_312), .B2(n_311), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_359), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_359), .B(n_17), .Y(n_394) );
NOR2xp33_ASAP7_75t_SL g395 ( .A(n_354), .B(n_278), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_275), .B1(n_310), .B2(n_284), .C(n_238), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_368), .A2(n_316), .B1(n_308), .B2(n_306), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_354), .A2(n_284), .B1(n_238), .B2(n_242), .C(n_253), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_368), .A2(n_284), .B1(n_308), .B2(n_306), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_316), .B1(n_308), .B2(n_306), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_357), .B(n_266), .Y(n_401) );
OR2x6_ASAP7_75t_L g402 ( .A(n_359), .B(n_281), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_357), .A2(n_263), .B1(n_316), .B2(n_308), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_351), .Y(n_404) );
OA21x2_ASAP7_75t_L g405 ( .A1(n_391), .A2(n_369), .B(n_366), .Y(n_405) );
AOI31xp33_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_355), .A3(n_363), .B(n_358), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_384), .B(n_351), .Y(n_407) );
INVx4_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_365), .B1(n_132), .B2(n_142), .C(n_270), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_404), .B(n_351), .Y(n_410) );
NAND4xp75_ASAP7_75t_L g411 ( .A(n_401), .B(n_365), .C(n_351), .D(n_26), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_393), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_382), .A2(n_365), .B1(n_316), .B2(n_306), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_132), .B1(n_142), .B2(n_118), .C(n_119), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_376), .B(n_351), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_372), .A2(n_289), .B1(n_263), .B2(n_292), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_394), .B(n_132), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_374), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_375), .B(n_210), .C(n_259), .D(n_253), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_377), .B(n_142), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_376), .B(n_142), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_402), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_378), .A2(n_119), .B1(n_121), .B2(n_289), .C(n_242), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_402), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_380), .A2(n_289), .B1(n_263), .B2(n_236), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_397), .A2(n_281), .B(n_292), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_392), .B(n_121), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_387), .B(n_259), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_383), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_399), .B(n_119), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_383), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_400), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_396), .B(n_121), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_390), .B(n_21), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_121), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_379), .A2(n_119), .B(n_121), .Y(n_446) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_393), .Y(n_447) );
AOI211xp5_ASAP7_75t_L g448 ( .A1(n_371), .A2(n_119), .B(n_121), .C(n_263), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_372), .A2(n_289), .B1(n_292), .B2(n_288), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_393), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_384), .B(n_121), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_407), .B(n_119), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_423), .B(n_24), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_448), .B(n_292), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_452), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_419), .B(n_27), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_425), .B(n_168), .C(n_169), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_426), .B(n_30), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_407), .B(n_31), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_451), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_447), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_415), .B(n_36), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_441), .B(n_45), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_415), .B(n_47), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_441), .B(n_48), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_453), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_444), .A2(n_428), .B(n_406), .C(n_409), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_422), .B(n_54), .C(n_56), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_450), .B(n_57), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_415), .B(n_58), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_410), .B(n_59), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_453), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_450), .B(n_64), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_437), .B(n_65), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_410), .B(n_66), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_437), .B(n_67), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_427), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_425), .B(n_70), .C(n_72), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_452), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_433), .A2(n_292), .B(n_288), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_410), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_440), .B(n_309), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_440), .B(n_309), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_309), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_431), .B(n_168), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_424), .B(n_168), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_442), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_418), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_438), .B(n_168), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_417), .Y(n_494) );
OAI211xp5_ASAP7_75t_SL g495 ( .A1(n_413), .A2(n_169), .B(n_197), .C(n_207), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
XOR2xp5_ASAP7_75t_L g497 ( .A(n_444), .B(n_263), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_417), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_427), .B(n_169), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_427), .B(n_169), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_424), .B(n_197), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_429), .B(n_197), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_435), .B(n_278), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_429), .B(n_197), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_405), .B(n_207), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_421), .Y(n_506) );
NOR2xp33_ASAP7_75t_SL g507 ( .A(n_408), .B(n_278), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_405), .B(n_207), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_405), .B(n_207), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_484), .B(n_421), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_491), .B(n_435), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_464), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_454), .B(n_430), .Y(n_515) );
NAND2xp33_ASAP7_75t_L g516 ( .A(n_497), .B(n_411), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_474), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_454), .B(n_443), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_485), .B(n_444), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_494), .B(n_434), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_492), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_457), .B(n_443), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_482), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_457), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_470), .B(n_408), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_470), .B(n_408), .C(n_432), .D(n_439), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_498), .B(n_434), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_469), .B(n_445), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_492), .B(n_445), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_506), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_475), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_480), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_496), .B(n_446), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_481), .B(n_414), .C(n_420), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_496), .B(n_446), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_480), .B(n_446), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_490), .B(n_411), .Y(n_538) );
AOI21x1_ASAP7_75t_L g539 ( .A1(n_456), .A2(n_449), .B(n_436), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_211), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_501), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_474), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_461), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_461), .B(n_416), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_508), .B(n_211), .Y(n_545) );
AND4x1_ASAP7_75t_L g546 ( .A(n_458), .B(n_266), .C(n_278), .D(n_281), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_501), .B(n_211), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_467), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_478), .B(n_465), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_467), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_502), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_478), .B(n_211), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_465), .Y(n_553) );
NOR2xp67_ASAP7_75t_SL g554 ( .A(n_456), .B(n_278), .Y(n_554) );
AOI322xp5_ASAP7_75t_L g555 ( .A1(n_473), .A2(n_266), .A3(n_281), .B1(n_288), .B2(n_292), .C1(n_471), .C2(n_466), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_473), .B(n_281), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_514), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_553), .B(n_489), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_515), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_525), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_512), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_524), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_533), .B(n_504), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_531), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_518), .B(n_489), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_517), .B(n_493), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_515), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_493), .Y(n_569) );
NOR2xp67_ASAP7_75t_L g570 ( .A(n_526), .B(n_459), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_533), .B(n_504), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_516), .A2(n_495), .B(n_497), .C(n_507), .Y(n_572) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_544), .B(n_488), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_539), .B(n_504), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_531), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_532), .B(n_509), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
XOR2x2_ASAP7_75t_L g578 ( .A(n_549), .B(n_455), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_510), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_541), .B(n_500), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_554), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_546), .B(n_488), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_520), .A2(n_468), .B1(n_479), .B2(n_477), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_513), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g586 ( .A(n_527), .B(n_500), .C(n_499), .D(n_472), .Y(n_586) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_516), .A2(n_499), .B(n_505), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_522), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_556), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_556), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_535), .B(n_476), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_542), .B(n_503), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_543), .B(n_505), .Y(n_593) );
AO21x1_ASAP7_75t_L g594 ( .A1(n_539), .A2(n_483), .B(n_509), .Y(n_594) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_544), .B(n_486), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_522), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_551), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_521), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_551), .B(n_486), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_523), .B(n_487), .Y(n_600) );
XNOR2x1_ASAP7_75t_L g601 ( .A(n_519), .B(n_487), .Y(n_601) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_538), .A2(n_266), .B(n_288), .C(n_548), .Y(n_602) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_536), .B(n_288), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_528), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_550), .A2(n_529), .B1(n_538), .B2(n_530), .Y(n_605) );
AO22x2_ASAP7_75t_L g606 ( .A1(n_530), .A2(n_537), .B1(n_536), .B2(n_523), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_534), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_555), .B(n_537), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_540), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_534), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_585), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_570), .B(n_602), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_605), .A2(n_606), .B1(n_608), .B2(n_586), .C(n_604), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_572), .B(n_574), .Y(n_614) );
XNOR2xp5_ASAP7_75t_L g615 ( .A(n_578), .B(n_601), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_573), .A2(n_605), .B1(n_606), .B2(n_591), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_577), .B(n_579), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_572), .B(n_574), .Y(n_619) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_602), .B(n_594), .C(n_580), .Y(n_620) );
AOI211xp5_ASAP7_75t_L g621 ( .A1(n_573), .A2(n_583), .B(n_587), .C(n_582), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_565), .Y(n_622) );
AOI322xp5_ASAP7_75t_L g623 ( .A1(n_613), .A2(n_568), .A3(n_595), .B1(n_560), .B2(n_598), .C1(n_561), .C2(n_597), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_621), .A2(n_562), .B1(n_558), .B2(n_557), .C(n_563), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_614), .B(n_580), .C(n_582), .Y(n_625) );
NAND4xp75_ASAP7_75t_L g626 ( .A(n_619), .B(n_567), .C(n_584), .D(n_571), .Y(n_626) );
AOI221x1_ASAP7_75t_SL g627 ( .A1(n_621), .A2(n_592), .B1(n_607), .B2(n_610), .C(n_575), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_615), .A2(n_590), .B1(n_589), .B2(n_566), .C1(n_559), .C2(n_599), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_611), .B(n_599), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_627), .A2(n_616), .B1(n_612), .B2(n_620), .C(n_617), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_624), .A2(n_564), .B1(n_609), .B2(n_622), .Y(n_631) );
NAND3xp33_ASAP7_75t_SL g632 ( .A(n_623), .B(n_618), .C(n_552), .Y(n_632) );
AOI31xp33_ASAP7_75t_L g633 ( .A1(n_628), .A2(n_564), .A3(n_581), .B(n_569), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_633), .A2(n_629), .B1(n_626), .B2(n_625), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_630), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_632), .B1(n_631), .B2(n_596), .Y(n_636) );
OR5x1_ASAP7_75t_L g637 ( .A(n_634), .B(n_603), .C(n_600), .D(n_593), .E(n_576), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_636), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_638), .B(n_637), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_639), .A2(n_588), .B1(n_600), .B2(n_545), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_640), .A2(n_540), .B(n_547), .Y(n_641) );
endmodule