module fake_jpeg_26886_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_0),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_84),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx2_ASAP7_75t_SL g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_53),
.B1(n_60),
.B2(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_72),
.B1(n_57),
.B2(n_62),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_60),
.B1(n_55),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_58),
.B1(n_69),
.B2(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_64),
.B1(n_63),
.B2(n_54),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_47),
.Y(n_106)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_94),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_72),
.B(n_51),
.C(n_56),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_72),
.B1(n_59),
.B2(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_59),
.B1(n_50),
.B2(n_61),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_110),
.B1(n_114),
.B2(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_46),
.C(n_45),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_85),
.A3(n_50),
.B1(n_21),
.B2(n_28),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_92),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_1),
.B(n_2),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_5),
.B(n_6),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_18),
.B1(n_44),
.B2(n_42),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_118),
.Y(n_131)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_126),
.B1(n_112),
.B2(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_9),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_13),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_112),
.B1(n_19),
.B2(n_26),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_17),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_34),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_37),
.C(n_38),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_135),
.C(n_147),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_142),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_144),
.C(n_145),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_139),
.C(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_129),
.Y(n_156)
);


endmodule