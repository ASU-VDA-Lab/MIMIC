module real_jpeg_21179_n_12 (n_5, n_4, n_8, n_0, n_325, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_325;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_0),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_98)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_3),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_3),
.B(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_3),
.B(n_146),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_5),
.A2(n_20),
.B1(n_21),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_5),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_104),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_104),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_57),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_41),
.B(n_45),
.C(n_46),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_8),
.B(n_41),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_8),
.A2(n_10),
.B(n_47),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_20),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_10),
.A2(n_20),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_33),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_61),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_24),
.B(n_63),
.C(n_197),
.Y(n_196)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_11),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_16),
.C(n_281),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_81),
.B(n_321),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_34),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_16),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_29),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_17),
.A2(n_23),
.B(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_18),
.B(n_102),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_27),
.Y(n_18)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_19),
.B(n_31),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_19),
.A2(n_23),
.B(n_31),
.Y(n_282)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_22),
.Y(n_132)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_23),
.B(n_103),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_24),
.A2(n_62),
.B(n_63),
.C(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_24),
.B(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_24),
.B(n_26),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_25),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_29),
.B(n_115),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_32),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_35),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_73),
.C(n_75),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_36),
.A2(n_37),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_54),
.C(n_58),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_38),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_38),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_38),
.A2(n_106),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_38),
.A2(n_58),
.B1(n_59),
.B2(n_106),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_50),
.B(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_39),
.A2(n_97),
.B(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_40),
.B(n_52),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_40),
.B(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_40),
.B(n_98),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_42),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_41),
.A2(n_53),
.B(n_65),
.Y(n_197)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_42),
.A2(n_49),
.B(n_53),
.C(n_161),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_46),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_46),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_46),
.B(n_52),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_48),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_50),
.B(n_53),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_50),
.A2(n_202),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_53),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_54),
.A2(n_55),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_67),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_69),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_62),
.B(n_72),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_62),
.A2(n_67),
.B(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_66),
.B(n_68),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_68),
.A2(n_141),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_69),
.B(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_73),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_73),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_73),
.A2(n_75),
.B1(n_245),
.B2(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_75),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_79),
.B(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_314),
.B(n_320),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_290),
.A3(n_309),
.B1(n_312),
.B2(n_313),
.C(n_325),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_268),
.B(n_289),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_249),
.B(n_267),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_148),
.B(n_231),
.C(n_248),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_134),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_87),
.B(n_134),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_111),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_100),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_89),
.B(n_100),
.C(n_111),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_90),
.B(n_96),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_91),
.A2(n_147),
.B(n_175),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_93),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_94),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_97),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_107),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_105),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_106),
.B(n_294),
.C(n_299),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_109),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_122),
.B1(n_123),
.B2(n_133),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_121),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_113),
.B(n_121),
.C(n_122),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_126),
.B(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_157),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_138),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_140),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_141),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_156),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_230),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_224),
.B(n_229),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_209),
.B(n_223),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_190),
.B(n_208),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_178),
.B(n_189),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_166),
.B(n_177),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_162),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B(n_176),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_180),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_199),
.B1(n_200),
.B2(n_207),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_194),
.A2(n_195),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_194),
.A2(n_195),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_194),
.A2(n_282),
.B(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_195),
.B(n_264),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_202),
.B(n_219),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_218),
.C(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_218),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_246),
.B2(n_247),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_240),
.C(n_247),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_238),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_250),
.B(n_251),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_266),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_262),
.B2(n_263),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_263),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_257),
.C(n_261),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_259),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_270),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_287),
.B2(n_288),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_278),
.B1(n_285),
.B2(n_286),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_273),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_286),
.C(n_288),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B(n_277),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_292),
.C(n_301),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_277),
.B(n_292),
.CI(n_301),
.CON(n_311),
.SN(n_311)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_279),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_280),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_302),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_294),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_304),
.C(n_308),
.Y(n_315)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_310),
.B(n_311),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_317),
.Y(n_319)
);


endmodule