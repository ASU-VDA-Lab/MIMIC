module fake_jpeg_24204_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_10),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_12),
.B(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_23),
.B(n_26),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_33),
.B(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_13),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_28),
.B1(n_18),
.B2(n_10),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_40),
.B1(n_25),
.B2(n_15),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_14),
.B(n_10),
.C(n_25),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_16),
.B(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_39),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_17),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_6),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_51),
.B(n_52),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_54),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_53),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_42),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_44),
.B(n_46),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_9),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_55),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_5),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_69),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_69),
.Y(n_74)
);

OAI31xp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_20),
.A3(n_11),
.B(n_2),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_71),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_20),
.Y(n_79)
);


endmodule