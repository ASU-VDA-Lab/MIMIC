module fake_jpeg_25905_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_30),
.C(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_40),
.Y(n_57)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_2),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_47),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_17),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_66),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_71),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

OA22x2_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_35),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_17),
.B1(n_24),
.B2(n_27),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_15),
.B1(n_20),
.B2(n_45),
.Y(n_101)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_48),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_67),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_61),
.B(n_74),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_102),
.B(n_39),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_70),
.C(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_94),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_79),
.B1(n_20),
.B2(n_15),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_50),
.B(n_46),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_110),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_108),
.C(n_9),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_78),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_16),
.CI(n_22),
.CON(n_126),
.SN(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_80),
.B(n_81),
.C(n_77),
.D(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_80),
.B1(n_79),
.B2(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_113),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_30),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_69),
.B1(n_82),
.B2(n_43),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_89),
.B(n_92),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_93),
.B(n_86),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_120),
.B(n_106),
.Y(n_128)
);

BUFx12f_ASAP7_75t_SL g130 ( 
.A(n_117),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_93),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_120),
.C(n_121),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_133),
.B(n_126),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_123),
.B(n_118),
.C(n_124),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_127),
.B1(n_131),
.B2(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_9),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_7),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_8),
.Y(n_142)
);


endmodule