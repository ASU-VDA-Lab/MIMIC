module real_jpeg_11579_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_41),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_68),
.B1(n_70),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_74),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_4),
.A2(n_41),
.B1(n_45),
.B2(n_74),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_237)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_32),
.B1(n_57),
.B2(n_58),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_32),
.B1(n_41),
.B2(n_45),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_6),
.A2(n_32),
.B1(n_68),
.B2(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_68),
.B1(n_70),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_160),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_7),
.A2(n_41),
.B1(n_45),
.B2(n_160),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_160),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_10),
.A2(n_68),
.B1(n_70),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_131),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_10),
.A2(n_41),
.B1(n_45),
.B2(n_131),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_131),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_11),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_11),
.B(n_76),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_11),
.B(n_30),
.C(n_44),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_11),
.A2(n_41),
.B1(n_45),
.B2(n_151),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_11),
.A2(n_84),
.B1(n_85),
.B2(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_11),
.B(n_107),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_12),
.A2(n_37),
.B1(n_68),
.B2(n_70),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_37),
.B1(n_41),
.B2(n_45),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_12),
.A2(n_37),
.B1(n_57),
.B2(n_58),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_14),
.A2(n_41),
.B1(n_45),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_14),
.A2(n_48),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_148)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_19),
.B(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_78),
.B2(n_79),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_52),
.C(n_64),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_22),
.A2(n_23),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_35),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_26),
.A2(n_85),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_28),
.B(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_30),
.B1(n_42),
.B2(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_29),
.B(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_33),
.A2(n_34),
.B1(n_121),
.B2(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_33),
.A2(n_36),
.B(n_123),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_33),
.A2(n_34),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_35),
.A2(n_84),
.B(n_237),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_38),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_39),
.A2(n_50),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_39),
.A2(n_88),
.B(n_102),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_39),
.A2(n_100),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_39),
.A2(n_49),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_39),
.A2(n_49),
.B1(n_209),
.B2(n_232),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_41),
.A2(n_55),
.B(n_204),
.C(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_41),
.B(n_228),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_45),
.B(n_54),
.C(n_58),
.Y(n_205)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_46),
.A2(n_104),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_47),
.A2(n_49),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_49),
.B(n_151),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_64),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_59),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_53),
.B(n_61),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_53),
.A2(n_154),
.B1(n_155),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_53),
.A2(n_155),
.B1(n_172),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_63)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_56),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_71),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_57),
.B(n_70),
.C(n_71),
.Y(n_152)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_58),
.A2(n_67),
.B(n_150),
.C(n_152),
.Y(n_149)
);

HAxp5_ASAP7_75t_SL g204 ( 
.A(n_58),
.B(n_151),
.CON(n_204),
.SN(n_204)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_62),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_62),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_62),
.A2(n_107),
.B1(n_181),
.B2(n_204),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_75),
.Y(n_64)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_65),
.A2(n_72),
.B1(n_73),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_65),
.A2(n_72),
.B1(n_130),
.B2(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_70),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_76),
.A2(n_93),
.B1(n_150),
.B2(n_159),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_97),
.B2(n_98),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_91),
.B1(n_92),
.B2(n_96),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_87),
.B1(n_96),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_120),
.B(n_122),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_84),
.A2(n_85),
.B1(n_235),
.B2(n_243),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_85),
.B(n_151),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_104),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_105),
.B(n_109),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_105),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_126),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.C(n_128),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_119),
.B(n_124),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_164),
.B(n_277),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_161),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_136),
.B(n_161),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_137),
.B(n_140),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_142),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.C(n_157),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_144),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_157),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_192),
.B(n_272),
.C(n_276),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_185),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.C(n_178),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_167),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_170),
.C(n_174),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_178),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_186),
.B(n_190),
.C(n_191),
.Y(n_273)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_266),
.B(n_271),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_221),
.B(n_265),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_211),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_211),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.C(n_207),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_198),
.A2(n_199),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_207),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_217),
.C(n_219),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_259),
.B(n_264),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_249),
.B(n_258),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_238),
.B(n_248),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_233),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_244),
.B(n_247),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_263)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);


endmodule