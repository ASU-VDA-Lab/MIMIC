module fake_ariane_2975_n_1909 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1909);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1909;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g172 ( 
.A(n_54),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_97),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_83),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_27),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_34),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_14),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_103),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_52),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_0),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_121),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_91),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_60),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_88),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_11),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_60),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_49),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_33),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_22),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_47),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_52),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_49),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_36),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_27),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_82),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_40),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_66),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_36),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_19),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_33),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_118),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_42),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_55),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_35),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_79),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_161),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_75),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_17),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_109),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_44),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_43),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_31),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_104),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_70),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_65),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_28),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_108),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_63),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_26),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_119),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_25),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_41),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_11),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_85),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_18),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_56),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_68),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_77),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_61),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_125),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_71),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_112),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_48),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_25),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_62),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_87),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_73),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_46),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_2),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_154),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_145),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_68),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_67),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_95),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_78),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_81),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_31),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_17),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_40),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_149),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_12),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_67),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_143),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_7),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_2),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_116),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_20),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_93),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_65),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_89),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_167),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_23),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_130),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_74),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_111),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_123),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_3),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_14),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_3),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_66),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_57),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_151),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_34),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_59),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_141),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_53),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_169),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_156),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_139),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_144),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_128),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_43),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_160),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_24),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_86),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_146),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_96),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_155),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_39),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_7),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_152),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_48),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_168),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_15),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_142),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_148),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_50),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_134),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_164),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_6),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_1),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_53),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_41),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_184),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_247),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_247),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_187),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_198),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_257),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_271),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_298),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_316),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_264),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_176),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_294),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_247),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_180),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_294),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_177),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_181),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_180),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_312),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_192),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_177),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_201),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_179),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_172),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_183),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_280),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_192),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_194),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_186),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_194),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_190),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_228),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_321),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_193),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_228),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_232),
.Y(n_384)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_179),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_232),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_195),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_211),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_236),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_196),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_199),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_236),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_209),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_182),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_246),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_211),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_211),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_246),
.B(n_4),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_290),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_212),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_251),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_172),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_251),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_255),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_255),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_203),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_172),
.B(n_4),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_260),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_214),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_260),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_R g411 ( 
.A(n_173),
.B(n_120),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_200),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_261),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_261),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_218),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_267),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_267),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_277),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_221),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_222),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_223),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_233),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_234),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_277),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_295),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_235),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_238),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_295),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_346),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_349),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_352),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_343),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_358),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_374),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_353),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_381),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_355),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_362),
.B(n_274),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_347),
.B(n_388),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_348),
.B(n_175),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_373),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_361),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_359),
.B(n_314),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_377),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_379),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_406),
.A2(n_325),
.B(n_302),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_362),
.B(n_320),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_382),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_R g459 ( 
.A(n_390),
.B(n_174),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_365),
.B(n_302),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_391),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_366),
.B(n_274),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_368),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_421),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_421),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_R g472 ( 
.A(n_393),
.B(n_400),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_375),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_394),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_R g476 ( 
.A(n_360),
.B(n_240),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_409),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_419),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_376),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_378),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_380),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_420),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_384),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_386),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_372),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_R g498 ( 
.A(n_363),
.B(n_242),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_422),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_395),
.A2(n_274),
.B(n_325),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_401),
.B(n_201),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_370),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_484),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_401),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_460),
.B(n_354),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_472),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_503),
.A2(n_326),
.B(n_407),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_423),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_403),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_403),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_435),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_466),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_469),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_453),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_404),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_500),
.B(n_489),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_448),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_466),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_473),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_404),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_484),
.B(n_427),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_405),
.Y(n_534)
);

AO22x2_ASAP7_75t_L g535 ( 
.A1(n_456),
.A2(n_357),
.B1(n_369),
.B2(n_364),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_489),
.B(n_405),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_489),
.B(n_408),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_429),
.B(n_326),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_429),
.B(n_290),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_452),
.B(n_408),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_432),
.B(n_290),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_484),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_432),
.B(n_335),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_466),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_454),
.B(n_396),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_460),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_466),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_442),
.B(n_335),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_482),
.B(n_410),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_364),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_SL g552 ( 
.A(n_457),
.B(n_185),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_482),
.B(n_410),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

BUFx6f_ASAP7_75t_SL g555 ( 
.A(n_505),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_483),
.B(n_413),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_436),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_462),
.A2(n_357),
.B1(n_398),
.B2(n_306),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_485),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_496),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_467),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_485),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_488),
.A2(n_428),
.B1(n_425),
.B2(n_424),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_496),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_462),
.B(n_387),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_486),
.B(n_413),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_496),
.B(n_191),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_467),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_496),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_496),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_496),
.Y(n_577)
);

CKINVDCx11_ASAP7_75t_R g578 ( 
.A(n_439),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_478),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_487),
.B(n_414),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_438),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_490),
.B(n_414),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_490),
.B(n_416),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_492),
.B(n_416),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_442),
.B(n_335),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_492),
.B(n_417),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_493),
.B(n_417),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_438),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_505),
.B(n_369),
.Y(n_591)
);

CKINVDCx11_ASAP7_75t_R g592 ( 
.A(n_444),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_493),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_497),
.B(n_418),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_497),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_480),
.B(n_350),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_430),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_470),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_456),
.B(n_351),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_491),
.B(n_397),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_438),
.B(n_424),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_441),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_502),
.B(n_415),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_445),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_445),
.B(n_425),
.Y(n_608)
);

AO22x2_ASAP7_75t_L g609 ( 
.A1(n_447),
.A2(n_412),
.B1(n_428),
.B2(n_185),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_449),
.B(n_399),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_449),
.B(n_412),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_451),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_451),
.B(n_426),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_488),
.B(n_197),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_488),
.B(n_372),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_447),
.B(n_402),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_494),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_494),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_494),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_459),
.B(n_191),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_499),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_476),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_499),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_499),
.B(n_402),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_504),
.B(n_371),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_471),
.B(n_407),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_431),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_504),
.B(n_201),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_504),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_455),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_455),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_433),
.B(n_385),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_434),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_481),
.B(n_443),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_481),
.B(n_249),
.Y(n_636)
);

INVxp33_ASAP7_75t_SL g637 ( 
.A(n_437),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_481),
.B(n_249),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_440),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_481),
.B(n_249),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_455),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_443),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_474),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_503),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_503),
.Y(n_645)
);

AND2x2_ASAP7_75t_SL g646 ( 
.A(n_474),
.B(n_185),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_443),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_498),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_474),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_441),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_443),
.Y(n_651)
);

BUFx8_ASAP7_75t_SL g652 ( 
.A(n_477),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_443),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_477),
.B(n_197),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_541),
.B(n_443),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_633),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_541),
.B(n_208),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_507),
.B(n_517),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_617),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_507),
.B(n_625),
.Y(n_661)
);

O2A1O1Ixp5_ASAP7_75t_L g662 ( 
.A1(n_533),
.A2(n_213),
.B(n_231),
.C(n_339),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_617),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_591),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_625),
.B(n_465),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_616),
.B(n_611),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_552),
.A2(n_465),
.B1(n_219),
.B2(n_340),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_582),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_517),
.B(n_208),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_200),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_616),
.B(n_611),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_551),
.B(n_202),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_616),
.B(n_465),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_648),
.B(n_243),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_619),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_511),
.B(n_465),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_519),
.B(n_465),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_609),
.A2(n_465),
.B1(n_223),
.B2(n_224),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_551),
.B(n_465),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_591),
.B(n_581),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_619),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_651),
.B(n_210),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_618),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_591),
.B(n_465),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_514),
.B(n_208),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_552),
.A2(n_219),
.B1(n_270),
.B2(n_241),
.Y(n_686)
);

AOI221xp5_ASAP7_75t_L g687 ( 
.A1(n_561),
.A2(n_535),
.B1(n_569),
.B2(n_215),
.C(n_216),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_581),
.B(n_213),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_644),
.B(n_332),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_584),
.B(n_213),
.Y(n_690)
);

INVx8_ASAP7_75t_L g691 ( 
.A(n_539),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_621),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_528),
.A2(n_479),
.B(n_477),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_623),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_622),
.B(n_208),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_629),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_559),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_584),
.B(n_589),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_547),
.B(n_202),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_580),
.B(n_248),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_529),
.B(n_596),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_605),
.B(n_248),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_627),
.B(n_248),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_582),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_SL g705 ( 
.A(n_598),
.B(n_231),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_590),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_613),
.B(n_206),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_645),
.A2(n_479),
.B(n_297),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_512),
.B(n_207),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_512),
.B(n_207),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_613),
.B(n_206),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_590),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_521),
.B(n_239),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_646),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_521),
.B(n_506),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_597),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_525),
.B(n_248),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_597),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_630),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_651),
.B(n_210),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_555),
.A2(n_229),
.B1(n_245),
.B2(n_237),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_642),
.B(n_647),
.Y(n_722)
);

BUFx12f_ASAP7_75t_L g723 ( 
.A(n_578),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_513),
.B(n_239),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_630),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_609),
.A2(n_224),
.B1(n_223),
.B2(n_287),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_516),
.B(n_215),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_577),
.A2(n_479),
.B(n_464),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_607),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_578),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_525),
.B(n_287),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_653),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_518),
.B(n_216),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_520),
.A2(n_252),
.B1(n_342),
.B2(n_341),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_529),
.B(n_217),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_612),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_524),
.B(n_217),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_531),
.B(n_250),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_525),
.B(n_287),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_558),
.B(n_250),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_600),
.B(n_253),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_562),
.B(n_253),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_509),
.B(n_297),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_555),
.A2(n_620),
.B1(n_533),
.B2(n_538),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_646),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_566),
.B(n_259),
.Y(n_746)
);

AND2x6_ASAP7_75t_SL g747 ( 
.A(n_626),
.B(n_259),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_526),
.B(n_244),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_579),
.B(n_263),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_610),
.B(n_254),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_583),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_557),
.B(n_256),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_593),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_595),
.B(n_263),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_602),
.B(n_527),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_620),
.A2(n_204),
.B1(n_338),
.B2(n_337),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_523),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_535),
.A2(n_224),
.B1(n_203),
.B2(n_220),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_532),
.B(n_268),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_523),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_615),
.B(n_268),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_600),
.B(n_258),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_530),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_546),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_538),
.B(n_332),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_624),
.B(n_269),
.Y(n_766)
);

INVx8_ASAP7_75t_L g767 ( 
.A(n_539),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_534),
.B(n_269),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_592),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_626),
.B(n_272),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_526),
.B(n_262),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_530),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_536),
.B(n_272),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_600),
.B(n_281),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_537),
.A2(n_475),
.B(n_464),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_550),
.B(n_281),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_559),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_545),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_522),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_553),
.B(n_286),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_556),
.B(n_286),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_570),
.B(n_288),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_585),
.B(n_288),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_601),
.B(n_266),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_538),
.A2(n_303),
.B1(n_188),
.B2(n_189),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_526),
.B(n_273),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_592),
.Y(n_787)
);

AND2x6_ASAP7_75t_SL g788 ( 
.A(n_626),
.B(n_292),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_586),
.B(n_292),
.Y(n_789)
);

NOR3x1_ASAP7_75t_L g790 ( 
.A(n_599),
.B(n_331),
.C(n_328),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_588),
.B(n_313),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_535),
.A2(n_538),
.B1(n_632),
.B2(n_631),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_545),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_574),
.B(n_275),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_567),
.B(n_313),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_548),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_548),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_594),
.B(n_315),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_563),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_637),
.B(n_278),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_608),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_564),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_315),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_563),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_567),
.B(n_323),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_628),
.B(n_323),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_540),
.A2(n_307),
.B1(n_291),
.B2(n_285),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_574),
.B(n_279),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_538),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_565),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_628),
.B(n_574),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_628),
.B(n_328),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_641),
.A2(n_220),
.B1(n_203),
.B2(n_331),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_539),
.B(n_283),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_565),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_571),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_641),
.A2(n_220),
.B1(n_203),
.B2(n_333),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_571),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_573),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_573),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_539),
.B(n_308),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_643),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_SL g823 ( 
.A(n_730),
.B(n_310),
.C(n_309),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_664),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_661),
.B(n_539),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_730),
.B(n_522),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_691),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_664),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_722),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_729),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_659),
.A2(n_637),
.B1(n_634),
.B2(n_542),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_722),
.B(n_655),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_663),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_729),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_719),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_666),
.B(n_542),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_722),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_764),
.B(n_723),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_691),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_698),
.A2(n_540),
.B1(n_568),
.B2(n_543),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_779),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_SL g842 ( 
.A(n_680),
.B(n_639),
.Y(n_842)
);

AND3x1_ASAP7_75t_SL g843 ( 
.A(n_687),
.B(n_329),
.C(n_336),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_663),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_732),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_675),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_671),
.B(n_542),
.Y(n_847)
);

AO221x1_ASAP7_75t_L g848 ( 
.A1(n_779),
.A2(n_220),
.B1(n_203),
.B2(n_652),
.C(n_543),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_701),
.B(n_560),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_751),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_670),
.B(n_639),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_801),
.B(n_542),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_735),
.B(n_515),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_691),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_675),
.Y(n_855)
);

NOR2x1p5_ASAP7_75t_L g856 ( 
.A(n_723),
.B(n_652),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_795),
.A2(n_549),
.B1(n_587),
.B2(n_544),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_811),
.B(n_653),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_714),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_706),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_811),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_691),
.Y(n_862)
);

NOR2x1p5_ASAP7_75t_L g863 ( 
.A(n_769),
.B(n_575),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_751),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_SL g865 ( 
.A(n_769),
.B(n_304),
.C(n_205),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_706),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_707),
.B(n_542),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_673),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_SL g869 ( 
.A(n_656),
.B(n_540),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_753),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_705),
.A2(n_549),
.B1(n_587),
.B2(n_544),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_787),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_716),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_753),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_767),
.Y(n_875)
);

INVx6_ASAP7_75t_L g876 ( 
.A(n_747),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_736),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_732),
.B(n_509),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_657),
.B(n_672),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_711),
.B(n_544),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_672),
.B(n_544),
.Y(n_881)
);

NOR3xp33_ASAP7_75t_SL g882 ( 
.A(n_787),
.B(n_330),
.C(n_327),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_767),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_712),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_R g885 ( 
.A(n_767),
.B(n_544),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_709),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_809),
.B(n_508),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_712),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_705),
.A2(n_549),
.B1(n_587),
.B2(n_568),
.Y(n_890)
);

NOR2x1p5_ASAP7_75t_L g891 ( 
.A(n_670),
.B(n_575),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_732),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_686),
.A2(n_220),
.B1(n_203),
.B2(n_576),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_R g894 ( 
.A(n_767),
.B(n_549),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_750),
.B(n_674),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_R g896 ( 
.A(n_657),
.B(n_549),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_718),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_715),
.B(n_568),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_795),
.B(n_587),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_735),
.B(n_515),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_806),
.B(n_587),
.Y(n_901)
);

BUFx4f_ASAP7_75t_L g902 ( 
.A(n_770),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_719),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_697),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_757),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_SL g907 ( 
.A(n_800),
.B(n_301),
.C(n_299),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_697),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_725),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_755),
.B(n_564),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_725),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_718),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_714),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_822),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_697),
.Y(n_915)
);

NAND2x2_ASAP7_75t_L g916 ( 
.A(n_741),
.B(n_774),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_777),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_760),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_770),
.Y(n_919)
);

NOR2xp67_ASAP7_75t_L g920 ( 
.A(n_784),
.B(n_572),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_822),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_760),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_770),
.B(n_745),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_658),
.B(n_508),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_809),
.B(n_508),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_763),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_709),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_777),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_777),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_699),
.B(n_636),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_788),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_763),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_778),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_745),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_713),
.B(n_636),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_669),
.B(n_508),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_752),
.B(n_761),
.Y(n_937)
);

INVx5_ASAP7_75t_L g938 ( 
.A(n_802),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_710),
.B(n_635),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_748),
.B(n_509),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_771),
.B(n_509),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_766),
.B(n_638),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_778),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_772),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_772),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_796),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_796),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_762),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_679),
.B(n_684),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_741),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_776),
.B(n_640),
.Y(n_951)
);

CKINVDCx6p67_ASAP7_75t_R g952 ( 
.A(n_786),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_774),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_SL g954 ( 
.A(n_794),
.B(n_226),
.C(n_225),
.Y(n_954)
);

AND2x2_ASAP7_75t_SL g955 ( 
.A(n_765),
.B(n_220),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_780),
.B(n_640),
.Y(n_956)
);

INVx3_ASAP7_75t_SL g957 ( 
.A(n_808),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_793),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_665),
.B(n_510),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_805),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_812),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_781),
.B(n_510),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_793),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_SL g964 ( 
.A(n_734),
.B(n_178),
.C(n_227),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_727),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_799),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_802),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_702),
.B(n_572),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_802),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_799),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_815),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_797),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_815),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_797),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_744),
.A2(n_510),
.B1(n_614),
.B2(n_654),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_765),
.B(n_554),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_807),
.B(n_230),
.C(n_265),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_717),
.B(n_554),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_816),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_782),
.B(n_510),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_816),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_731),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_R g983 ( 
.A(n_814),
.B(n_554),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_700),
.B(n_276),
.C(n_282),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_783),
.B(n_643),
.Y(n_985)
);

AO22x1_ASAP7_75t_L g986 ( 
.A1(n_790),
.A2(n_614),
.B1(n_654),
.B2(n_554),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_660),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_818),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_818),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_739),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_743),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_683),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_695),
.B(n_703),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_685),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_667),
.A2(n_614),
.B1(n_654),
.B2(n_649),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_789),
.B(n_649),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_785),
.A2(n_614),
.B1(n_654),
.B2(n_318),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_688),
.A2(n_319),
.B1(n_289),
.B2(n_293),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_721),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_819),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_SL g1001 ( 
.A(n_733),
.B(n_305),
.C(n_311),
.Y(n_1001)
);

INVx5_ASAP7_75t_L g1002 ( 
.A(n_819),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_791),
.B(n_614),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_820),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_743),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_660),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_690),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_798),
.B(n_604),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_758),
.B(n_604),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_683),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_820),
.Y(n_1011)
);

AOI31xp67_ASAP7_75t_L g1012 ( 
.A1(n_959),
.A2(n_724),
.A3(n_768),
.B(n_773),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_937),
.A2(n_955),
.B1(n_834),
.B2(n_850),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_835),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_854),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_959),
.A2(n_708),
.B(n_682),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_950),
.B(n_726),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_830),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_840),
.A2(n_682),
.B(n_720),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_1003),
.A2(n_682),
.B(n_720),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_965),
.B(n_792),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_935),
.A2(n_720),
.B(n_775),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_829),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_965),
.B(n_960),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_825),
.A2(n_676),
.B(n_677),
.Y(n_1025)
);

AOI31xp67_ASAP7_75t_L g1026 ( 
.A1(n_912),
.A2(n_880),
.A3(n_867),
.B(n_887),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_854),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_1008),
.A2(n_693),
.B(n_662),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_864),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_1009),
.A2(n_728),
.B(n_743),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_910),
.A2(n_689),
.B(n_696),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_868),
.A2(n_704),
.B(n_668),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_829),
.B(n_692),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_912),
.A2(n_694),
.B(n_696),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_950),
.B(n_737),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_869),
.A2(n_689),
.B(n_694),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_837),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1007),
.B(n_738),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_951),
.A2(n_692),
.B(n_803),
.Y(n_1039)
);

AOI211x1_ASAP7_75t_L g1040 ( 
.A1(n_824),
.A2(n_749),
.B(n_742),
.C(n_746),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_870),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_849),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_837),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_955),
.A2(n_759),
.B(n_740),
.C(n_754),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_908),
.B(n_915),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_868),
.A2(n_810),
.B(n_804),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_874),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_877),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_858),
.B(n_681),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_858),
.B(n_681),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_908),
.B(n_821),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_908),
.B(n_678),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_879),
.B(n_756),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_879),
.B(n_828),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_961),
.B(n_813),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_L g1056 ( 
.A1(n_956),
.A2(n_817),
.B(n_650),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_SL g1057 ( 
.A1(n_992),
.A2(n_606),
.B(n_654),
.Y(n_1057)
);

AO22x2_ASAP7_75t_L g1058 ( 
.A1(n_853),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_962),
.A2(n_650),
.B(n_604),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_SL g1060 ( 
.A(n_827),
.B(n_604),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_886),
.B(n_650),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_SL g1062 ( 
.A1(n_839),
.A2(n_655),
.B(n_606),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_980),
.A2(n_650),
.B(n_606),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_869),
.A2(n_334),
.B(n_322),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_L g1065 ( 
.A(n_885),
.B(n_332),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_1010),
.A2(n_5),
.B(n_8),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_886),
.B(n_927),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_927),
.B(n_9),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_859),
.B(n_9),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_953),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_836),
.A2(n_332),
.B(n_464),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_841),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_831),
.A2(n_324),
.B1(n_317),
.B2(n_182),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_898),
.A2(n_852),
.B(n_942),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_847),
.A2(n_332),
.B(n_464),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_948),
.B(n_163),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_985),
.A2(n_332),
.B(n_464),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_919),
.B(n_13),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_859),
.B(n_13),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_898),
.A2(n_475),
.B(n_464),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_851),
.B(n_162),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_996),
.A2(n_332),
.B(n_441),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_903),
.A2(n_475),
.B(n_441),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_884),
.Y(n_1084)
);

CKINVDCx11_ASAP7_75t_R g1085 ( 
.A(n_872),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_975),
.A2(n_332),
.B(n_441),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_SL g1087 ( 
.A1(n_889),
.A2(n_15),
.B(n_16),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_845),
.A2(n_332),
.B(n_441),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_903),
.A2(n_475),
.B(n_317),
.Y(n_1089)
);

AO21x1_ASAP7_75t_L g1090 ( 
.A1(n_893),
.A2(n_925),
.B(n_887),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_845),
.A2(n_475),
.B(n_317),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_977),
.A2(n_317),
.B(n_182),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_913),
.B(n_16),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_905),
.A2(n_20),
.B(n_21),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_920),
.A2(n_317),
.B(n_182),
.C(n_475),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_892),
.A2(n_317),
.B(n_182),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_909),
.A2(n_930),
.B(n_938),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_892),
.A2(n_900),
.B(n_925),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_909),
.A2(n_182),
.B(n_157),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_964),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_999),
.B(n_28),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_906),
.A2(n_30),
.B(n_32),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_861),
.B(n_923),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_835),
.A2(n_153),
.B(n_147),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_911),
.A2(n_135),
.B(n_133),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_938),
.A2(n_132),
.B(n_131),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_908),
.B(n_30),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_832),
.Y(n_1108)
);

AOI211x1_ASAP7_75t_L g1109 ( 
.A1(n_986),
.A2(n_32),
.B(n_35),
.C(n_37),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_911),
.A2(n_126),
.B(n_124),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_860),
.A2(n_115),
.B(n_114),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_833),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_899),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_915),
.B(n_38),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_964),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_866),
.A2(n_106),
.B(n_100),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_923),
.B(n_45),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_826),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_826),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_SL g1120 ( 
.A(n_827),
.B(n_99),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_918),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_873),
.A2(n_94),
.B(n_92),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_902),
.B(n_923),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_938),
.A2(n_84),
.B(n_80),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_888),
.A2(n_76),
.B(n_72),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_897),
.A2(n_947),
.B(n_972),
.Y(n_1126)
);

INVx4_ASAP7_75t_SL g1127 ( 
.A(n_832),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_944),
.A2(n_50),
.B(n_51),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_945),
.A2(n_51),
.B(n_54),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_946),
.A2(n_55),
.B(n_57),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_827),
.B(n_58),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_839),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_922),
.A2(n_58),
.B(n_59),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_861),
.B(n_61),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_913),
.B(n_71),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_938),
.A2(n_63),
.B(n_64),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_934),
.B(n_64),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_926),
.A2(n_69),
.B(n_70),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_974),
.A2(n_1000),
.B(n_921),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_844),
.A2(n_855),
.B(n_846),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_934),
.B(n_891),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_914),
.A2(n_979),
.B(n_973),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_902),
.B(n_876),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_SL g1144 ( 
.A(n_931),
.B(n_838),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_839),
.B(n_862),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_932),
.A2(n_988),
.B(n_943),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_987),
.B(n_1006),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_876),
.B(n_838),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_876),
.B(n_838),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_933),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_915),
.B(n_917),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_SL g1152 ( 
.A1(n_958),
.A2(n_963),
.B(n_981),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_863),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_842),
.B(n_939),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

AO221x2_ASAP7_75t_L g1156 ( 
.A1(n_893),
.A2(n_998),
.B1(n_843),
.B2(n_977),
.C(n_842),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_970),
.A2(n_989),
.B(n_971),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_924),
.A2(n_936),
.B(n_890),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_987),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1006),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_969),
.A2(n_995),
.B(n_878),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_939),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_969),
.A2(n_881),
.B(n_857),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_924),
.A2(n_901),
.A3(n_936),
.B(n_1005),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_857),
.A2(n_904),
.B(n_929),
.Y(n_1165)
);

AOI221x1_ASAP7_75t_L g1166 ( 
.A1(n_1011),
.A2(n_993),
.B1(n_915),
.B2(n_928),
.C(n_967),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_904),
.A2(n_929),
.B(n_827),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_878),
.A2(n_871),
.B(n_997),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_848),
.A2(n_983),
.B(n_1004),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1071),
.A2(n_1004),
.B(n_1002),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1150),
.B(n_939),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1071),
.A2(n_1002),
.B(n_1004),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1075),
.A2(n_1002),
.B(n_1004),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_1077),
.A2(n_1001),
.B(n_954),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1127),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1075),
.A2(n_1002),
.B(n_1005),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1077),
.A2(n_983),
.B(n_1011),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1082),
.A2(n_1011),
.B(n_856),
.Y(n_1178)
);

AO21x1_ASAP7_75t_L g1179 ( 
.A1(n_1013),
.A2(n_998),
.B(n_941),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1108),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1082),
.A2(n_1011),
.B(n_883),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_SL g1182 ( 
.A1(n_1152),
.A2(n_994),
.B(n_928),
.Y(n_1182)
);

OAI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1101),
.A2(n_957),
.B1(n_916),
.B2(n_990),
.C(n_982),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1156),
.A2(n_916),
.B1(n_993),
.B2(n_949),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1100),
.A2(n_957),
.B(n_907),
.C(n_968),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1044),
.A2(n_907),
.B(n_954),
.C(n_984),
.Y(n_1186)
);

OAI221xp5_ASAP7_75t_L g1187 ( 
.A1(n_1101),
.A2(n_823),
.B1(n_984),
.B2(n_882),
.C(n_865),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1070),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1014),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1086),
.A2(n_1001),
.B(n_941),
.Y(n_1190)
);

NAND2x1_ASAP7_75t_L g1191 ( 
.A(n_1015),
.B(n_967),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1014),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1086),
.A2(n_883),
.B(n_917),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1044),
.A2(n_843),
.B(n_940),
.C(n_882),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1042),
.B(n_1035),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1048),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1024),
.B(n_952),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1021),
.B(n_949),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1038),
.B(n_968),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1108),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1072),
.B(n_968),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1036),
.A2(n_1031),
.B(n_1074),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1127),
.B(n_949),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_SL g1204 ( 
.A1(n_1146),
.A2(n_928),
.B(n_917),
.Y(n_1204)
);

BUFx2_ASAP7_75t_SL g1205 ( 
.A(n_1143),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1022),
.A2(n_883),
.B(n_928),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1022),
.A2(n_883),
.B(n_967),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_SL g1208 ( 
.A1(n_1167),
.A2(n_1102),
.B(n_1094),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1059),
.A2(n_967),
.B(n_917),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1059),
.A2(n_1063),
.B(n_1088),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1063),
.A2(n_976),
.B(n_839),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1034),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1156),
.A2(n_832),
.B1(n_978),
.B2(n_896),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1025),
.A2(n_865),
.B(n_823),
.Y(n_1214)
);

CKINVDCx6p67_ASAP7_75t_R g1215 ( 
.A(n_1085),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1067),
.B(n_832),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1039),
.A2(n_896),
.B(n_976),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1156),
.A2(n_832),
.B1(n_991),
.B2(n_885),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1127),
.B(n_862),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1158),
.A2(n_894),
.B(n_875),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1150),
.B(n_875),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1163),
.A2(n_875),
.B(n_1097),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1068),
.A2(n_1040),
.B1(n_1117),
.B2(n_1058),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1088),
.A2(n_1016),
.B(n_1019),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1049),
.B(n_1050),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1123),
.B(n_1108),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1018),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1085),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1080),
.A2(n_1065),
.B(n_1165),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1016),
.A2(n_1019),
.B(n_1030),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1030),
.A2(n_1028),
.B(n_1020),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1119),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1078),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1028),
.A2(n_1020),
.B(n_1091),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1065),
.A2(n_1083),
.B(n_1099),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1029),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1058),
.A2(n_1017),
.B1(n_1049),
.B2(n_1050),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1091),
.A2(n_1096),
.B(n_1168),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1117),
.A2(n_1053),
.B1(n_1144),
.B2(n_1054),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1134),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1045),
.A2(n_1151),
.B(n_1168),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1045),
.A2(n_1151),
.B(n_1161),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1096),
.A2(n_1111),
.B(n_1125),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1134),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1100),
.A2(n_1115),
.B(n_1133),
.C(n_1114),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1058),
.A2(n_1049),
.B1(n_1050),
.B2(n_1117),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1034),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1103),
.B(n_1154),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1090),
.A2(n_1095),
.A3(n_1166),
.B(n_1089),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1033),
.A2(n_1103),
.B1(n_1055),
.B2(n_1112),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1128),
.A2(n_1129),
.B(n_1130),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1041),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1033),
.B(n_1047),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1095),
.A2(n_1052),
.B(n_1051),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1145),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1084),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1111),
.A2(n_1122),
.B(n_1116),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1128),
.A2(n_1130),
.B(n_1129),
.Y(n_1258)
);

NOR2xp67_ASAP7_75t_L g1259 ( 
.A(n_1153),
.B(n_1148),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1116),
.A2(n_1125),
.B(n_1122),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1104),
.A2(n_1110),
.B(n_1105),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1149),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1121),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1033),
.B(n_1103),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1142),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1069),
.A2(n_1093),
.B(n_1135),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1155),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1110),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1161),
.A2(n_1098),
.B(n_1051),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1145),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1023),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1141),
.B(n_1043),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_L g1273 ( 
.A(n_1079),
.B(n_1137),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1157),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1157),
.Y(n_1275)
);

BUFx8_ASAP7_75t_L g1276 ( 
.A(n_1023),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1023),
.B(n_1043),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1098),
.A2(n_1142),
.B(n_1126),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1037),
.B(n_1043),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1037),
.B(n_1159),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1037),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1169),
.A2(n_1057),
.B(n_1126),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1112),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1037),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1139),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1147),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1162),
.B(n_1015),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1160),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1015),
.B(n_1027),
.Y(n_1289)
);

OR2x6_ASAP7_75t_L g1290 ( 
.A(n_1032),
.B(n_1046),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1139),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1132),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1145),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1052),
.A2(n_1092),
.B(n_1140),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1081),
.B(n_1076),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1027),
.B(n_1132),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1169),
.A2(n_1140),
.B(n_1124),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1106),
.A2(n_1138),
.B(n_1073),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1132),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1027),
.B(n_1132),
.Y(n_1300)
);

AO21x1_ASAP7_75t_L g1301 ( 
.A1(n_1107),
.A2(n_1114),
.B(n_1113),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1131),
.A2(n_1107),
.B(n_1136),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1115),
.A2(n_1061),
.B(n_1012),
.Y(n_1303)
);

BUFx2_ASAP7_75t_SL g1304 ( 
.A(n_1145),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1164),
.B(n_1131),
.Y(n_1305)
);

OAI222xp33_ASAP7_75t_L g1306 ( 
.A1(n_1064),
.A2(n_1109),
.B1(n_1066),
.B2(n_1087),
.C1(n_1164),
.C2(n_1026),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1120),
.A2(n_1145),
.B(n_1060),
.C(n_1164),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1062),
.A2(n_1075),
.B(n_1071),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1164),
.A2(n_1075),
.B(n_1071),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1071),
.A2(n_1075),
.B(n_1077),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1077),
.A2(n_1082),
.B(n_1056),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1143),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1101),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1156),
.A2(n_353),
.B1(n_355),
.B2(n_343),
.Y(n_1314)
);

AOI332xp33_ASAP7_75t_L g1315 ( 
.A1(n_1048),
.A2(n_179),
.A3(n_177),
.B1(n_202),
.B2(n_200),
.B3(n_216),
.C1(n_215),
.C2(n_207),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1071),
.A2(n_1075),
.B(n_1077),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1077),
.A2(n_1082),
.B(n_1056),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1108),
.B(n_829),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1101),
.A2(n_561),
.B1(n_541),
.B2(n_452),
.C(n_461),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1101),
.A2(n_546),
.B1(n_601),
.B2(n_701),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1044),
.A2(n_895),
.B(n_661),
.C(n_1013),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1021),
.B(n_853),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1044),
.A2(n_895),
.B(n_661),
.C(n_1013),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1071),
.A2(n_1075),
.B(n_1077),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1042),
.B(n_541),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1127),
.Y(n_1326)
);

BUFx2_ASAP7_75t_R g1327 ( 
.A(n_1118),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1042),
.B(n_541),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1014),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1048),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1108),
.B(n_829),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1255),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1276),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1255),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1189),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1319),
.A2(n_1240),
.B1(n_1320),
.B2(n_1244),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1321),
.A2(n_1323),
.B(n_1185),
.C(n_1194),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1237),
.A2(n_1314),
.B1(n_1313),
.B2(n_1246),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1196),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1223),
.A2(n_1187),
.B1(n_1315),
.B2(n_1266),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1325),
.B(n_1328),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1313),
.A2(n_1239),
.B1(n_1290),
.B2(n_1273),
.Y(n_1342)
);

AOI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1295),
.A2(n_1323),
.B(n_1321),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1313),
.A2(n_1290),
.B1(n_1322),
.B2(n_1179),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1192),
.Y(n_1345)
);

CKINVDCx6p67_ASAP7_75t_R g1346 ( 
.A(n_1215),
.Y(n_1346)
);

AOI221xp5_ASAP7_75t_L g1347 ( 
.A1(n_1245),
.A2(n_1186),
.B1(n_1214),
.B2(n_1194),
.C(n_1183),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1225),
.B(n_1233),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1304),
.B(n_1175),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1199),
.B(n_1216),
.Y(n_1350)
);

AOI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1301),
.A2(n_1186),
.B(n_1208),
.Y(n_1351)
);

AOI22x1_ASAP7_75t_L g1352 ( 
.A1(n_1202),
.A2(n_1289),
.B1(n_1204),
.B2(n_1182),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1195),
.B(n_1286),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1290),
.A2(n_1205),
.B1(n_1201),
.B2(n_1312),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1327),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1225),
.B(n_1264),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1276),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1290),
.A2(n_1322),
.B1(n_1179),
.B2(n_1301),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1171),
.A2(n_1198),
.B1(n_1184),
.B2(n_1330),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1171),
.A2(n_1198),
.B1(n_1250),
.B2(n_1312),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1235),
.A2(n_1229),
.B(n_1245),
.Y(n_1361)
);

INVx8_ASAP7_75t_L g1362 ( 
.A(n_1281),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1262),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1281),
.Y(n_1364)
);

NOR2xp67_ASAP7_75t_SL g1365 ( 
.A(n_1255),
.B(n_1180),
.Y(n_1365)
);

AOI221xp5_ASAP7_75t_L g1366 ( 
.A1(n_1227),
.A2(n_1267),
.B1(n_1236),
.B2(n_1256),
.C(n_1252),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1215),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1232),
.A2(n_1188),
.B1(n_1213),
.B2(n_1197),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1263),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1264),
.B(n_1262),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1283),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1253),
.B(n_1288),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1226),
.B(n_1248),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1307),
.A2(n_1222),
.B(n_1241),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1329),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1228),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1226),
.B(n_1248),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1232),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1270),
.Y(n_1379)
);

INVxp33_ASAP7_75t_L g1380 ( 
.A(n_1259),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1265),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1228),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1226),
.B(n_1248),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1306),
.A2(n_1272),
.B1(n_1280),
.B2(n_1307),
.C(n_1274),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1218),
.A2(n_1203),
.B1(n_1221),
.B2(n_1248),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_R g1386 ( 
.A(n_1270),
.B(n_1293),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1280),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1254),
.A2(n_1203),
.B1(n_1220),
.B2(n_1305),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1289),
.A2(n_1305),
.B1(n_1318),
.B2(n_1331),
.Y(n_1389)
);

AO22x1_ASAP7_75t_L g1390 ( 
.A1(n_1276),
.A2(n_1326),
.B1(n_1175),
.B2(n_1203),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1279),
.Y(n_1391)
);

AND2x6_ASAP7_75t_L g1392 ( 
.A(n_1270),
.B(n_1293),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1289),
.A2(n_1331),
.B1(n_1318),
.B2(n_1293),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1275),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1271),
.B(n_1279),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1175),
.A2(n_1326),
.B1(n_1254),
.B2(n_1174),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1221),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1271),
.B(n_1284),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1287),
.A2(n_1303),
.B1(n_1300),
.B2(n_1296),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1254),
.A2(n_1220),
.B1(n_1326),
.B2(n_1303),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1287),
.A2(n_1219),
.B1(n_1200),
.B2(n_1180),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1303),
.A2(n_1174),
.B1(n_1294),
.B2(n_1190),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1180),
.A2(n_1200),
.B1(n_1284),
.B2(n_1277),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1292),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1219),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1265),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1219),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1294),
.A2(n_1190),
.B1(n_1180),
.B2(n_1200),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1296),
.A2(n_1300),
.B1(n_1191),
.B2(n_1200),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1302),
.A2(n_1298),
.B(n_1209),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1296),
.A2(n_1300),
.B1(n_1292),
.B2(n_1299),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1294),
.A2(n_1190),
.B1(n_1285),
.B2(n_1247),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1292),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_L g1414 ( 
.A(n_1242),
.B(n_1217),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1292),
.B(n_1299),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1212),
.A2(n_1302),
.B1(n_1291),
.B2(n_1258),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1299),
.B(n_1178),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1299),
.B(n_1249),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1178),
.B(n_1249),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1278),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1251),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1211),
.B(n_1269),
.Y(n_1422)
);

NAND2xp33_ASAP7_75t_SL g1423 ( 
.A(n_1291),
.B(n_1317),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1251),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1269),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1251),
.B(n_1258),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1211),
.B(n_1207),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1206),
.B(n_1207),
.Y(n_1428)
);

CKINVDCx14_ASAP7_75t_R g1429 ( 
.A(n_1206),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1258),
.B(n_1209),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1282),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1282),
.B(n_1176),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1238),
.A2(n_1298),
.B(n_1231),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1311),
.B(n_1317),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1311),
.A2(n_1317),
.B1(n_1268),
.B2(n_1257),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1309),
.B(n_1311),
.C(n_1230),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1260),
.A2(n_1243),
.B(n_1297),
.C(n_1238),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1176),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1193),
.A2(n_1297),
.B1(n_1172),
.B2(n_1173),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1170),
.A2(n_1172),
.B1(n_1173),
.B2(n_1309),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1230),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1231),
.A2(n_1234),
.B(n_1316),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1170),
.A2(n_1234),
.B(n_1193),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1224),
.B(n_1210),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1210),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1224),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1181),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1177),
.Y(n_1448)
);

CKINVDCx6p67_ASAP7_75t_R g1449 ( 
.A(n_1177),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1310),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1308),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1324),
.A2(n_1319),
.B1(n_895),
.B2(n_1320),
.C(n_1101),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_SL g1453 ( 
.A(n_1308),
.B(n_580),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1319),
.A2(n_895),
.B(n_1323),
.C(n_1321),
.Y(n_1454)
);

AND2x6_ASAP7_75t_SL g1455 ( 
.A(n_1201),
.B(n_838),
.Y(n_1455)
);

INVx4_ASAP7_75t_L g1456 ( 
.A(n_1281),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1276),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1319),
.A2(n_1240),
.B1(n_895),
.B2(n_1320),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1244),
.B(n_1101),
.Y(n_1459)
);

AOI222xp33_ASAP7_75t_L g1460 ( 
.A1(n_1319),
.A2(n_687),
.B1(n_1101),
.B2(n_1058),
.C1(n_280),
.C2(n_321),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1325),
.B(n_1328),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1264),
.B(n_1225),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_R g1463 ( 
.A(n_1270),
.B(n_1293),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1244),
.B(n_1322),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1262),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1196),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1325),
.B(n_1328),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1452),
.A2(n_1458),
.B1(n_1337),
.B2(n_1454),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1390),
.B(n_1349),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1460),
.A2(n_1338),
.B1(n_1340),
.B2(n_1336),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1355),
.A2(n_1367),
.B1(n_1376),
.B2(n_1382),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1337),
.A2(n_1347),
.B1(n_1342),
.B2(n_1338),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1343),
.A2(n_1358),
.B1(n_1351),
.B2(n_1344),
.C(n_1459),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1363),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1358),
.A2(n_1342),
.B1(n_1344),
.B2(n_1341),
.Y(n_1475)
);

BUFx5_ASAP7_75t_L g1476 ( 
.A(n_1392),
.Y(n_1476)
);

OAI33xp33_ASAP7_75t_L g1477 ( 
.A1(n_1464),
.A2(n_1467),
.A3(n_1461),
.B1(n_1353),
.B2(n_1466),
.B3(n_1369),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1368),
.A2(n_1359),
.B1(n_1350),
.B2(n_1360),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1378),
.A2(n_1359),
.B1(n_1354),
.B2(n_1357),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1362),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1384),
.B(n_1403),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1380),
.A2(n_1366),
.B1(n_1397),
.B2(n_1387),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1362),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1465),
.A2(n_1372),
.B1(n_1371),
.B2(n_1385),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1407),
.A2(n_1383),
.B1(n_1373),
.B2(n_1377),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1429),
.A2(n_1377),
.B1(n_1383),
.B2(n_1407),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1386),
.A2(n_1463),
.B1(n_1457),
.B2(n_1349),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1333),
.A2(n_1361),
.B1(n_1457),
.B2(n_1370),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1457),
.A2(n_1346),
.B1(n_1364),
.B2(n_1456),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1407),
.A2(n_1356),
.B1(n_1400),
.B2(n_1462),
.Y(n_1490)
);

OAI211xp5_ASAP7_75t_L g1491 ( 
.A1(n_1402),
.A2(n_1435),
.B(n_1352),
.C(n_1374),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1462),
.B(n_1395),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1418),
.A2(n_1402),
.B(n_1399),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1400),
.A2(n_1388),
.B1(n_1389),
.B2(n_1375),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1455),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1388),
.A2(n_1405),
.B1(n_1396),
.B2(n_1456),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1362),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1405),
.A2(n_1364),
.B1(n_1392),
.B2(n_1335),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1398),
.B(n_1391),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1413),
.Y(n_1500)
);

BUFx12f_ASAP7_75t_L g1501 ( 
.A(n_1404),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1453),
.A2(n_1447),
.B(n_1439),
.Y(n_1502)
);

OAI211xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1435),
.A2(n_1433),
.B(n_1394),
.C(n_1437),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1386),
.A2(n_1463),
.B1(n_1349),
.B2(n_1401),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1414),
.A2(n_1410),
.B(n_1437),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1404),
.B(n_1379),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1379),
.B(n_1411),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1345),
.A2(n_1393),
.B1(n_1419),
.B2(n_1381),
.Y(n_1508)
);

OAI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1408),
.A2(n_1412),
.B1(n_1434),
.B2(n_1415),
.C(n_1416),
.Y(n_1509)
);

OAI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1408),
.A2(n_1412),
.B1(n_1416),
.B2(n_1423),
.C(n_1409),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1332),
.A2(n_1334),
.B1(n_1403),
.B2(n_1425),
.Y(n_1511)
);

OAI211xp5_ASAP7_75t_L g1512 ( 
.A1(n_1444),
.A2(n_1420),
.B(n_1450),
.C(n_1436),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1381),
.Y(n_1513)
);

O2A1O1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1422),
.A2(n_1450),
.B(n_1334),
.C(n_1332),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1440),
.A2(n_1431),
.B1(n_1432),
.B2(n_1447),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1444),
.B(n_1420),
.C(n_1445),
.Y(n_1516)
);

AOI211xp5_ASAP7_75t_L g1517 ( 
.A1(n_1439),
.A2(n_1417),
.B(n_1422),
.C(n_1426),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1406),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1430),
.A2(n_1440),
.B(n_1421),
.Y(n_1519)
);

OAI211xp5_ASAP7_75t_L g1520 ( 
.A1(n_1424),
.A2(n_1443),
.B(n_1446),
.C(n_1441),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1428),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1365),
.A2(n_1427),
.B(n_1438),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1449),
.A2(n_1448),
.B1(n_1451),
.B2(n_1427),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1451),
.A2(n_1441),
.B1(n_1428),
.B2(n_1442),
.Y(n_1524)
);

AOI222xp33_ASAP7_75t_L g1525 ( 
.A1(n_1451),
.A2(n_1319),
.B1(n_1458),
.B2(n_687),
.C1(n_1058),
.C2(n_1460),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1442),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1442),
.A2(n_1452),
.B1(n_1320),
.B2(n_1458),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1458),
.A2(n_1452),
.B1(n_1336),
.B2(n_1117),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1361),
.A2(n_1454),
.B(n_1323),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_1340),
.B2(n_1058),
.C(n_1452),
.Y(n_1530)
);

OAI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1460),
.A2(n_1319),
.B1(n_895),
.B2(n_1320),
.C(n_1452),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_687),
.B2(n_1058),
.C1(n_1460),
.C2(n_1101),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1348),
.B(n_1356),
.Y(n_1533)
);

NAND4xp25_ASAP7_75t_L g1534 ( 
.A(n_1454),
.B(n_1319),
.C(n_461),
.D(n_1460),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1361),
.A2(n_1454),
.B(n_1323),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1452),
.A2(n_1319),
.B1(n_1458),
.B2(n_1337),
.Y(n_1536)
);

OAI211xp5_ASAP7_75t_L g1537 ( 
.A1(n_1454),
.A2(n_1319),
.B(n_1347),
.C(n_1315),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1460),
.A2(n_1454),
.B(n_1319),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1339),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1340),
.A2(n_1058),
.B1(n_1452),
.B2(n_1458),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1420),
.Y(n_1541)
);

AOI222xp33_ASAP7_75t_L g1542 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_687),
.B2(n_1058),
.C1(n_1460),
.C2(n_1101),
.Y(n_1542)
);

AOI222xp33_ASAP7_75t_L g1543 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_687),
.B2(n_1058),
.C1(n_1460),
.C2(n_1101),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1452),
.A2(n_1319),
.B1(n_1458),
.B2(n_1337),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1460),
.A2(n_1058),
.B1(n_1458),
.B2(n_1319),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1348),
.B(n_1356),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1348),
.B(n_1356),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1420),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1373),
.B(n_1377),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1458),
.A2(n_1452),
.B1(n_1336),
.B2(n_1117),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1452),
.A2(n_1319),
.B1(n_1458),
.B2(n_1337),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1373),
.B(n_1377),
.Y(n_1552)
);

AOI222xp33_ASAP7_75t_L g1553 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_687),
.B2(n_1058),
.C1(n_1460),
.C2(n_1101),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1460),
.A2(n_1058),
.B1(n_1458),
.B2(n_1319),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1373),
.B(n_1377),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1454),
.A2(n_1319),
.B(n_1347),
.C(n_1315),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1452),
.A2(n_1319),
.B1(n_1458),
.B2(n_1337),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1460),
.A2(n_1058),
.B1(n_1458),
.B2(n_1319),
.Y(n_1558)
);

AND2x6_ASAP7_75t_SL g1559 ( 
.A(n_1459),
.B(n_838),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_1340),
.B2(n_1058),
.C(n_1452),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1460),
.A2(n_1058),
.B1(n_1458),
.B2(n_1319),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1460),
.A2(n_1058),
.B1(n_1458),
.B2(n_1319),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1452),
.A2(n_1319),
.B1(n_1458),
.B2(n_1337),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1458),
.A2(n_1319),
.B1(n_1340),
.B2(n_1058),
.C(n_1452),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1460),
.A2(n_1058),
.B1(n_1458),
.B2(n_1319),
.Y(n_1565)
);

AOI21xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1367),
.A2(n_637),
.B(n_1458),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1348),
.B(n_1356),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1348),
.B(n_1356),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1414),
.A2(n_1268),
.B(n_1261),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1362),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1505),
.Y(n_1571)
);

NAND2xp33_ASAP7_75t_SL g1572 ( 
.A(n_1468),
.B(n_1536),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1526),
.B(n_1521),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1521),
.B(n_1517),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1535),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1493),
.B(n_1505),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1548),
.Y(n_1578)
);

OR2x6_ASAP7_75t_SL g1579 ( 
.A(n_1544),
.B(n_1551),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1557),
.B(n_1563),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1548),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1516),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1525),
.A2(n_1554),
.B1(n_1545),
.B2(n_1565),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1545),
.A2(n_1565),
.B1(n_1562),
.B2(n_1561),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1519),
.B(n_1512),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1502),
.A2(n_1491),
.B(n_1508),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1569),
.B(n_1533),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1569),
.B(n_1507),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1513),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1518),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1567),
.B(n_1568),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1539),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1515),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1520),
.Y(n_1595)
);

NOR2xp67_ASAP7_75t_R g1596 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1481),
.B(n_1523),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1476),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1490),
.B(n_1508),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1524),
.B(n_1509),
.Y(n_1600)
);

OAI221xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1538),
.A2(n_1554),
.B1(n_1558),
.B2(n_1561),
.C(n_1562),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1503),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1490),
.B(n_1522),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1524),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1476),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1514),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1511),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1510),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1558),
.A2(n_1532),
.B1(n_1542),
.B2(n_1543),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1527),
.B(n_1475),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_L g1612 ( 
.A(n_1487),
.B(n_1469),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1609),
.A2(n_1553),
.B1(n_1534),
.B2(n_1540),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_R g1614 ( 
.A(n_1572),
.B(n_1483),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1574),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1574),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_R g1617 ( 
.A(n_1580),
.B(n_1495),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1578),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1610),
.A2(n_1479),
.B1(n_1531),
.B2(n_1472),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1576),
.B(n_1482),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1598),
.Y(n_1622)
);

AND2x2_ASAP7_75t_SL g1623 ( 
.A(n_1577),
.B(n_1586),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1609),
.A2(n_1470),
.B1(n_1564),
.B2(n_1560),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1590),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1576),
.A2(n_1550),
.B(n_1528),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_L g1628 ( 
.A(n_1572),
.B(n_1530),
.C(n_1556),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1598),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1580),
.B(n_1471),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1578),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1608),
.A2(n_1470),
.B1(n_1528),
.B2(n_1550),
.C(n_1477),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1590),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1579),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1610),
.A2(n_1478),
.B1(n_1481),
.B2(n_1484),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1578),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1585),
.B(n_1488),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1610),
.A2(n_1478),
.B1(n_1484),
.B2(n_1504),
.Y(n_1639)
);

BUFx4f_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1608),
.A2(n_1537),
.B1(n_1482),
.B2(n_1566),
.C(n_1504),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1591),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1573),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_SL g1644 ( 
.A(n_1585),
.B(n_1496),
.C(n_1474),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1601),
.A2(n_1496),
.B1(n_1498),
.B2(n_1485),
.C(n_1486),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1593),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1579),
.B(n_1489),
.Y(n_1647)
);

OA211x2_ASAP7_75t_L g1648 ( 
.A1(n_1576),
.A2(n_1498),
.B(n_1499),
.C(n_1485),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1585),
.A2(n_1506),
.B(n_1483),
.C(n_1480),
.Y(n_1649)
);

NAND4xp25_ASAP7_75t_L g1650 ( 
.A(n_1583),
.B(n_1570),
.C(n_1480),
.D(n_1492),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_SL g1652 ( 
.A1(n_1610),
.A2(n_1549),
.B1(n_1552),
.B2(n_1559),
.Y(n_1652)
);

INVx5_ASAP7_75t_L g1653 ( 
.A(n_1571),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1579),
.A2(n_1497),
.B1(n_1570),
.B2(n_1611),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1587),
.Y(n_1655)
);

NOR2x1p5_ASAP7_75t_L g1656 ( 
.A(n_1634),
.B(n_1606),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1622),
.B(n_1605),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1623),
.B(n_1588),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1619),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1619),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1618),
.B(n_1594),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1620),
.A2(n_1595),
.B(n_1611),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1615),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1637),
.B(n_1582),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1631),
.B(n_1594),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1582),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1630),
.B(n_1579),
.Y(n_1667)
);

NAND4xp25_ASAP7_75t_L g1668 ( 
.A(n_1628),
.B(n_1583),
.C(n_1601),
.D(n_1584),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1626),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1623),
.B(n_1588),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1622),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1623),
.B(n_1577),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1626),
.B(n_1588),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1622),
.B(n_1605),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1621),
.B(n_1606),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1622),
.B(n_1588),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1642),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1616),
.B(n_1595),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1629),
.B(n_1588),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1633),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1629),
.B(n_1588),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1624),
.B(n_1577),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1636),
.B(n_1577),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1653),
.B(n_1612),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1634),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1646),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1629),
.B(n_1573),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1653),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1653),
.B(n_1571),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1646),
.B(n_1581),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1686),
.B(n_1672),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1676),
.B(n_1634),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1674),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_1589),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1676),
.B(n_1679),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1674),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1659),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1659),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1679),
.B(n_1602),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1667),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1659),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1667),
.B(n_1647),
.Y(n_1704)
);

NAND4xp25_ASAP7_75t_L g1705 ( 
.A(n_1662),
.B(n_1613),
.C(n_1641),
.D(n_1625),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1656),
.B(n_1649),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1661),
.B(n_1589),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1661),
.B(n_1602),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1661),
.B(n_1665),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1665),
.B(n_1602),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1656),
.A2(n_1592),
.B(n_1589),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1663),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1686),
.B(n_1589),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1663),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1664),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1656),
.B(n_1651),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1660),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1665),
.B(n_1638),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1673),
.Y(n_1719)
);

NAND2x1_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1651),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1664),
.B(n_1607),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1686),
.B(n_1592),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1666),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1660),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1672),
.B(n_1614),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1660),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1666),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1672),
.B(n_1607),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1669),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1658),
.B(n_1670),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1698),
.Y(n_1731)
);

NAND2xp33_ASAP7_75t_SL g1732 ( 
.A(n_1720),
.B(n_1662),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1698),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1699),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1730),
.B(n_1658),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1730),
.B(n_1658),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1730),
.B(n_1658),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1699),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1715),
.B(n_1723),
.Y(n_1739)
);

AND2x2_ASAP7_75t_SL g1740 ( 
.A(n_1704),
.B(n_1640),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1706),
.B(n_1670),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1692),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1693),
.B(n_1670),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1705),
.A2(n_1608),
.B1(n_1644),
.B2(n_1611),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1692),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1727),
.B(n_1669),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1700),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1700),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1701),
.B(n_1669),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1693),
.B(n_1670),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1697),
.B(n_1684),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1708),
.B(n_1684),
.Y(n_1752)
);

INVx4_ASAP7_75t_L g1753 ( 
.A(n_1716),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1677),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1703),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1710),
.B(n_1683),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1703),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1718),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1683),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1717),
.Y(n_1760)
);

CKINVDCx16_ASAP7_75t_R g1761 ( 
.A(n_1696),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1717),
.Y(n_1762)
);

OAI31xp33_ASAP7_75t_L g1763 ( 
.A1(n_1702),
.A2(n_1668),
.A3(n_1597),
.B(n_1654),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_L g1764 ( 
.A(n_1725),
.B(n_1689),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1696),
.B(n_1677),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1695),
.B(n_1683),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1713),
.B(n_1677),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1712),
.B(n_1681),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1724),
.Y(n_1769)
);

NOR3xp33_ASAP7_75t_L g1770 ( 
.A(n_1728),
.B(n_1668),
.C(n_1632),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

NAND4xp75_ASAP7_75t_L g1772 ( 
.A(n_1694),
.B(n_1648),
.C(n_1627),
.D(n_1586),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1713),
.B(n_1677),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1770),
.B(n_1722),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1731),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1731),
.Y(n_1776)
);

NOR3xp33_ASAP7_75t_SL g1777 ( 
.A(n_1732),
.B(n_1761),
.C(n_1741),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1743),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1770),
.B(n_1722),
.Y(n_1779)
);

OAI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1763),
.A2(n_1744),
.B1(n_1758),
.B2(n_1635),
.C(n_1772),
.Y(n_1780)
);

AOI32xp33_ASAP7_75t_L g1781 ( 
.A1(n_1758),
.A2(n_1575),
.A3(n_1709),
.B1(n_1639),
.B2(n_1673),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1733),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1761),
.B(n_1716),
.Y(n_1783)
);

XNOR2x2_ASAP7_75t_L g1784 ( 
.A(n_1772),
.B(n_1650),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1733),
.Y(n_1785)
);

NAND3x2_ASAP7_75t_L g1786 ( 
.A(n_1743),
.B(n_1716),
.C(n_1657),
.Y(n_1786)
);

AOI211x1_ASAP7_75t_L g1787 ( 
.A1(n_1743),
.A2(n_1714),
.B(n_1682),
.C(n_1680),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1750),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1734),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1763),
.A2(n_1597),
.B(n_1586),
.Y(n_1790)
);

OAI21xp33_ASAP7_75t_L g1791 ( 
.A1(n_1739),
.A2(n_1719),
.B(n_1707),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1734),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1739),
.B(n_1707),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1673),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1753),
.B(n_1720),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1755),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1755),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1766),
.B(n_1719),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1735),
.B(n_1688),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1740),
.A2(n_1648),
.B1(n_1600),
.B2(n_1650),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1759),
.B(n_1655),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1740),
.A2(n_1597),
.B1(n_1600),
.B2(n_1685),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1764),
.A2(n_1740),
.B(n_1768),
.Y(n_1803)
);

OAI322xp33_ASAP7_75t_L g1804 ( 
.A1(n_1752),
.A2(n_1600),
.A3(n_1617),
.B1(n_1597),
.B2(n_1729),
.C1(n_1726),
.C2(n_1691),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1751),
.B(n_1655),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1735),
.A2(n_1597),
.B1(n_1600),
.B2(n_1685),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1738),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1738),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1747),
.Y(n_1809)
);

OAI31xp33_ASAP7_75t_L g1810 ( 
.A1(n_1780),
.A2(n_1750),
.A3(n_1645),
.B(n_1685),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1777),
.B(n_1735),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1774),
.Y(n_1812)
);

INVxp33_ASAP7_75t_L g1813 ( 
.A(n_1777),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1790),
.A2(n_1779),
.B(n_1803),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_1750),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1804),
.A2(n_1749),
.B1(n_1752),
.B2(n_1762),
.C(n_1771),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1784),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1784),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1808),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1778),
.Y(n_1820)
);

AOI31xp33_ASAP7_75t_L g1821 ( 
.A1(n_1783),
.A2(n_1736),
.A3(n_1737),
.B(n_1754),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1808),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1800),
.A2(n_1584),
.B1(n_1599),
.B2(n_1586),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1807),
.Y(n_1824)
);

OAI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1783),
.A2(n_1766),
.B(n_1754),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1778),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1806),
.A2(n_1599),
.B1(n_1586),
.B2(n_1603),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1793),
.B(n_1751),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1809),
.Y(n_1829)
);

OAI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1781),
.A2(n_1788),
.B(n_1791),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1788),
.Y(n_1831)
);

NAND2x1_ASAP7_75t_L g1832 ( 
.A(n_1795),
.B(n_1753),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1775),
.B(n_1736),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1786),
.A2(n_1736),
.B(n_1737),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1802),
.A2(n_1753),
.B1(n_1685),
.B2(n_1782),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1811),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1812),
.B(n_1776),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1828),
.B(n_1789),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1820),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1817),
.B(n_1753),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_R g1841 ( 
.A(n_1819),
.B(n_1792),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1842)
);

AOI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1813),
.A2(n_1795),
.B(n_1797),
.C(n_1737),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1817),
.B(n_1768),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1818),
.B(n_1787),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1820),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1826),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1826),
.Y(n_1848)
);

NOR3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1814),
.B(n_1805),
.C(n_1801),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1831),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1831),
.Y(n_1851)
);

NOR4xp25_ASAP7_75t_L g1852 ( 
.A(n_1818),
.B(n_1748),
.C(n_1762),
.D(n_1760),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1824),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1824),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1829),
.Y(n_1855)
);

NAND5xp2_ASAP7_75t_L g1856 ( 
.A(n_1843),
.B(n_1813),
.C(n_1811),
.D(n_1834),
.E(n_1830),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1836),
.B(n_1833),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1852),
.A2(n_1810),
.B(n_1822),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_SL g1859 ( 
.A1(n_1840),
.A2(n_1822),
.B(n_1829),
.C(n_1815),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1841),
.B(n_1835),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1845),
.A2(n_1821),
.B(n_1825),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1844),
.A2(n_1816),
.B1(n_1823),
.B2(n_1827),
.C(n_1833),
.Y(n_1862)
);

OAI211xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1849),
.A2(n_1832),
.B(n_1794),
.C(n_1798),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1844),
.B(n_1832),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1840),
.B(n_1849),
.Y(n_1865)
);

AOI211xp5_ASAP7_75t_L g1866 ( 
.A1(n_1837),
.A2(n_1833),
.B(n_1752),
.C(n_1745),
.Y(n_1866)
);

BUFx8_ASAP7_75t_SL g1867 ( 
.A(n_1853),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1858),
.A2(n_1850),
.B1(n_1847),
.B2(n_1846),
.C(n_1839),
.Y(n_1868)
);

AOI32xp33_ASAP7_75t_L g1869 ( 
.A1(n_1863),
.A2(n_1855),
.A3(n_1854),
.B1(n_1851),
.B2(n_1848),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1857),
.Y(n_1870)
);

OAI211xp5_ASAP7_75t_L g1871 ( 
.A1(n_1859),
.A2(n_1842),
.B(n_1838),
.C(n_1754),
.Y(n_1871)
);

O2A1O1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1865),
.A2(n_1749),
.B(n_1748),
.C(n_1757),
.Y(n_1872)
);

O2A1O1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1861),
.A2(n_1769),
.B(n_1760),
.C(n_1757),
.Y(n_1873)
);

OAI211xp5_ASAP7_75t_L g1874 ( 
.A1(n_1864),
.A2(n_1799),
.B(n_1773),
.C(n_1765),
.Y(n_1874)
);

AOI21xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1860),
.A2(n_1689),
.B(n_1747),
.Y(n_1875)
);

AOI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1856),
.A2(n_1742),
.B(n_1745),
.C(n_1756),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1862),
.A2(n_1746),
.B(n_1769),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1866),
.A2(n_1771),
.B1(n_1742),
.B2(n_1745),
.C(n_1746),
.Y(n_1878)
);

XNOR2xp5_ASAP7_75t_L g1879 ( 
.A(n_1870),
.B(n_1867),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1871),
.A2(n_1773),
.B(n_1767),
.Y(n_1880)
);

NAND4xp25_ASAP7_75t_SL g1881 ( 
.A(n_1869),
.B(n_1773),
.C(n_1767),
.D(n_1765),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1872),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1876),
.B(n_1742),
.Y(n_1883)
);

OAI31xp33_ASAP7_75t_L g1884 ( 
.A1(n_1877),
.A2(n_1685),
.A3(n_1756),
.B(n_1767),
.Y(n_1884)
);

NAND4xp75_ASAP7_75t_L g1885 ( 
.A(n_1882),
.B(n_1868),
.C(n_1878),
.D(n_1875),
.Y(n_1885)
);

OAI211xp5_ASAP7_75t_L g1886 ( 
.A1(n_1880),
.A2(n_1873),
.B(n_1874),
.C(n_1765),
.Y(n_1886)
);

AOI221x1_ASAP7_75t_L g1887 ( 
.A1(n_1883),
.A2(n_1879),
.B1(n_1881),
.B2(n_1884),
.C(n_1729),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1879),
.Y(n_1888)
);

NAND3x1_ASAP7_75t_L g1889 ( 
.A(n_1882),
.B(n_1671),
.C(n_1726),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1879),
.Y(n_1890)
);

OAI21xp33_ASAP7_75t_L g1891 ( 
.A1(n_1890),
.A2(n_1682),
.B(n_1680),
.Y(n_1891)
);

OAI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1887),
.A2(n_1671),
.B(n_1689),
.C(n_1682),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1886),
.A2(n_1586),
.B1(n_1575),
.B2(n_1497),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1889),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1886),
.A2(n_1687),
.B1(n_1604),
.B2(n_1571),
.C(n_1575),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1894),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1891),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1892),
.B(n_1888),
.Y(n_1898)
);

NOR2x1_ASAP7_75t_L g1899 ( 
.A(n_1898),
.B(n_1885),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1899),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1900),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1900),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1902),
.B(n_1896),
.Y(n_1903)
);

OAI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1902),
.A2(n_1897),
.B1(n_1895),
.B2(n_1893),
.Y(n_1904)
);

AOI222xp33_ASAP7_75t_L g1905 ( 
.A1(n_1903),
.A2(n_1901),
.B1(n_1640),
.B2(n_1690),
.C1(n_1599),
.C2(n_1678),
.Y(n_1905)
);

NOR2xp67_ASAP7_75t_L g1906 ( 
.A(n_1904),
.B(n_1497),
.Y(n_1906)
);

XNOR2xp5_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1652),
.Y(n_1907)
);

OAI221xp5_ASAP7_75t_R g1908 ( 
.A1(n_1907),
.A2(n_1905),
.B1(n_1596),
.B2(n_1671),
.C(n_1675),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1497),
.B(n_1690),
.C(n_1596),
.Y(n_1909)
);


endmodule