module fake_jpeg_30797_n_70 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_39),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_5),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_47),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_31),
.C(n_27),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_46),
.C(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_48),
.B1(n_9),
.B2(n_10),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_22),
.C(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_6),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_18),
.C(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_20),
.B1(n_15),
.B2(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

XNOR2x1_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_6),
.C(n_7),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_9),
.C(n_11),
.Y(n_58)
);

XOR2x2_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_12),
.Y(n_62)
);

OAI321xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_11),
.A3(n_12),
.B1(n_50),
.B2(n_54),
.C(n_58),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_68),
.B(n_67),
.Y(n_70)
);


endmodule