module real_jpeg_33786_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_290;
wire n_239;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_0),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_0),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_1),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_1),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_1),
.B(n_374),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_1),
.B(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_SL g502 ( 
.A(n_1),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_2),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

NAND2x1_ASAP7_75t_SL g137 ( 
.A(n_2),
.B(n_138),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_2),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_248),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_R g285 ( 
.A(n_2),
.B(n_286),
.Y(n_285)
);

AND2x4_ASAP7_75t_SL g55 ( 
.A(n_3),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_3),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_3),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_3),
.B(n_43),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_84),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_166),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_4),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_6),
.B(n_43),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_6),
.B(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_6),
.A2(n_282),
.B(n_284),
.Y(n_281)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_6),
.Y(n_345)
);

NAND2x1_ASAP7_75t_SL g376 ( 
.A(n_6),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_6),
.B(n_282),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g485 ( 
.A(n_6),
.B(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_6),
.B(n_515),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_8),
.Y(n_344)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_9),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_10),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_10),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_10),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_10),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_10),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_10),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_10),
.B(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_11),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_11),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_11),
.Y(n_464)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_13),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_13),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_13),
.B(n_82),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_13),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_13),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_13),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_13),
.B(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_14),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_15),
.B(n_43),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_15),
.B(n_40),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_15),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_15),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_15),
.B(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_15),
.B(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_15),
.B(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_47),
.Y(n_46)
);

AND2x4_ASAP7_75t_SL g90 ( 
.A(n_17),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_17),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_17),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_17),
.B(n_245),
.Y(n_244)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_167),
.B(n_552),
.C(n_558),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

AOI221xp5_ASAP7_75t_L g558 ( 
.A1(n_20),
.A2(n_21),
.B1(n_554),
.B2(n_557),
.C(n_559),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_153),
.C(n_165),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_130),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_22),
.B(n_130),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.C(n_99),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_23),
.B(n_75),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_49),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_25),
.B(n_64),
.C(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_38),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_32),
.B(n_36),
.C(n_38),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_32),
.A2(n_37),
.B1(n_129),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_32),
.A2(n_37),
.B1(n_207),
.B2(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_35),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_37),
.B(n_123),
.C(n_129),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_37),
.B(n_200),
.C(n_207),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.C(n_45),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_42),
.B(n_120),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_42),
.B(n_158),
.CI(n_159),
.CON(n_157),
.SN(n_157)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_44),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_45),
.B(n_201),
.C(n_205),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_45),
.A2(n_46),
.B1(n_205),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_63),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_51),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_53),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_54)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_61),
.B1(n_65),
.B2(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_57),
.Y(n_380)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_61),
.C(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_62),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_58),
.A2(n_62),
.B1(n_228),
.B2(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_65),
.C(n_70),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_61),
.B(n_109),
.C(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_61),
.B(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_62),
.B(n_90),
.C(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_62),
.B(n_228),
.C(n_230),
.Y(n_227)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_80),
.C(n_85),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_65),
.B(n_340),
.C(n_346),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_65),
.A2(n_78),
.B1(n_340),
.B2(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_69),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_69),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_74),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_74),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_89),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_76),
.B(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_79),
.B(n_89),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_84),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_124),
.C(n_126),
.Y(n_123)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_86),
.B(n_160),
.Y(n_181)
);

XOR2x2_ASAP7_75t_L g431 ( 
.A(n_86),
.B(n_244),
.Y(n_431)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_88),
.Y(n_294)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_88),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_88),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.C(n_95),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_90),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_92),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_92),
.A2(n_230),
.B1(n_355),
.B2(n_357),
.Y(n_354)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_118),
.C(n_122),
.Y(n_100)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_102),
.B(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_116),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_103),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_105),
.B(n_116),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_113),
.Y(n_105)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_109),
.A2(n_110),
.B1(n_302),
.B2(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_119),
.B(n_122),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_123),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_149),
.B1(n_150),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_126),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_126),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_126),
.B(n_187),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_126),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_126),
.A2(n_182),
.B1(n_439),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_128),
.Y(n_286)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_134),
.C(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_143),
.C(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_149),
.B(n_235),
.C(n_246),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_149),
.A2(n_150),
.B1(n_246),
.B2(n_247),
.Y(n_308)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_154),
.B(n_165),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_162),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g564 ( 
.A(n_157),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g562 ( 
.A(n_165),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_167),
.B(n_553),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_257),
.B(n_548),
.Y(n_167)
);

NAND2x1_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_212),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_170),
.A2(n_550),
.B(n_551),
.Y(n_549)
);

NOR2x1_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_171),
.B(n_173),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_209),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_174),
.B(n_210),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_176),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_193),
.C(n_198),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_191),
.Y(n_178)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_182),
.B(n_439),
.Y(n_438)
);

XOR2x1_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_191),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_186),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_187),
.B(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_187),
.A2(n_233),
.B1(n_334),
.B2(n_335),
.Y(n_370)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_190),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_203),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_206),
.Y(n_389)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_255),
.Y(n_212)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_213),
.B(n_255),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.C(n_220),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_218),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_234),
.C(n_250),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_221),
.A2(n_222),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.C(n_231),
.Y(n_222)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_227),
.B(n_231),
.Y(n_325)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_228),
.Y(n_356)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_251),
.B1(n_252),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_235),
.A2(n_236),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.C(n_244),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_240),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_279),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_245),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_249),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_358),
.B(n_539),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_310),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_261),
.B(n_264),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_261),
.B(n_264),
.Y(n_547)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.C(n_275),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_266),
.A2(n_271),
.B1(n_272),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_313),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_298),
.C(n_306),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_287),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g412 ( 
.A(n_278),
.B(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_280),
.A2(n_281),
.B1(n_287),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g402 ( 
.A(n_281),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_285),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_287),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.C(n_295),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.C(n_305),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_302),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_305),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_311),
.A2(n_541),
.B(n_547),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_315),
.B(n_316),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_312),
.B(n_315),
.C(n_316),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.C(n_326),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_319),
.A2(n_320),
.B1(n_323),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_327),
.B(n_419),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_351),
.C(n_354),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_328),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_339),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_364),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_332),
.A2(n_333),
.B1(n_339),
.B2(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_338),
.Y(n_527)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_340),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_345),
.B(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_346),
.B(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_354),
.Y(n_408)
);

XOR2x2_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

NAND3xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_415),
.C(n_421),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_406),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_360),
.B(n_406),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_366),
.C(n_382),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_362),
.A2(n_363),
.B1(n_384),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_366),
.B(n_424),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_424),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.C(n_371),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_367),
.B(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_372),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.C(n_381),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_373),
.B(n_376),
.Y(n_472)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_381),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_397),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_402),
.C(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_390),
.C(n_396),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_386),
.A2(n_387),
.B1(n_390),
.B2(n_391),
.Y(n_445)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_392),
.B(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_402),
.B2(n_405),
.Y(n_397)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_398),
.Y(n_411)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_402),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_410),
.C(n_412),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_416),
.A2(n_544),
.B(n_545),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_417),
.B(n_418),
.Y(n_545)
);

OAI21x1_ASAP7_75t_SL g421 ( 
.A1(n_422),
.A2(n_446),
.B(n_538),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_426),
.B(n_427),
.Y(n_422)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_423),
.B(n_426),
.C(n_427),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.C(n_443),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_444),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.C(n_438),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_432),
.B1(n_433),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_475),
.B(n_537),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_473),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_448),
.B(n_473),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_453),
.C(n_470),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_493),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_453),
.A2(n_454),
.B1(n_471),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_460),
.C(n_465),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_455),
.A2(n_456),
.B1(n_460),
.B2(n_461),
.Y(n_480)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_465),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

OAI21x1_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_495),
.B(n_536),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_492),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_492),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.C(n_484),
.Y(n_477)
);

XNOR2x2_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_533),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_481),
.A2(n_482),
.B1(n_484),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_484),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_489),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_489),
.Y(n_499)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_530),
.B(n_535),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_516),
.B(n_529),
.Y(n_496)
);

NOR2x1_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_509),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_498),
.B(n_509),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_499),
.B(n_502),
.C(n_504),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_501),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_514),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_514),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_523),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_522),
.B(n_528),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_521),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_521),
.Y(n_528)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_532),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_543),
.B(n_546),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_542),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_549),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_556),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_557),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_560),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_562),
.Y(n_560)
);


endmodule