module fake_jpeg_22215_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_42),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_18),
.C(n_31),
.Y(n_63)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_3),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_4),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_17),
.B1(n_15),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_52),
.B1(n_54),
.B2(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_16),
.B1(n_20),
.B2(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_17),
.B1(n_15),
.B2(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_65),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_8),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_33),
.A2(n_18),
.B1(n_32),
.B2(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_40),
.B1(n_47),
.B2(n_31),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_23),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_55),
.B(n_5),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_32),
.B1(n_27),
.B2(n_26),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_95),
.B(n_29),
.C(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_7),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_107),
.B1(n_80),
.B2(n_93),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_23),
.A3(n_51),
.B1(n_49),
.B2(n_29),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_88),
.C(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_29),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_11),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_111),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_4),
.Y(n_111)
);

AO21x2_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_6),
.B(n_7),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_72),
.B1(n_93),
.B2(n_81),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_6),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_75),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_121),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_125),
.B1(n_109),
.B2(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_116),
.B1(n_122),
.B2(n_108),
.Y(n_132)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_113),
.B(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_73),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_98),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_92),
.C(n_78),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_104),
.C(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_133),
.B1(n_143),
.B2(n_117),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_112),
.B1(n_99),
.B2(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_131),
.C(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_141),
.B1(n_144),
.B2(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_82),
.B(n_72),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_115),
.B1(n_76),
.B2(n_126),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_150),
.C(n_135),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_150),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_118),
.C(n_119),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_153),
.C(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_132),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_126),
.B1(n_120),
.B2(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_120),
.C(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_161),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_133),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_130),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_138),
.C(n_137),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_130),
.C(n_106),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_170),
.B(n_172),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_8),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_76),
.C(n_75),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_175),
.C(n_167),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_177),
.B(n_6),
.C(n_86),
.D(n_110),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_164),
.C(n_12),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_86),
.Y(n_179)
);


endmodule