module real_aes_7407_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g222 ( .A1(n_0), .A2(n_223), .B(n_226), .C(n_230), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_1), .B(n_214), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_2), .B(n_224), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_3), .A2(n_184), .B(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_4), .A2(n_216), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g171 ( .A(n_5), .Y(n_171) );
AND2x6_ASAP7_75t_L g189 ( .A(n_5), .B(n_169), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_5), .B(n_515), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_6), .A2(n_189), .B(n_191), .C(n_280), .Y(n_279) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_7), .A2(n_20), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g209 ( .A(n_8), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_9), .B(n_224), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_10), .A2(n_33), .B1(n_158), .B2(n_161), .Y(n_157) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_11), .A2(n_23), .B1(n_91), .B2(n_95), .Y(n_94) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_12), .A2(n_191), .B(n_194), .C(n_202), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_13), .A2(n_25), .B1(n_143), .B2(n_145), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_14), .A2(n_62), .B1(n_102), .B2(n_107), .Y(n_101) );
AOI22xp33_ASAP7_75t_SL g150 ( .A1(n_15), .A2(n_64), .B1(n_151), .B2(n_154), .Y(n_150) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_16), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_17), .A2(n_191), .B(n_202), .C(n_294), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_18), .A2(n_184), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g187 ( .A(n_19), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_21), .A2(n_242), .B(n_243), .C(n_247), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_22), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_22), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_23), .A2(n_39), .B1(n_51), .B2(n_508), .C(n_509), .Y(n_507) );
INVxp67_ASAP7_75t_L g510 ( .A(n_23), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_24), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_26), .B(n_183), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_27), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_27), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_28), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_29), .B(n_224), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_30), .B(n_184), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_31), .B(n_121), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_32), .A2(n_242), .B(n_247), .C(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g227 ( .A(n_34), .Y(n_227) );
INVx1_ASAP7_75t_L g270 ( .A(n_35), .Y(n_270) );
OAI22xp5_ASAP7_75t_SL g502 ( .A1(n_36), .A2(n_71), .B1(n_260), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_36), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_37), .B(n_184), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_38), .Y(n_211) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_39), .A2(n_61), .B1(n_91), .B2(n_95), .Y(n_98) );
INVxp67_ASAP7_75t_L g511 ( .A(n_39), .Y(n_511) );
INVx1_ASAP7_75t_L g169 ( .A(n_40), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_41), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_42), .B(n_184), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_43), .B(n_214), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_44), .A2(n_201), .B(n_257), .C(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g208 ( .A(n_45), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_46), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_47), .B(n_224), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_48), .A2(n_52), .B1(n_125), .B2(n_129), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_49), .B(n_225), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_49), .A2(n_493), .B1(n_506), .B2(n_512), .Y(n_492) );
INVx1_ASAP7_75t_L g521 ( .A(n_49), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_50), .A2(n_76), .B1(n_135), .B2(n_138), .Y(n_134) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_51), .A2(n_68), .B1(n_91), .B2(n_92), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_53), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_54), .B(n_196), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_55), .A2(n_191), .B(n_247), .C(n_310), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_56), .Y(n_255) );
INVx1_ASAP7_75t_L g497 ( .A(n_57), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_58), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_59), .B(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_60), .Y(n_249) );
INVx2_ASAP7_75t_L g206 ( .A(n_63), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_65), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_66), .B(n_229), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_67), .B(n_184), .Y(n_240) );
INVx1_ASAP7_75t_L g244 ( .A(n_69), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_70), .A2(n_80), .B1(n_81), .B2(n_163), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_70), .Y(n_163) );
INVxp67_ASAP7_75t_L g260 ( .A(n_71), .Y(n_260) );
INVx1_ASAP7_75t_L g91 ( .A(n_72), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_72), .Y(n_93) );
INVx1_ASAP7_75t_L g277 ( .A(n_73), .Y(n_277) );
INVx1_ASAP7_75t_L g311 ( .A(n_74), .Y(n_311) );
AND2x2_ASAP7_75t_L g272 ( .A(n_75), .B(n_205), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_164), .B1(n_172), .B2(n_487), .C(n_491), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
OAI322xp33_ASAP7_75t_L g491 ( .A1(n_80), .A2(n_492), .A3(n_516), .B1(n_517), .B2(n_518), .C1(n_521), .C2(n_522), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_SL g82 ( .A(n_83), .B(n_132), .Y(n_82) );
INVxp67_ASAP7_75t_L g517 ( .A(n_83), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_111), .Y(n_83) );
OAI21xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_86), .B(n_101), .Y(n_84) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x6_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
AND2x4_ASAP7_75t_L g108 ( .A(n_89), .B(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_94), .Y(n_89) );
AND2x2_ASAP7_75t_L g106 ( .A(n_90), .B(n_98), .Y(n_106) );
INVx2_ASAP7_75t_L g119 ( .A(n_90), .Y(n_119) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_93), .Y(n_95) );
OR2x2_ASAP7_75t_L g118 ( .A(n_94), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g123 ( .A(n_94), .B(n_119), .Y(n_123) );
INVx2_ASAP7_75t_L g128 ( .A(n_94), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_94), .Y(n_131) );
AND2x6_ASAP7_75t_L g137 ( .A(n_96), .B(n_117), .Y(n_137) );
AND2x2_ASAP7_75t_L g144 ( .A(n_96), .B(n_141), .Y(n_144) );
AND2x4_ASAP7_75t_L g153 ( .A(n_96), .B(n_123), .Y(n_153) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_99), .Y(n_96) );
AND2x2_ASAP7_75t_L g116 ( .A(n_97), .B(n_100), .Y(n_116) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g140 ( .A(n_98), .B(n_110), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_98), .B(n_100), .Y(n_148) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g105 ( .A(n_100), .Y(n_105) );
INVx1_ASAP7_75t_L g110 ( .A(n_100), .Y(n_110) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g127 ( .A(n_105), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g126 ( .A(n_106), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g129 ( .A(n_106), .B(n_130), .Y(n_129) );
BUFx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_120), .C(n_124), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x6_ASAP7_75t_L g122 ( .A(n_116), .B(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g160 ( .A(n_116), .B(n_141), .Y(n_160) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g141 ( .A(n_119), .B(n_128), .Y(n_141) );
BUFx4f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g156 ( .A(n_123), .B(n_140), .Y(n_156) );
BUFx4f_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVxp67_ASAP7_75t_L g516 ( .A(n_132), .Y(n_516) );
NOR2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_149), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_142), .Y(n_133) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx11_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g146 ( .A(n_141), .B(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g161 ( .A(n_147), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_157), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx8_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_SL g165 ( .A(n_166), .B(n_170), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND3x1_ASAP7_75t_SL g506 ( .A(n_167), .B(n_170), .C(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g512 ( .A(n_167), .B(n_513), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_167), .A2(n_489), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_168), .B(n_171), .Y(n_520) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_176), .B(n_423), .Y(n_175) );
NOR5xp2_ASAP7_75t_L g176 ( .A(n_177), .B(n_354), .C(n_383), .D(n_403), .E(n_410), .Y(n_176) );
OAI211xp5_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_234), .B(n_298), .C(n_341), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_179), .A2(n_426), .B1(n_428), .B2(n_429), .Y(n_425) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_213), .Y(n_179) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_180), .Y(n_301) );
AND2x4_ASAP7_75t_L g334 ( .A(n_180), .B(n_335), .Y(n_334) );
INVx5_ASAP7_75t_L g352 ( .A(n_180), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_180), .B(n_353), .Y(n_361) );
AND2x2_ASAP7_75t_L g373 ( .A(n_180), .B(n_238), .Y(n_373) );
AND2x2_ASAP7_75t_L g469 ( .A(n_180), .B(n_337), .Y(n_469) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_210), .Y(n_180) );
AOI21xp5_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_190), .B(n_203), .Y(n_181) );
BUFx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_189), .Y(n_184) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_185), .B(n_189), .Y(n_278) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
INVx1_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g192 ( .A(n_187), .Y(n_192) );
INVx1_ASAP7_75t_L g285 ( .A(n_187), .Y(n_285) );
INVx1_ASAP7_75t_L g193 ( .A(n_188), .Y(n_193) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_188), .Y(n_197) );
INVx3_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
INVx1_ASAP7_75t_L g296 ( .A(n_188), .Y(n_296) );
BUFx3_ASAP7_75t_L g202 ( .A(n_189), .Y(n_202) );
INVx4_ASAP7_75t_SL g232 ( .A(n_189), .Y(n_232) );
INVx5_ASAP7_75t_L g221 ( .A(n_191), .Y(n_221) );
AND2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
BUFx3_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_192), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_198), .B(n_200), .Y(n_194) );
INVx2_ASAP7_75t_L g199 ( .A(n_196), .Y(n_199) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx4_ASAP7_75t_L g258 ( .A(n_197), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_199), .A2(n_244), .B(n_245), .C(n_246), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_199), .A2(n_246), .B(n_270), .C(n_271), .Y(n_269) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_199), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_200), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_202), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g212 ( .A(n_205), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_205), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_205), .A2(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AND2x2_ASAP7_75t_L g217 ( .A(n_206), .B(n_207), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g335 ( .A(n_213), .Y(n_335) );
AND2x2_ASAP7_75t_L g353 ( .A(n_213), .B(n_307), .Y(n_353) );
AND2x2_ASAP7_75t_L g372 ( .A(n_213), .B(n_306), .Y(n_372) );
AND2x2_ASAP7_75t_L g412 ( .A(n_213), .B(n_352), .Y(n_412) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_218), .B(n_233), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_215), .B(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_215), .A2(n_276), .B(n_286), .Y(n_275) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_215), .A2(n_308), .B(n_316), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_215), .B(n_317), .Y(n_316) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_216), .A2(n_292), .B(n_293), .Y(n_291) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B(n_222), .C(n_232), .Y(n_219) );
INVx2_ASAP7_75t_L g242 ( .A(n_221), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_221), .A2(n_232), .B(n_255), .C(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_224), .B(n_260), .Y(n_259) );
INVx5_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx4_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_231), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
INVxp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_262), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AOI322xp5_ASAP7_75t_L g471 ( .A1(n_237), .A2(n_273), .A3(n_326), .B1(n_334), .B2(n_388), .C1(n_472), .C2(n_475), .Y(n_471) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_250), .Y(n_237) );
INVx5_ASAP7_75t_L g303 ( .A(n_238), .Y(n_303) );
AND2x2_ASAP7_75t_L g320 ( .A(n_238), .B(n_305), .Y(n_320) );
BUFx2_ASAP7_75t_L g398 ( .A(n_238), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_238), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g475 ( .A(n_238), .B(n_382), .Y(n_475) );
OR2x6_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_250), .B(n_264), .Y(n_329) );
INVx1_ASAP7_75t_L g356 ( .A(n_250), .Y(n_356) );
AND2x2_ASAP7_75t_L g369 ( .A(n_250), .B(n_289), .Y(n_369) );
AND2x2_ASAP7_75t_L g470 ( .A(n_250), .B(n_388), .Y(n_470) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g324 ( .A(n_251), .B(n_264), .Y(n_324) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
OR2x2_ASAP7_75t_L g339 ( .A(n_251), .B(n_289), .Y(n_339) );
AND2x2_ASAP7_75t_L g349 ( .A(n_251), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_251), .B(n_275), .Y(n_378) );
INVxp67_ASAP7_75t_L g402 ( .A(n_251), .Y(n_402) );
AND2x2_ASAP7_75t_L g409 ( .A(n_251), .B(n_273), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_251), .B(n_289), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_251), .B(n_274), .Y(n_435) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_261), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_257), .A2(n_311), .B(n_312), .C(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_273), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_264), .B(n_290), .Y(n_379) );
OR2x2_ASAP7_75t_L g401 ( .A(n_264), .B(n_274), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_264), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_264), .B(n_369), .Y(n_420) );
OAI211xp5_ASAP7_75t_SL g424 ( .A1(n_264), .A2(n_425), .B(n_430), .C(n_439), .Y(n_424) );
AND2x2_ASAP7_75t_L g485 ( .A(n_264), .B(n_289), .Y(n_485) );
INVx5_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g338 ( .A(n_265), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_265), .B(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_265), .B(n_333), .Y(n_345) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_265), .Y(n_347) );
OR2x2_ASAP7_75t_L g358 ( .A(n_265), .B(n_274), .Y(n_358) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_265), .B(n_349), .Y(n_363) );
AND2x2_ASAP7_75t_L g388 ( .A(n_265), .B(n_274), .Y(n_388) );
AND2x2_ASAP7_75t_L g408 ( .A(n_265), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g446 ( .A(n_265), .B(n_273), .Y(n_446) );
OR2x2_ASAP7_75t_L g449 ( .A(n_265), .B(n_435), .Y(n_449) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_272), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_289), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_274), .A2(n_393), .B(n_396), .C(n_402), .Y(n_392) );
INVx5_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_275), .B(n_289), .Y(n_323) );
AND2x2_ASAP7_75t_L g327 ( .A(n_275), .B(n_290), .Y(n_327) );
OR2x2_ASAP7_75t_L g333 ( .A(n_275), .B(n_289), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_279), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_283), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_283), .A2(n_295), .B(n_297), .Y(n_294) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_SL g350 ( .A(n_289), .Y(n_350) );
OR2x2_ASAP7_75t_L g478 ( .A(n_289), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_318), .B(n_321), .C(n_330), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI31xp33_ASAP7_75t_L g403 ( .A1(n_300), .A2(n_404), .A3(n_406), .B(n_407), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_301), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_302), .B(n_334), .Y(n_340) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_303), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g360 ( .A(n_303), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g365 ( .A(n_303), .B(n_335), .Y(n_365) );
AND2x2_ASAP7_75t_L g375 ( .A(n_303), .B(n_334), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_303), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g395 ( .A(n_303), .B(n_352), .Y(n_395) );
AND2x2_ASAP7_75t_L g400 ( .A(n_303), .B(n_372), .Y(n_400) );
OR2x2_ASAP7_75t_L g419 ( .A(n_303), .B(n_305), .Y(n_419) );
OR2x2_ASAP7_75t_L g421 ( .A(n_303), .B(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_303), .Y(n_468) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g368 ( .A(n_305), .B(n_335), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_305), .B(n_352), .Y(n_391) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_315), .Y(n_308) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g428 ( .A(n_320), .B(n_352), .Y(n_428) );
AOI322xp5_ASAP7_75t_L g430 ( .A1(n_320), .A2(n_334), .A3(n_372), .B1(n_431), .B2(n_432), .C1(n_433), .C2(n_436), .Y(n_430) );
INVx1_ASAP7_75t_L g438 ( .A(n_320), .Y(n_438) );
NAND2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_SL g432 ( .A(n_322), .Y(n_432) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OR2x2_ASAP7_75t_L g384 ( .A(n_323), .B(n_329), .Y(n_384) );
INVx1_ASAP7_75t_L g415 ( .A(n_323), .Y(n_415) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI32xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .A3(n_336), .B1(n_338), .B2(n_340), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AOI21xp33_ASAP7_75t_SL g370 ( .A1(n_333), .A2(n_348), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g385 ( .A(n_334), .Y(n_385) );
AND2x4_ASAP7_75t_L g382 ( .A(n_335), .B(n_352), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_335), .B(n_418), .Y(n_417) );
AOI322xp5_ASAP7_75t_L g447 ( .A1(n_336), .A2(n_363), .A3(n_382), .B1(n_415), .B2(n_448), .C1(n_450), .C2(n_451), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_336), .A2(n_413), .B1(n_477), .B2(n_478), .C(n_480), .Y(n_476) );
AND2x2_ASAP7_75t_L g364 ( .A(n_337), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g344 ( .A(n_339), .Y(n_344) );
OR2x2_ASAP7_75t_L g416 ( .A(n_339), .B(n_401), .Y(n_416) );
OAI31xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .A3(n_346), .B(n_351), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_342), .A2(n_375), .B1(n_376), .B2(n_380), .Y(n_374) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g387 ( .A(n_344), .B(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_346), .A2(n_387), .B1(n_440), .B2(n_443), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g429 ( .A(n_349), .B(n_398), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_349), .B(n_388), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_350), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g463 ( .A(n_350), .B(n_401), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_351), .A2(n_446), .B1(n_459), .B2(n_462), .Y(n_458) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
AND2x2_ASAP7_75t_L g450 ( .A(n_352), .B(n_372), .Y(n_450) );
OR2x2_ASAP7_75t_L g452 ( .A(n_352), .B(n_419), .Y(n_452) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_352), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_353), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_353), .B(n_398), .Y(n_406) );
OAI211xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B(n_362), .C(n_374), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_366), .B2(n_369), .C(n_370), .Y(n_362) );
INVxp67_ASAP7_75t_L g474 ( .A(n_365), .Y(n_474) );
INVx1_ASAP7_75t_L g441 ( .A(n_366), .Y(n_441) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x2_ASAP7_75t_L g405 ( .A(n_367), .B(n_372), .Y(n_405) );
INVx1_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_368), .B(n_395), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g437 ( .A(n_372), .Y(n_437) );
AND2x2_ASAP7_75t_L g443 ( .A(n_372), .B(n_398), .Y(n_443) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g431 ( .A(n_379), .Y(n_431) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_382), .B(n_418), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_386), .B2(n_389), .C(n_392), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g479 ( .A(n_388), .Y(n_479) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_395), .B(n_454), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_401), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g444 ( .A1(n_399), .A2(n_445), .B(n_447), .C(n_453), .Y(n_444) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g456 ( .A(n_401), .Y(n_456) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_416), .B2(n_417), .C1(n_420), .C2(n_421), .Y(n_410) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g486 ( .A(n_417), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_418), .B(n_461), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_418), .A2(n_465), .B1(n_467), .B2(n_470), .Y(n_464) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
NOR4xp25_ASAP7_75t_L g423 ( .A(n_424), .B(n_444), .C(n_457), .D(n_476), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_426), .B(n_456), .Y(n_466) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g433 ( .A(n_431), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_434), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_464), .C(n_471), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g473 ( .A(n_469), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_483), .B(n_486), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_494), .A2(n_506), .B1(n_512), .B2(n_521), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_499), .B1(n_504), .B2(n_505), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_495), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_499), .Y(n_505) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVxp67_ASAP7_75t_L g515 ( .A(n_507), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
endmodule