module fake_jpeg_30955_n_104 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_10),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_23),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_15),
.B1(n_13),
.B2(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_17),
.B1(n_15),
.B2(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_14),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_37),
.B(n_17),
.C(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_37),
.B1(n_36),
.B2(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_47),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_13),
.B1(n_22),
.B2(n_23),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_19),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_34),
.B(n_29),
.C(n_11),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_45),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_34),
.A3(n_12),
.B1(n_16),
.B2(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_56),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_12),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_45),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_51),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_71),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

AO221x1_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_73),
.B1(n_45),
.B2(n_49),
.C(n_46),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_55),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_48),
.C(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_60),
.B1(n_57),
.B2(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_1),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_74),
.B1(n_76),
.B2(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_84),
.B1(n_21),
.B2(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_38),
.C(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_48),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_88),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_33),
.C(n_21),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_90),
.C(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_79),
.B1(n_84),
.B2(n_5),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_6),
.C(n_8),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_2),
.C(n_3),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_94),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_6),
.B1(n_8),
.B2(n_5),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_88),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_98),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_2),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_3),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_5),
.Y(n_104)
);


endmodule