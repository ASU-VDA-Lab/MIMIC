module fake_jpeg_14694_n_243 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_33),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_47),
.B(n_51),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_17),
.B1(n_32),
.B2(n_21),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_27),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_67),
.B1(n_35),
.B2(n_1),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_65),
.B1(n_35),
.B2(n_43),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_26),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_0),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_29),
.B1(n_30),
.B2(n_26),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_66),
.B1(n_59),
.B2(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_90),
.Y(n_112)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_94),
.C(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_92),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_45),
.B1(n_42),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_40),
.B1(n_45),
.B2(n_42),
.Y(n_122)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_98),
.Y(n_108)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_49),
.B1(n_66),
.B2(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_45),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_51),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_111),
.B1(n_122),
.B2(n_95),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_67),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_113),
.C(n_121),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_16),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_107),
.B(n_0),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_43),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_81),
.C(n_101),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_42),
.B1(n_62),
.B2(n_20),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_99),
.B1(n_73),
.B2(n_82),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_62),
.B(n_31),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_84),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_75),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_74),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_86),
.B(n_71),
.C(n_93),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_83),
.B1(n_85),
.B2(n_74),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_84),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_138),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_79),
.B1(n_124),
.B2(n_112),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_24),
.B1(n_3),
.B2(n_4),
.Y(n_173)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_145),
.Y(n_162)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_77),
.B1(n_75),
.B2(n_69),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_62),
.B1(n_23),
.B2(n_20),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_109),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_125),
.C(n_102),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_167),
.C(n_169),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_118),
.C(n_114),
.Y(n_161)
);

OAI322xp33_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_131),
.A3(n_152),
.B1(n_143),
.B2(n_135),
.C1(n_147),
.C2(n_144),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_122),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_108),
.B1(n_123),
.B2(n_23),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_151),
.B1(n_133),
.B2(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_98),
.C(n_62),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_34),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_132),
.B(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_146),
.B1(n_148),
.B2(n_142),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_172),
.B1(n_163),
.B2(n_162),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_13),
.C(n_15),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_87),
.B1(n_24),
.B2(n_31),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_31),
.B1(n_34),
.B2(n_25),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_184),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_31),
.B1(n_25),
.B2(n_5),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_2),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_191),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_169),
.B1(n_167),
.B2(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_174),
.B1(n_165),
.B2(n_11),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_25),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_8),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_154),
.C(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_180),
.C(n_176),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_161),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_201),
.B(n_182),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_176),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_13),
.C(n_15),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_190),
.C(n_192),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_206),
.B(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_209),
.C(n_215),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_175),
.C(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_176),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_193),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_195),
.B1(n_204),
.B2(n_194),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_208),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_217),
.B(n_207),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_209),
.B(n_196),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_225),
.C(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_197),
.C(n_200),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_223),
.B(n_225),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_201),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_221),
.C(n_223),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_231),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_238),
.B(n_231),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_239),
.A2(n_240),
.B(n_233),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_224),
.B(n_15),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);


endmodule