module fake_jpeg_2644_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_23),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_11),
.Y(n_44)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_47),
.B1(n_51),
.B2(n_48),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_38),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_56),
.B1(n_60),
.B2(n_59),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_76),
.B1(n_77),
.B2(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_48),
.B(n_39),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_40),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_56),
.B1(n_39),
.B2(n_47),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_65),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_50),
.B1(n_63),
.B2(n_37),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_50),
.B1(n_37),
.B2(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_38),
.B1(n_41),
.B2(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_93),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_73),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_60),
.C(n_68),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_95),
.C(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_41),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_43),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_45),
.C(n_66),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_102),
.C(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_75),
.B(n_72),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_62),
.B1(n_75),
.B2(n_57),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_105),
.B1(n_111),
.B2(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_75),
.B1(n_34),
.B2(n_33),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_0),
.CI(n_1),
.CON(n_109),
.SN(n_109)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_112),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_31),
.B(n_30),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_124),
.B(n_17),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_99),
.C(n_112),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_126),
.B1(n_109),
.B2(n_5),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_27),
.C(n_26),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_125),
.B1(n_2),
.B2(n_6),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_104),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_24),
.B(n_21),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_109),
.B1(n_4),
.B2(n_5),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_7),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_123),
.B1(n_115),
.B2(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_120),
.C(n_121),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_7),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_132),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_134),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_141),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_127),
.B(n_140),
.C(n_137),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_8),
.B(n_9),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_10),
.B(n_13),
.Y(n_145)
);

AOI321xp33_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_10),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_14),
.Y(n_147)
);


endmodule