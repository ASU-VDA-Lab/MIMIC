module real_jpeg_806_n_5 (n_4, n_0, n_1, n_2, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_5;

wire n_17;
wire n_12;
wire n_8;
wire n_18;
wire n_11;
wire n_14;
wire n_13;
wire n_6;
wire n_7;
wire n_16;
wire n_15;
wire n_10;
wire n_9;

INVx1_ASAP7_75t_SL g10 ( 
.A(n_0),
.Y(n_10)
);

OR2x4_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_12),
.Y(n_11)
);

AO21x1_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_17),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_3),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_10),
.Y(n_9)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g5 ( 
.A(n_6),
.Y(n_5)
);

AOI22xp33_ASAP7_75t_SL g6 ( 
.A1(n_7),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_11),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);


endmodule