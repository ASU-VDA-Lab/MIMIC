module fake_jpeg_18327_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_3),
.B(n_7),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NAND2x1_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_13),
.B1(n_8),
.B2(n_9),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_18),
.B1(n_13),
.B2(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_25),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B1(n_33),
.B2(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_23),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_42),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_33),
.B(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_41),
.B1(n_37),
.B2(n_42),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B(n_5),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_31),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_6),
.B(n_11),
.C(n_39),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_11),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_11),
.Y(n_50)
);


endmodule