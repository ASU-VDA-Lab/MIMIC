module fake_jpeg_7713_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_28),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_47),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_18),
.B1(n_26),
.B2(n_17),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_37),
.B1(n_18),
.B2(n_26),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_30),
.B1(n_28),
.B2(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_25),
.B1(n_20),
.B2(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_63),
.B1(n_68),
.B2(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_24),
.B1(n_29),
.B2(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_61),
.B1(n_20),
.B2(n_22),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_24),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_25),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_29),
.B1(n_18),
.B2(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_27),
.Y(n_93)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_81),
.B1(n_83),
.B2(n_61),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_26),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_22),
.B1(n_19),
.B2(n_31),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_57),
.B1(n_70),
.B2(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_47),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_32),
.B1(n_26),
.B2(n_50),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_48),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_48),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_100),
.B(n_87),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_46),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_0),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_68),
.B1(n_62),
.B2(n_56),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_106),
.B1(n_108),
.B2(n_112),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_72),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_45),
.B1(n_57),
.B2(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_104),
.B1(n_113),
.B2(n_118),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_59),
.B1(n_57),
.B2(n_48),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_49),
.B1(n_50),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_32),
.B1(n_66),
.B2(n_54),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_132),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_112),
.Y(n_154)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_131),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_78),
.B1(n_90),
.B2(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_111),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_42),
.C(n_51),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_92),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_106),
.B1(n_109),
.B2(n_116),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_134),
.B1(n_104),
.B2(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_93),
.B1(n_73),
.B2(n_54),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_73),
.B1(n_66),
.B2(n_89),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_95),
.A2(n_60),
.B1(n_64),
.B2(n_51),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_66),
.B1(n_89),
.B2(n_71),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_64),
.B(n_60),
.C(n_71),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_142),
.B(n_26),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_40),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_42),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_94),
.A2(n_98),
.B1(n_96),
.B2(n_118),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_100),
.C(n_110),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_167),
.C(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_153),
.B1(n_159),
.B2(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_94),
.B1(n_96),
.B2(n_112),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_159),
.Y(n_190)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_163),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_94),
.B1(n_96),
.B2(n_95),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_0),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_138),
.B(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_51),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_95),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_51),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_11),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_141),
.B1(n_120),
.B2(n_133),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_189),
.B1(n_32),
.B2(n_79),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_185),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_124),
.B1(n_142),
.B2(n_137),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_188),
.C(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_122),
.B1(n_126),
.B2(n_132),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_174),
.B1(n_175),
.B2(n_187),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_153),
.B1(n_155),
.B2(n_160),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_126),
.C(n_121),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_163),
.B1(n_148),
.B2(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_134),
.C(n_131),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_193),
.C(n_149),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_120),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_160),
.B(n_153),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_138),
.B(n_139),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_161),
.B(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_198),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

NOR4xp25_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_173),
.C(n_171),
.D(n_164),
.Y(n_199)
);

AOI211xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_181),
.B(n_32),
.C(n_10),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_206),
.C(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_212),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_181),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_151),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_150),
.B(n_146),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_151),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_205),
.B1(n_174),
.B2(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_216),
.B1(n_218),
.B2(n_194),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_156),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_165),
.C(n_41),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_79),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_32),
.C(n_3),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_183),
.C(n_172),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_231),
.B1(n_236),
.B2(n_9),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_238),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_196),
.B1(n_182),
.B2(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_235),
.C(n_202),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_183),
.B1(n_173),
.B2(n_176),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_233),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_32),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_214),
.C(n_211),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_208),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_16),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_244),
.C(n_246),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_251),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_225),
.C(n_237),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_15),
.Y(n_248)
);

FAx1_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_12),
.CI(n_9),
.CON(n_262),
.SN(n_262)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_2),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_13),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_13),
.CI(n_12),
.CON(n_251),
.SN(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_252),
.B(n_232),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_12),
.B1(n_9),
.B2(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_225),
.C(n_228),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_241),
.Y(n_268)
);

AOI211xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_231),
.B(n_229),
.C(n_236),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_245),
.B1(n_247),
.B2(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_265),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_234),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_228),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_270),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_273),
.A3(n_243),
.B1(n_249),
.B2(n_6),
.C1(n_7),
.C2(n_2),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_248),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_243),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_249),
.C(n_6),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_250),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_272),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_253),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_255),
.B1(n_245),
.B2(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_282),
.Y(n_284)
);

OAI31xp33_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_263),
.A3(n_249),
.B(n_262),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_288),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_278),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_292),
.B(n_289),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.C(n_291),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_287),
.B(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_283),
.Y(n_298)
);


endmodule