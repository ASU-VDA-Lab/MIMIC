module real_jpeg_1588_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_58),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_0),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_0),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_2),
.B(n_65),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_167),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_2),
.A2(n_32),
.B(n_33),
.C(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_38),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_217),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_52),
.C(n_55),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_2),
.B(n_94),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_2),
.B(n_83),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_126),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_126),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_6),
.A2(n_44),
.B1(n_55),
.B2(n_56),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_7),
.A2(n_47),
.B1(n_65),
.B2(n_66),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_159)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g343 ( 
.A(n_11),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_11),
.B(n_345),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_60),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_12),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_13),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_166),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_166),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_166),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_15),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_16),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_104),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_16),
.A2(n_39),
.B1(n_40),
.B2(n_104),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_16),
.A2(n_55),
.B1(n_56),
.B2(n_104),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_17),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_17),
.A2(n_39),
.B1(n_40),
.B2(n_68),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_343),
.B(n_344),
.Y(n_19)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_338),
.B(n_341),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_330),
.B(n_334),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_317),
.B(n_329),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_142),
.B(n_314),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_129),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_105),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_26),
.B(n_105),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_86),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_61),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_28),
.A2(n_29),
.B(n_48),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_28),
.B(n_61),
.C(n_86),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_48),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_30),
.A2(n_45),
.B1(n_46),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_30),
.A2(n_43),
.B1(n_45),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_30),
.A2(n_45),
.B1(n_80),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_30),
.A2(n_183),
.B(n_185),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_30),
.A2(n_185),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_31),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_31),
.A2(n_38),
.B1(n_184),
.B2(n_201),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_31),
.A2(n_38),
.B(n_321),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B(n_37),
.C(n_38),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_34),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g187 ( 
.A1(n_33),
.A2(n_66),
.A3(n_72),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_34),
.B(n_73),
.Y(n_189)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_38),
.B(n_163),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_39),
.A2(n_42),
.B(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_40),
.B(n_262),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_45),
.A2(n_122),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_45),
.A2(n_162),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_54),
.B1(n_57),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_49),
.A2(n_54),
.B1(n_210),
.B2(n_244),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_49),
.A2(n_212),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_50),
.A2(n_83),
.B1(n_99),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_50),
.A2(n_83),
.B1(n_120),
.B2(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_50),
.A2(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_50),
.B(n_213),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_54),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_54),
.A2(n_233),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_55),
.B(n_273),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_77),
.B2(n_85),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_63),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g140 ( 
.A(n_63),
.B(n_78),
.C(n_82),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_63),
.B(n_133),
.C(n_140),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_71),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_75)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_66),
.A2(n_69),
.B(n_217),
.C(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_124),
.B(n_127),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_70),
.A2(n_125),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_70),
.A2(n_167),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_70),
.A2(n_167),
.B1(n_324),
.B2(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_70),
.A2(n_167),
.B(n_332),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_71),
.A2(n_101),
.B(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_81),
.A2(n_82),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_82),
.B(n_134),
.C(n_138),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_83),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_100),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_88),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_90),
.B1(n_100),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_89),
.A2(n_90),
.B1(n_97),
.B2(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_94),
.B(n_95),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_91),
.A2(n_94),
.B1(n_117),
.B2(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_91),
.A2(n_217),
.B(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_92),
.A2(n_93),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_92),
.A2(n_93),
.B1(n_192),
.B2(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_92),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_92),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_92),
.A2(n_93),
.B1(n_248),
.B2(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_93),
.A2(n_207),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_93),
.B(n_221),
.Y(n_250)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_94),
.A2(n_220),
.B(n_277),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_97),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_121),
.C(n_123),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_114),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_128),
.B(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_129),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_130),
.B(n_141),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_135),
.Y(n_323)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_139),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_168),
.B(n_313),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_144),
.B(n_147),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_153),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.C(n_164),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_155),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_156),
.B(n_158),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_157),
.Y(n_232)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_194),
.B(n_312),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_170),
.B(n_172),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.C(n_179),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_173),
.B(n_177),
.Y(n_297)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_186),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_180),
.B(n_182),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_186),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI31xp33_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_294),
.A3(n_304),
.B(n_309),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_238),
.B(n_293),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_222),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_197),
.B(n_222),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_208),
.C(n_214),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_198),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_203),
.C(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_208),
.B(n_214),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_218),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_223),
.B(n_235),
.C(n_237),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_224),
.B(n_229),
.C(n_230),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_288),
.B(n_292),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_257),
.B(n_287),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_251),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_251),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_247),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_255),
.C(n_256),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_269),
.B(n_286),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_265),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_280),
.B(n_285),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_275),
.B(n_279),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_278),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_283),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_298),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_308),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_328),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_327),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_322),
.B1(n_325),
.B2(n_326),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_320),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_325),
.C(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_331),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_331),
.B(n_339),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_336),
.B(n_340),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);


endmodule