module fake_netlist_6_884_n_1644 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1644);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1644;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

BUFx2_ASAP7_75t_SL g154 ( 
.A(n_32),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_27),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_79),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_41),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_14),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_53),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_26),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_55),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_92),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_66),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_41),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_37),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_37),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_120),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_18),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_56),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_147),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_28),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_146),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_32),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_27),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_76),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_73),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_9),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_95),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_58),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_94),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_10),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_68),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_28),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_75),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_25),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_24),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_107),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_64),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_23),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_57),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_49),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_5),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_11),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_20),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_130),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_49),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_96),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_11),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_22),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_69),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_23),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_84),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_9),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_10),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_142),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_100),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_46),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_67),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_117),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_110),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_45),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_71),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_2),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_62),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_39),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_132),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_22),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_70),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_44),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_16),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_35),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_12),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_35),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_65),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_103),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_24),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_1),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_91),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_42),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_128),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_29),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_34),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_89),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_151),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_31),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_136),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_54),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_26),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_60),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_139),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_33),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_85),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_78),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_140),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_152),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_39),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_104),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_221),
.B(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_198),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_197),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_202),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_209),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_203),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_208),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_162),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_211),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_154),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_217),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_209),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_209),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_269),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_224),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_209),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_226),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_231),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_172),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_160),
.B(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_172),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_233),
.Y(n_325)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_162),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_200),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_201),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_280),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_206),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_205),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_206),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_237),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_221),
.B(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_242),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_216),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_168),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_254),
.Y(n_341)
);

BUFx6f_ASAP7_75t_SL g342 ( 
.A(n_153),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_176),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_160),
.B(n_6),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_247),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_171),
.B(n_191),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_168),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_259),
.B(n_6),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_291),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_250),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_210),
.B(n_141),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_153),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_248),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_171),
.B(n_7),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_191),
.B(n_272),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_253),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_230),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_153),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_230),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_R g364 ( 
.A(n_155),
.B(n_8),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_300),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_170),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_189),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_238),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_238),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_190),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_155),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_157),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_305),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_R g379 ( 
.A(n_351),
.B(n_156),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_302),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_303),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_314),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_210),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_329),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_304),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_308),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_287),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_355),
.B(n_182),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_192),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_373),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_369),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_309),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_287),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_332),
.A2(n_165),
.B1(n_278),
.B2(n_298),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_368),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_311),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_156),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_354),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_272),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_338),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_313),
.B(n_195),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_307),
.A2(n_227),
.B1(n_292),
.B2(n_289),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_324),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_374),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_317),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_341),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_319),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_320),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_347),
.B(n_256),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_357),
.B(n_158),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_349),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_325),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_331),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_333),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_334),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_337),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_355),
.B(n_182),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_337),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_368),
.B(n_161),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_339),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_370),
.B(n_161),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_398),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_336),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_431),
.B(n_316),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_394),
.B(n_159),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_370),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_345),
.Y(n_456)
);

BUFx10_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_356),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_378),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_396),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_410),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_414),
.B(n_316),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_381),
.B(n_366),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_376),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_376),
.Y(n_469)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_394),
.A2(n_323),
.B1(n_344),
.B2(n_301),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_391),
.B(n_330),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_377),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_415),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_394),
.A2(n_301),
.B1(n_335),
.B2(n_348),
.Y(n_477)
);

INVx4_ASAP7_75t_SL g478 ( 
.A(n_414),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_388),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_363),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_403),
.B(n_330),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_404),
.A2(n_167),
.B1(n_178),
.B2(n_299),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_404),
.B(n_163),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_404),
.B(n_362),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_383),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_407),
.B(n_359),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_404),
.B(n_312),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_385),
.B(n_173),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_399),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_416),
.A2(n_246),
.B1(n_180),
.B2(n_286),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_427),
.B(n_365),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_385),
.B(n_174),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_412),
.B(n_371),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_378),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_378),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_371),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_429),
.B(n_182),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_416),
.B(n_177),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_430),
.B(n_164),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_388),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_395),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_380),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_436),
.B(n_342),
.Y(n_511)
);

BUFx4f_ASAP7_75t_L g512 ( 
.A(n_388),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_416),
.A2(n_251),
.B1(n_187),
.B2(n_283),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_380),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_440),
.B(n_164),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_433),
.B(n_183),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_433),
.A2(n_277),
.B1(n_212),
.B2(n_261),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_433),
.A2(n_243),
.B1(n_240),
.B2(n_215),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_408),
.B(n_379),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_408),
.B(n_166),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_434),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_434),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_384),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_426),
.B(n_166),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_384),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_389),
.Y(n_528)
);

INVx6_ASAP7_75t_L g529 ( 
.A(n_433),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_389),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_411),
.B(n_339),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_L g532 ( 
.A(n_444),
.B(n_446),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

AO21x2_ASAP7_75t_L g534 ( 
.A1(n_444),
.A2(n_220),
.B(n_194),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_390),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_446),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_390),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_406),
.B(n_184),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_397),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_401),
.B(n_175),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_425),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_425),
.B(n_213),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

AND2x2_ASAP7_75t_SL g546 ( 
.A(n_402),
.B(n_175),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_442),
.B(n_342),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_R g550 ( 
.A(n_406),
.B(n_169),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_420),
.B(n_399),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_417),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_409),
.B(n_342),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_413),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_445),
.A2(n_270),
.B1(n_267),
.B2(n_441),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_413),
.B(n_239),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_421),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_421),
.B(n_249),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_422),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_405),
.B(n_169),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_432),
.B(n_179),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_386),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_405),
.B(n_364),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_441),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_443),
.B(n_268),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_423),
.B(n_175),
.Y(n_568)
);

INVxp33_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_423),
.B(n_297),
.C(n_290),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_423),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_424),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_424),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_424),
.B(n_350),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_437),
.B(n_274),
.Y(n_576)
);

AOI21x1_ASAP7_75t_L g577 ( 
.A1(n_437),
.A2(n_439),
.B(n_438),
.Y(n_577)
);

OAI21xp33_ASAP7_75t_SL g578 ( 
.A1(n_438),
.A2(n_353),
.B(n_352),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_438),
.A2(n_175),
.B1(n_207),
.B2(n_244),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_439),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_418),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_428),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_439),
.B(n_353),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_435),
.B(n_204),
.C(n_214),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_447),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_537),
.B(n_179),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_577),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_479),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_577),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_449),
.A2(n_288),
.B(n_294),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_479),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_520),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_501),
.B(n_175),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_479),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_501),
.B(n_207),
.Y(n_596)
);

AOI221xp5_ASAP7_75t_L g597 ( 
.A1(n_533),
.A2(n_263),
.B1(n_298),
.B2(n_292),
.C(n_289),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_523),
.B(n_350),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_546),
.B(n_207),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_545),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_546),
.B(n_244),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_538),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_531),
.B(n_244),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_449),
.B(n_176),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_448),
.B(n_181),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_531),
.B(n_181),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_545),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_557),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_541),
.B(n_352),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_498),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_559),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_538),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_449),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_478),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_534),
.A2(n_176),
.B1(n_279),
.B2(n_278),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_457),
.B(n_185),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_467),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_574),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_498),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_478),
.B(n_176),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_471),
.B(n_477),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_478),
.B(n_176),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_478),
.B(n_176),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_583),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_559),
.Y(n_627)
);

NOR3xp33_ASAP7_75t_L g628 ( 
.A(n_458),
.B(n_252),
.C(n_193),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_492),
.A2(n_497),
.B(n_452),
.C(n_486),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_569),
.B(n_196),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_536),
.B(n_176),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_554),
.B(n_186),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_534),
.A2(n_264),
.B1(n_265),
.B2(n_271),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_457),
.B(n_260),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_583),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_554),
.B(n_260),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_536),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_456),
.A2(n_507),
.B(n_491),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_527),
.B(n_262),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_454),
.B(n_266),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_527),
.B(n_528),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_452),
.A2(n_296),
.B(n_295),
.C(n_293),
.Y(n_642)
);

BUFx12f_ASAP7_75t_L g643 ( 
.A(n_581),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_451),
.B(n_266),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_527),
.B(n_276),
.Y(n_645)
);

AOI22x1_ASAP7_75t_L g646 ( 
.A1(n_536),
.A2(n_296),
.B1(n_295),
.B2(n_293),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_540),
.A2(n_276),
.B1(n_282),
.B2(n_281),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_528),
.B(n_282),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_487),
.B(n_457),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_488),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_494),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_528),
.B(n_199),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_494),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_457),
.B(n_241),
.Y(n_654)
);

BUFx4_ASAP7_75t_L g655 ( 
.A(n_581),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_560),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_475),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_475),
.B(n_285),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_452),
.B(n_245),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_452),
.B(n_236),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_540),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_494),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_568),
.B(n_235),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_475),
.B(n_285),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_486),
.B(n_234),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_526),
.B(n_232),
.Y(n_667)
);

AND2x2_ASAP7_75t_SL g668 ( 
.A(n_568),
.B(n_98),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_552),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_552),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_552),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_581),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_523),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_564),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_464),
.B(n_257),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_571),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_550),
.B(n_229),
.C(n_219),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_564),
.B(n_218),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_548),
.B(n_466),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_568),
.B(n_222),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_566),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_475),
.B(n_279),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_566),
.B(n_225),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_522),
.B(n_223),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_573),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_509),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_509),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_470),
.B(n_275),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_483),
.B(n_275),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_524),
.B(n_273),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_489),
.B(n_273),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_514),
.B(n_271),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_514),
.B(n_265),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_506),
.B(n_264),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_524),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_534),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_516),
.B(n_15),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_503),
.B(n_15),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_515),
.B(n_81),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_515),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_483),
.B(n_16),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_453),
.B(n_17),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_493),
.B(n_17),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_525),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_504),
.A2(n_21),
.B(n_30),
.C(n_36),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_530),
.B(n_88),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_535),
.B(n_83),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_562),
.B(n_21),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_535),
.B(n_90),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_539),
.B(n_36),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_561),
.B(n_38),
.C(n_40),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_529),
.B(n_102),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_517),
.A2(n_93),
.B(n_131),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_529),
.A2(n_80),
.B1(n_125),
.B2(n_123),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_539),
.B(n_38),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_539),
.B(n_42),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_539),
.B(n_43),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_529),
.B(n_549),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_455),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_556),
.B(n_105),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_529),
.B(n_72),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_549),
.B(n_106),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_549),
.B(n_134),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_543),
.B(n_121),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_581),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_582),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_543),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_549),
.B(n_119),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_511),
.B(n_43),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_455),
.B(n_115),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

INVx8_ASAP7_75t_L g732 ( 
.A(n_539),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_455),
.B(n_108),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_551),
.B(n_50),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_459),
.Y(n_735)
);

BUFx12f_ASAP7_75t_L g736 ( 
.A(n_582),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_459),
.B(n_51),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_582),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_605),
.B(n_556),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_696),
.A2(n_551),
.B1(n_485),
.B2(n_513),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_585),
.B(n_484),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_718),
.A2(n_512),
.B(n_481),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_708),
.A2(n_565),
.B(n_553),
.C(n_556),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_605),
.B(n_584),
.C(n_472),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_623),
.A2(n_616),
.B1(n_668),
.B2(n_697),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_611),
.B(n_563),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_587),
.A2(n_461),
.B(n_465),
.Y(n_747)
);

AOI21x1_ASAP7_75t_L g748 ( 
.A1(n_604),
.A2(n_544),
.B(n_460),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_650),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_592),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_668),
.B(n_582),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_614),
.A2(n_638),
.B(n_629),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_673),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_614),
.A2(n_512),
.B(n_481),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_614),
.A2(n_512),
.B(n_481),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_649),
.B(n_521),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_615),
.B(n_500),
.Y(n_757)
);

AO21x1_ASAP7_75t_L g758 ( 
.A1(n_599),
.A2(n_558),
.B(n_576),
.Y(n_758)
);

NAND3xp33_ASAP7_75t_L g759 ( 
.A(n_586),
.B(n_691),
.C(n_644),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_589),
.A2(n_474),
.B(n_450),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_620),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_626),
.B(n_500),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_588),
.B(n_567),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_618),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_592),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_593),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_626),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_601),
.A2(n_462),
.B(n_450),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_643),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_697),
.A2(n_518),
.B(n_519),
.C(n_570),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_635),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_618),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_664),
.A2(n_578),
.B(n_567),
.C(n_575),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_695),
.B(n_496),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_635),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_609),
.B(n_495),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_641),
.A2(n_502),
.B(n_500),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_630),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_664),
.A2(n_578),
.B(n_567),
.C(n_575),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_600),
.B(n_607),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_608),
.B(n_500),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_610),
.B(n_459),
.Y(n_782)
);

OAI21xp33_ASAP7_75t_L g783 ( 
.A1(n_586),
.A2(n_555),
.B(n_567),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_612),
.B(n_543),
.Y(n_784)
);

AO22x1_ASAP7_75t_L g785 ( 
.A1(n_698),
.A2(n_542),
.B1(n_543),
.B2(n_462),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_712),
.A2(n_502),
.B(n_499),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_588),
.A2(n_567),
.B1(n_579),
.B2(n_543),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_593),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_603),
.A2(n_460),
.B(n_473),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_684),
.A2(n_570),
.B(n_499),
.C(n_547),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_725),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_602),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_591),
.B(n_499),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_721),
.A2(n_482),
.B(n_510),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_649),
.B(n_580),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_602),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_627),
.B(n_656),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_580),
.Y(n_798)
);

OAI321xp33_ASAP7_75t_L g799 ( 
.A1(n_696),
.A2(n_480),
.A3(n_508),
.B1(n_505),
.B2(n_463),
.C(n_468),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_594),
.A2(n_476),
.B(n_505),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_674),
.B(n_580),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_596),
.A2(n_723),
.B(n_722),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_616),
.A2(n_580),
.B1(n_572),
.B2(n_547),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_681),
.B(n_572),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_R g805 ( 
.A(n_657),
.B(n_572),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_686),
.B(n_687),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_613),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_728),
.A2(n_473),
.B(n_490),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_700),
.B(n_572),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_684),
.A2(n_547),
.B(n_468),
.C(n_463),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_618),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_704),
.B(n_547),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_606),
.B(n_469),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_727),
.A2(n_542),
.B(n_52),
.Y(n_815)
);

AND2x2_ASAP7_75t_SL g816 ( 
.A(n_658),
.B(n_51),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_732),
.B(n_52),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_637),
.A2(n_53),
.B1(n_542),
.B2(n_595),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_679),
.B(n_542),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_720),
.A2(n_542),
.B(n_652),
.Y(n_820)
);

AND2x6_ASAP7_75t_SL g821 ( 
.A(n_698),
.B(n_542),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_669),
.A2(n_670),
.B(n_671),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_598),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_654),
.B(n_621),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_719),
.Y(n_825)
);

O2A1O1Ixp5_ASAP7_75t_L g826 ( 
.A1(n_680),
.A2(n_678),
.B(n_683),
.C(n_625),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_714),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_632),
.B(n_636),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_669),
.A2(n_670),
.B(n_671),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_633),
.A2(n_734),
.B1(n_716),
.B2(n_715),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_710),
.A2(n_717),
.B1(n_715),
.B2(n_716),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_690),
.B(n_688),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_639),
.B(n_645),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_648),
.A2(n_631),
.B(n_699),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_631),
.A2(n_709),
.B(n_706),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_710),
.A2(n_717),
.B(n_642),
.C(n_693),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_707),
.A2(n_730),
.B(n_733),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_633),
.A2(n_701),
.B1(n_694),
.B2(n_667),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_640),
.B(n_598),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_654),
.B(n_675),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_622),
.A2(n_624),
.B(n_666),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_675),
.A2(n_694),
.B1(n_644),
.B2(n_667),
.Y(n_842)
);

NOR2x1_ASAP7_75t_L g843 ( 
.A(n_725),
.B(n_738),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_640),
.B(n_692),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_659),
.B(n_661),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_732),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_732),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_711),
.A2(n_628),
.B1(n_701),
.B2(n_713),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_651),
.A2(n_663),
.B(n_653),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_651),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_662),
.A2(n_647),
.B(n_737),
.C(n_597),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_676),
.B(n_685),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_617),
.B(n_634),
.Y(n_854)
);

INVxp33_ASAP7_75t_SL g855 ( 
.A(n_665),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_729),
.A2(n_646),
.B1(n_731),
.B2(n_685),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_705),
.A2(n_689),
.B(n_702),
.C(n_590),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_703),
.B(n_682),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_677),
.A2(n_726),
.B(n_738),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_726),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_672),
.A2(n_655),
.B(n_643),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_736),
.A2(n_449),
.B(n_467),
.Y(n_862)
);

OAI21xp33_ASAP7_75t_L g863 ( 
.A1(n_736),
.A2(n_447),
.B(n_431),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_618),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_585),
.B(n_447),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_605),
.B(n_447),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_585),
.B(n_609),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_605),
.B(n_447),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_605),
.B(n_447),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_698),
.B(n_489),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_673),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_605),
.B(n_447),
.Y(n_874)
);

CKINVDCx6p67_ASAP7_75t_R g875 ( 
.A(n_643),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_619),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_605),
.B(n_447),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_L g878 ( 
.A(n_679),
.B(n_447),
.C(n_458),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_708),
.A2(n_447),
.B(n_623),
.C(n_664),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_619),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_623),
.A2(n_447),
.B1(n_629),
.B2(n_414),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_605),
.B(n_447),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_649),
.A2(n_532),
.B1(n_447),
.B2(n_605),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_585),
.B(n_447),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_605),
.B(n_447),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_587),
.A2(n_589),
.B(n_629),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_605),
.B(n_447),
.Y(n_890)
);

AOI22x1_ASAP7_75t_L g891 ( 
.A1(n_637),
.A2(n_638),
.B1(n_735),
.B2(n_719),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_605),
.B(n_447),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_605),
.B(n_447),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_618),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_605),
.B(n_447),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_592),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_718),
.A2(n_449),
.B(n_467),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_611),
.B(n_447),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_618),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_696),
.A2(n_447),
.B1(n_623),
.B2(n_668),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_842),
.A2(n_838),
.B(n_840),
.C(n_866),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_868),
.B(n_870),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_887),
.B(n_874),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_877),
.B(n_885),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_752),
.A2(n_802),
.B(n_837),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_882),
.A2(n_739),
.B(n_747),
.Y(n_909)
);

BUFx5_ASAP7_75t_L g910 ( 
.A(n_844),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_860),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_912)
);

OAI21x1_ASAP7_75t_L g913 ( 
.A1(n_808),
.A2(n_891),
.B(n_786),
.Y(n_913)
);

NAND2x1_ASAP7_75t_L g914 ( 
.A(n_772),
.B(n_809),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_850),
.A2(n_777),
.B(n_748),
.Y(n_915)
);

AOI21xp33_ASAP7_75t_L g916 ( 
.A1(n_838),
.A2(n_903),
.B(n_890),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_761),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_760),
.A2(n_835),
.B(n_889),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_888),
.B(n_892),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_869),
.A2(n_880),
.B(n_871),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_893),
.B(n_895),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_820),
.A2(n_834),
.B(n_742),
.Y(n_922)
);

OAI21x1_ASAP7_75t_SL g923 ( 
.A1(n_758),
.A2(n_846),
.B(n_862),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_865),
.B(n_867),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_903),
.B(n_878),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_754),
.A2(n_755),
.B(n_828),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_768),
.A2(n_789),
.B(n_800),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_741),
.B(n_832),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_886),
.B(n_824),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_776),
.B(n_858),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_901),
.B(n_833),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_883),
.A2(n_899),
.B(n_896),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_884),
.A2(n_900),
.B(n_897),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_745),
.A2(n_879),
.B(n_836),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_839),
.B(n_847),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_759),
.B(n_744),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_774),
.B(n_778),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_768),
.A2(n_826),
.B(n_789),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_783),
.A2(n_849),
.B(n_854),
.C(n_852),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_830),
.A2(n_831),
.B1(n_740),
.B2(n_751),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_845),
.B(n_767),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_771),
.B(n_775),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_799),
.A2(n_800),
.B(n_841),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_876),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_881),
.B(n_814),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_740),
.B(n_830),
.C(n_863),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_812),
.B(n_772),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_853),
.A2(n_784),
.B(n_779),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_770),
.A2(n_827),
.B1(n_816),
.B2(n_806),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_773),
.A2(n_757),
.B(n_813),
.Y(n_950)
);

AO31x2_ASAP7_75t_L g951 ( 
.A1(n_811),
.A2(n_790),
.A3(n_743),
.B(n_818),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_757),
.A2(n_804),
.B(n_801),
.Y(n_952)
);

AND2x6_ASAP7_75t_SL g953 ( 
.A(n_817),
.B(n_839),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_R g954 ( 
.A(n_749),
.B(n_751),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_799),
.A2(n_762),
.B(n_803),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_857),
.A2(n_819),
.B(n_782),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_780),
.B(n_797),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_798),
.A2(n_810),
.B(n_825),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_860),
.B(n_861),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_764),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_847),
.B(n_848),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_753),
.B(n_855),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_788),
.B(n_807),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_812),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_825),
.A2(n_781),
.B(n_851),
.Y(n_965)
);

AND3x2_ASAP7_75t_L g966 ( 
.A(n_873),
.B(n_823),
.C(n_763),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_796),
.A2(n_795),
.B(n_750),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_765),
.A2(n_898),
.B(n_792),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_766),
.A2(n_787),
.B(n_856),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_L g970 ( 
.A1(n_756),
.A2(n_753),
.B1(n_746),
.B2(n_791),
.C(n_859),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_894),
.A2(n_815),
.B(n_843),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_763),
.B(n_894),
.Y(n_972)
);

AND3x2_ASAP7_75t_L g973 ( 
.A(n_769),
.B(n_875),
.C(n_872),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_793),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_860),
.B(n_817),
.Y(n_975)
);

AO21x1_ASAP7_75t_L g976 ( 
.A1(n_793),
.A2(n_809),
.B(n_821),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_764),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_812),
.A2(n_785),
.B(n_902),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_902),
.B(n_764),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_864),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_812),
.A2(n_864),
.B(n_902),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_817),
.B(n_847),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_864),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_848),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_848),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_769),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_805),
.A2(n_829),
.B(n_822),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_838),
.A2(n_903),
.B(n_745),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_866),
.B(n_447),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_838),
.A2(n_842),
.B(n_903),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_812),
.B(n_772),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_851),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_842),
.B(n_838),
.C(n_447),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_749),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_842),
.B(n_838),
.C(n_447),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_761),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_842),
.A2(n_838),
.B(n_840),
.C(n_866),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_887),
.B(n_866),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_887),
.B(n_866),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_749),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_839),
.B(n_847),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_867),
.B(n_585),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_842),
.A2(n_838),
.B(n_840),
.C(n_866),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_887),
.B(n_866),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_1007)
);

NAND2x1p5_ASAP7_75t_L g1008 ( 
.A(n_812),
.B(n_772),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_860),
.B(n_732),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_867),
.B(n_585),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_887),
.B(n_866),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_759),
.B(n_901),
.Y(n_1013)
);

OAI22x1_ASAP7_75t_L g1014 ( 
.A1(n_842),
.A2(n_759),
.B1(n_824),
.B2(n_561),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_887),
.B(n_866),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_753),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_842),
.A2(n_838),
.B1(n_840),
.B2(n_759),
.Y(n_1017)
);

AOI221x1_ASAP7_75t_L g1018 ( 
.A1(n_838),
.A2(n_903),
.B1(n_840),
.B2(n_830),
.C(n_759),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_887),
.B(n_866),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_842),
.A2(n_838),
.B(n_840),
.C(n_866),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_840),
.A2(n_838),
.B(n_868),
.C(n_866),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_866),
.B(n_868),
.Y(n_1022)
);

INVx6_ASAP7_75t_L g1023 ( 
.A(n_860),
.Y(n_1023)
);

INVxp67_ASAP7_75t_SL g1024 ( 
.A(n_764),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_867),
.B(n_585),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_761),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_842),
.A2(n_838),
.B(n_840),
.C(n_866),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_746),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_768),
.A2(n_889),
.B(n_789),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_822),
.A2(n_829),
.B(n_794),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_753),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_842),
.B(n_840),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_866),
.B(n_868),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_753),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_911),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_917),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_944),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_931),
.B(n_930),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_989),
.A2(n_997),
.B(n_994),
.C(n_988),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_1033),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_SL g1043 ( 
.A(n_990),
.B(n_988),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_1036),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_928),
.B(n_1004),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_908),
.A2(n_909),
.B(n_918),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1010),
.B(n_1025),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_982),
.B(n_959),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_1016),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_935),
.B(n_1003),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_907),
.B(n_919),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_998),
.Y(n_1052)
);

AOI222xp33_ASAP7_75t_L g1053 ( 
.A1(n_940),
.A2(n_946),
.B1(n_1034),
.B2(n_1020),
.C1(n_1029),
.C2(n_904),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_982),
.B(n_959),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_907),
.B(n_919),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_1030),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_937),
.B(n_1022),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_970),
.B(n_906),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_1023),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_906),
.B(n_1000),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1001),
.B(n_1006),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_984),
.B(n_961),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_990),
.A2(n_934),
.B(n_1005),
.Y(n_1064)
);

AOI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_1017),
.A2(n_999),
.B(n_925),
.Y(n_1065)
);

AND3x1_ASAP7_75t_SL g1066 ( 
.A(n_980),
.B(n_983),
.C(n_1028),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1006),
.B(n_1011),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_934),
.A2(n_916),
.B(n_956),
.C(n_969),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_921),
.B(n_905),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_921),
.A2(n_1035),
.B1(n_1015),
.B2(n_1011),
.Y(n_1070)
);

BUFx10_ASAP7_75t_L g1071 ( 
.A(n_1002),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1015),
.A2(n_1019),
.B1(n_939),
.B2(n_957),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_1019),
.A2(n_916),
.B(n_925),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_924),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_929),
.B(n_924),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_975),
.B(n_1013),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_957),
.B(n_941),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_982),
.B(n_959),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_961),
.B(n_1009),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_949),
.A2(n_945),
.B1(n_936),
.B2(n_942),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_926),
.A2(n_922),
.B(n_938),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_953),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_938),
.A2(n_943),
.B(n_915),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_964),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1021),
.A2(n_949),
.B(n_956),
.C(n_969),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_945),
.B(n_1018),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_984),
.B(n_1014),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_962),
.B(n_954),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_972),
.B(n_996),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_976),
.A2(n_955),
.B(n_978),
.C(n_967),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_947),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1023),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_972),
.B(n_1009),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_947),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_977),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_984),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_974),
.B(n_963),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_986),
.B(n_985),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_966),
.B(n_960),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_979),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1031),
.B(n_910),
.Y(n_1102)
);

AND2x6_ASAP7_75t_L g1103 ( 
.A(n_979),
.B(n_910),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1024),
.B(n_971),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_955),
.A2(n_923),
.B(n_927),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_967),
.A2(n_968),
.B(n_927),
.C(n_1031),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_991),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_973),
.B(n_910),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_910),
.B(n_951),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_910),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_951),
.B(n_948),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1008),
.A2(n_914),
.B1(n_951),
.B2(n_950),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1008),
.B(n_958),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_965),
.B(n_952),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_981),
.B(n_987),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_920),
.B(n_932),
.C(n_933),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_913),
.A2(n_912),
.B(n_992),
.C(n_995),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_1007),
.B(n_1012),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_1026),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1027),
.A2(n_990),
.B(n_988),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1032),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_911),
.Y(n_1122)
);

BUFx4_ASAP7_75t_SL g1123 ( 
.A(n_996),
.Y(n_1123)
);

INVx6_ASAP7_75t_L g1124 ( 
.A(n_911),
.Y(n_1124)
);

BUFx4f_ASAP7_75t_L g1125 ( 
.A(n_911),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_930),
.B(n_928),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_940),
.A2(n_989),
.B1(n_997),
.B2(n_994),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1033),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1033),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_989),
.B(n_907),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_994),
.A2(n_838),
.B(n_997),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1033),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_989),
.B(n_447),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_908),
.A2(n_614),
.B(n_449),
.Y(n_1134)
);

AO32x1_ASAP7_75t_L g1135 ( 
.A1(n_949),
.A2(n_838),
.A3(n_903),
.B1(n_830),
.B2(n_882),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_996),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1033),
.Y(n_1137)
);

NOR2x1_ASAP7_75t_SL g1138 ( 
.A(n_964),
.B(n_984),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_993),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_994),
.A2(n_838),
.B1(n_842),
.B2(n_997),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_984),
.B(n_1033),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_982),
.B(n_959),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_989),
.B(n_906),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_908),
.A2(n_614),
.B(n_449),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1033),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_987),
.A2(n_992),
.B(n_912),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_993),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_SL g1148 ( 
.A1(n_954),
.A2(n_855),
.B1(n_751),
.B2(n_665),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_930),
.B(n_928),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_931),
.B(n_930),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_935),
.B(n_1003),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_984),
.B(n_1033),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_990),
.A2(n_838),
.B(n_840),
.C(n_988),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_989),
.B(n_906),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1033),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_1002),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1033),
.Y(n_1157)
);

BUFx12f_ASAP7_75t_L g1158 ( 
.A(n_911),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_989),
.B(n_907),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1104),
.B(n_1088),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1133),
.A2(n_1127),
.B1(n_1043),
.B2(n_1140),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1123),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1039),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1104),
.B(n_1088),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1109),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1052),
.Y(n_1166)
);

BUFx4f_ASAP7_75t_SL g1167 ( 
.A(n_1158),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1111),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1136),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1041),
.A2(n_1072),
.B(n_1127),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1087),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1143),
.A2(n_1154),
.B1(n_1130),
.B2(n_1159),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1087),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1119),
.Y(n_1174)
);

CKINVDCx8_ASAP7_75t_R g1175 ( 
.A(n_1037),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_SL g1176 ( 
.A1(n_1043),
.A2(n_1064),
.B1(n_1089),
.B2(n_1083),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1075),
.B(n_1051),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1042),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1128),
.Y(n_1179)
);

INVx3_ASAP7_75t_SL g1180 ( 
.A(n_1124),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1130),
.A2(n_1159),
.B1(n_1061),
.B2(n_1062),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1058),
.B(n_1110),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1102),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1048),
.B(n_1054),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1074),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1131),
.A2(n_1053),
.B1(n_1065),
.B2(n_1073),
.Y(n_1186)
);

AO21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1131),
.A2(n_1065),
.B(n_1113),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1060),
.A2(n_1067),
.B1(n_1069),
.B2(n_1150),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1053),
.A2(n_1073),
.B1(n_1148),
.B2(n_1072),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1051),
.B(n_1055),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1129),
.Y(n_1191)
);

INVx8_ASAP7_75t_L g1192 ( 
.A(n_1080),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1114),
.A2(n_1082),
.B(n_1046),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1047),
.A2(n_1126),
.B1(n_1149),
.B2(n_1045),
.Y(n_1194)
);

AO21x1_ASAP7_75t_L g1195 ( 
.A1(n_1081),
.A2(n_1105),
.B(n_1120),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1153),
.A2(n_1081),
.B(n_1070),
.Y(n_1196)
);

AO21x1_ASAP7_75t_SL g1197 ( 
.A1(n_1120),
.A2(n_1055),
.B(n_1121),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1057),
.B(n_1069),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1070),
.A2(n_1040),
.B1(n_1076),
.B2(n_1056),
.Y(n_1199)
);

CKINVDCx6p67_ASAP7_75t_R g1200 ( 
.A(n_1071),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1106),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1103),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1044),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1077),
.B(n_1098),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1090),
.A2(n_1048),
.B1(n_1078),
.B2(n_1054),
.Y(n_1205)
);

AOI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1118),
.A2(n_1112),
.B(n_1144),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1084),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1101),
.B(n_1094),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1139),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1101),
.B(n_1086),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1084),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1118),
.A2(n_1112),
.B(n_1134),
.Y(n_1212)
);

OA21x2_ASAP7_75t_L g1213 ( 
.A1(n_1117),
.A2(n_1091),
.B(n_1116),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1048),
.A2(n_1142),
.B1(n_1078),
.B2(n_1054),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1147),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1101),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1078),
.B(n_1142),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_SL g1218 ( 
.A1(n_1142),
.A2(n_1108),
.B1(n_1157),
.B2(n_1124),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1137),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1145),
.A2(n_1155),
.B1(n_1049),
.B2(n_1132),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1135),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1125),
.A2(n_1156),
.B1(n_1071),
.B2(n_1079),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1135),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1135),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1118),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1115),
.Y(n_1226)
);

BUFx2_ASAP7_75t_R g1227 ( 
.A(n_1093),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1103),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1099),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1037),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1103),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1050),
.A2(n_1151),
.B1(n_1100),
.B2(n_1096),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1141),
.A2(n_1152),
.B1(n_1080),
.B2(n_1100),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1080),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1059),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1066),
.A2(n_1156),
.B1(n_1125),
.B2(n_1037),
.Y(n_1236)
);

INVx6_ASAP7_75t_L g1237 ( 
.A(n_1085),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1085),
.B(n_1095),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_SL g1239 ( 
.A1(n_1138),
.A2(n_1107),
.B(n_1068),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1092),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1097),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1063),
.B(n_1122),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_1122),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1074),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1074),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1133),
.A2(n_838),
.B1(n_997),
.B2(n_994),
.Y(n_1246)
);

INVxp33_ASAP7_75t_L g1247 ( 
.A(n_1132),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1042),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1133),
.B(n_1075),
.Y(n_1249)
);

OAI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_1133),
.A2(n_842),
.B(n_447),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1075),
.B(n_1017),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1123),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1146),
.A2(n_992),
.B(n_912),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1133),
.B(n_1075),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1132),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1133),
.A2(n_842),
.B1(n_1154),
.B2(n_1143),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1132),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1042),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1133),
.A2(n_838),
.B1(n_997),
.B2(n_994),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_L g1260 ( 
.A(n_1136),
.B(n_725),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1109),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1038),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1075),
.B(n_1017),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1201),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_1196),
.A2(n_1195),
.B(n_1201),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1183),
.B(n_1168),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1185),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1192),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1184),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1221),
.B(n_1223),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1244),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1224),
.A2(n_1207),
.A3(n_1211),
.B(n_1171),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1193),
.A2(n_1170),
.B(n_1206),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1165),
.Y(n_1274)
);

AO21x2_ASAP7_75t_L g1275 ( 
.A1(n_1193),
.A2(n_1170),
.B(n_1206),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1251),
.A2(n_1263),
.B1(n_1256),
.B2(n_1254),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1261),
.Y(n_1277)
);

OR2x6_ASAP7_75t_L g1278 ( 
.A(n_1184),
.B(n_1225),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1261),
.B(n_1171),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_SL g1280 ( 
.A1(n_1250),
.A2(n_1249),
.B(n_1204),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1173),
.B(n_1197),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1226),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1177),
.B(n_1190),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1226),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1244),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1212),
.A2(n_1253),
.B(n_1213),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1182),
.Y(n_1289)
);

OR2x6_ASAP7_75t_L g1290 ( 
.A(n_1184),
.B(n_1160),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1197),
.B(n_1187),
.Y(n_1291)
);

OR2x6_ASAP7_75t_L g1292 ( 
.A(n_1160),
.B(n_1164),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1182),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1187),
.B(n_1210),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1210),
.B(n_1251),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1263),
.B(n_1190),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1213),
.A2(n_1202),
.B(n_1239),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1228),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_SL g1299 ( 
.A(n_1175),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1228),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1160),
.B(n_1164),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1245),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1186),
.A2(n_1161),
.B(n_1259),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1177),
.B(n_1189),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1231),
.B(n_1163),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1231),
.A2(n_1172),
.A3(n_1262),
.B(n_1166),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1181),
.A2(n_1188),
.B(n_1236),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1245),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1217),
.Y(n_1309)
);

CKINVDCx12_ASAP7_75t_R g1310 ( 
.A(n_1208),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1217),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1255),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1246),
.B(n_1198),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1241),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1199),
.B(n_1229),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1176),
.B(n_1194),
.C(n_1218),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1296),
.B(n_1208),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1284),
.B(n_1169),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1306),
.B(n_1219),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1302),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1306),
.B(n_1272),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1296),
.B(n_1214),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1302),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1296),
.B(n_1205),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1276),
.B(n_1232),
.C(n_1222),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1295),
.B(n_1216),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1314),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1303),
.A2(n_1247),
.B(n_1220),
.Y(n_1328)
);

NOR2x1_ASAP7_75t_R g1329 ( 
.A(n_1268),
.B(n_1162),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1295),
.B(n_1216),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_L g1331 ( 
.A(n_1307),
.B(n_1280),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1290),
.B(n_1174),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1303),
.A2(n_1234),
.B1(n_1203),
.B2(n_1219),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1306),
.B(n_1257),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1284),
.B(n_1312),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1308),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1313),
.B(n_1169),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1305),
.B(n_1216),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1314),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1313),
.B(n_1215),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1305),
.B(n_1216),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1306),
.B(n_1241),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1299),
.B(n_1162),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1292),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1270),
.B(n_1240),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1270),
.B(n_1174),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1270),
.B(n_1309),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1267),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1309),
.B(n_1311),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1308),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1290),
.B(n_1174),
.Y(n_1351)
);

NAND2x1_ASAP7_75t_L g1352 ( 
.A(n_1292),
.B(n_1237),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1306),
.B(n_1209),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1311),
.B(n_1282),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1310),
.B(n_1252),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1335),
.B(n_1271),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1348),
.B(n_1271),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1331),
.B(n_1276),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1331),
.B(n_1316),
.C(n_1303),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1317),
.B(n_1287),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1325),
.A2(n_1303),
.B1(n_1316),
.B2(n_1333),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1328),
.B(n_1303),
.C(n_1265),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1333),
.B(n_1265),
.C(n_1315),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1332),
.B(n_1351),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1337),
.B(n_1200),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1354),
.B(n_1282),
.Y(n_1366)
);

OAI221xp5_ASAP7_75t_L g1367 ( 
.A1(n_1318),
.A2(n_1260),
.B1(n_1315),
.B2(n_1175),
.C(n_1180),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1336),
.B(n_1283),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1347),
.B(n_1294),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1347),
.B(n_1294),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1350),
.B(n_1283),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1320),
.B(n_1323),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1349),
.B(n_1264),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1332),
.B(n_1233),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1329),
.A2(n_1290),
.B(n_1292),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1343),
.B(n_1200),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1346),
.B(n_1264),
.Y(n_1377)
);

OAI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1340),
.A2(n_1304),
.B(n_1285),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1338),
.B(n_1291),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1327),
.Y(n_1380)
);

OAI221xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1319),
.A2(n_1304),
.B1(n_1290),
.B2(n_1292),
.C(n_1301),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1338),
.B(n_1341),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1327),
.B(n_1279),
.Y(n_1383)
);

AOI21xp33_ASAP7_75t_L g1384 ( 
.A1(n_1334),
.A2(n_1265),
.B(n_1304),
.Y(n_1384)
);

AOI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1322),
.A2(n_1286),
.B1(n_1235),
.B2(n_1298),
.C(n_1300),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1341),
.B(n_1291),
.Y(n_1386)
);

NAND4xp25_ASAP7_75t_L g1387 ( 
.A(n_1334),
.B(n_1248),
.C(n_1178),
.D(n_1179),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1326),
.B(n_1265),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1324),
.A2(n_1281),
.B1(n_1269),
.B2(n_1265),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1339),
.B(n_1279),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1355),
.A2(n_1269),
.B(n_1281),
.Y(n_1391)
);

OAI221xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1319),
.A2(n_1290),
.B1(n_1292),
.B2(n_1301),
.C(n_1278),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1326),
.B(n_1272),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1330),
.B(n_1272),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1321),
.A2(n_1288),
.B(n_1297),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1342),
.B(n_1289),
.C(n_1293),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1342),
.A2(n_1274),
.B1(n_1277),
.B2(n_1266),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1380),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1395),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1393),
.B(n_1394),
.Y(n_1400)
);

OR2x6_ASAP7_75t_SL g1401 ( 
.A(n_1363),
.B(n_1321),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1364),
.B(n_1344),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1395),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1368),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1388),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1371),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1363),
.B(n_1353),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1372),
.B(n_1353),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1393),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1394),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1366),
.B(n_1369),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1383),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1395),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1370),
.B(n_1382),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1370),
.B(n_1273),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1382),
.B(n_1273),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1390),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1395),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1373),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1377),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1397),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1374),
.B(n_1332),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1358),
.B(n_1332),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1379),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1386),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_1345),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1359),
.A2(n_1290),
.B1(n_1301),
.B2(n_1292),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1397),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1396),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1427),
.B(n_1386),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1422),
.Y(n_1433)
);

NAND2x1_ASAP7_75t_L g1434 ( 
.A(n_1427),
.B(n_1375),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1422),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1427),
.B(n_1389),
.Y(n_1436)
);

NOR2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1427),
.B(n_1359),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1399),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1422),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1421),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1421),
.Y(n_1441)
);

NAND2xp67_ASAP7_75t_L g1442 ( 
.A(n_1416),
.B(n_1242),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1399),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1407),
.B(n_1396),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1423),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1427),
.B(n_1391),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1400),
.B(n_1391),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1399),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1400),
.B(n_1351),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1423),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1407),
.B(n_1430),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1399),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1408),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1407),
.B(n_1356),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1430),
.B(n_1378),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1430),
.B(n_1360),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1400),
.B(n_1351),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1420),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1404),
.B(n_1384),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1404),
.B(n_1384),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1408),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1403),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1408),
.B(n_1410),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1419),
.B(n_1351),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1419),
.B(n_1375),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1426),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1431),
.B(n_1352),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1444),
.A2(n_1401),
.B1(n_1361),
.B2(n_1387),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1451),
.B(n_1431),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1440),
.Y(n_1473)
);

NOR2xp67_ASAP7_75t_L g1474 ( 
.A(n_1436),
.B(n_1419),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_SL g1475 ( 
.A(n_1446),
.B(n_1329),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1451),
.B(n_1431),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1440),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1438),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1444),
.B(n_1410),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1460),
.B(n_1410),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1455),
.B(n_1406),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1441),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1456),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1447),
.B(n_1419),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1458),
.Y(n_1487)
);

OAI31xp33_ASAP7_75t_L g1488 ( 
.A1(n_1437),
.A2(n_1361),
.A3(n_1429),
.B(n_1367),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1406),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1416),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1447),
.B(n_1446),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1416),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1458),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1437),
.A2(n_1401),
.B1(n_1381),
.B2(n_1392),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1454),
.B(n_1412),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1459),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1445),
.B(n_1417),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1450),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1436),
.B(n_1466),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1459),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1438),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1443),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1450),
.Y(n_1504)
);

OAI32xp33_ASAP7_75t_L g1505 ( 
.A1(n_1468),
.A2(n_1401),
.A3(n_1429),
.B1(n_1409),
.B2(n_1428),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1460),
.B(n_1362),
.C(n_1385),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1462),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1461),
.B(n_1417),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1461),
.B(n_1409),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1462),
.B(n_1405),
.Y(n_1510)
);

NAND2xp33_ASAP7_75t_SL g1511 ( 
.A(n_1434),
.B(n_1252),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1471),
.A2(n_1466),
.B1(n_1424),
.B2(n_1362),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1485),
.B(n_1449),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1469),
.B(n_1470),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1511),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1504),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1491),
.B(n_1453),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1472),
.B(n_1453),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1449),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1473),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1500),
.B(n_1457),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1472),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1500),
.B(n_1457),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1481),
.B(n_1414),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1474),
.B(n_1432),
.Y(n_1525)
);

CKINVDCx16_ASAP7_75t_R g1526 ( 
.A(n_1475),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1477),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1511),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1494),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1476),
.A2(n_1434),
.B(n_1468),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1486),
.B(n_1432),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1499),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1476),
.B(n_1464),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1468),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1482),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1508),
.B(n_1464),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1489),
.B(n_1495),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1414),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1479),
.B(n_1467),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1498),
.B(n_1414),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1483),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1479),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1486),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1510),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1487),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1493),
.B(n_1376),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1468),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1529),
.B(n_1505),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1546),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1529),
.A2(n_1546),
.B(n_1515),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1545),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1512),
.A2(n_1424),
.B1(n_1402),
.B2(n_1490),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1517),
.B(n_1465),
.Y(n_1553)
);

NAND2x1p5_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1424),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1532),
.B(n_1507),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1526),
.A2(n_1387),
.B1(n_1424),
.B2(n_1509),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1520),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_1528),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1514),
.A2(n_1488),
.B(n_1480),
.C(n_1492),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1520),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1534),
.A2(n_1480),
.B(n_1365),
.C(n_1496),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1517),
.B(n_1501),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1526),
.A2(n_1424),
.B1(n_1402),
.B2(n_1465),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1516),
.B(n_1167),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1534),
.A2(n_1275),
.B1(n_1357),
.B2(n_1415),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1518),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1522),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1522),
.B(n_1398),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1534),
.A2(n_1402),
.B1(n_1419),
.B2(n_1426),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1521),
.B(n_1411),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1567),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1548),
.A2(n_1534),
.B1(n_1543),
.B2(n_1542),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1568),
.B(n_1516),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1554),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1550),
.B(n_1516),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_R g1579 ( 
.A(n_1565),
.B(n_1243),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1563),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1558),
.B(n_1523),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1516),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1549),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1557),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1548),
.B(n_1523),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1519),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1551),
.B(n_1519),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1569),
.B(n_1562),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1555),
.B(n_1537),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1561),
.B(n_1518),
.Y(n_1591)
);

AOI32xp33_ASAP7_75t_L g1592 ( 
.A1(n_1591),
.A2(n_1559),
.A3(n_1552),
.B1(n_1566),
.B2(n_1570),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1591),
.A2(n_1566),
.B1(n_1572),
.B2(n_1565),
.C(n_1544),
.Y(n_1593)
);

OAI211xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1574),
.A2(n_1556),
.B(n_1564),
.C(n_1527),
.Y(n_1594)
);

AOI222xp33_ASAP7_75t_L g1595 ( 
.A1(n_1578),
.A2(n_1547),
.B1(n_1541),
.B2(n_1535),
.C1(n_1544),
.C2(n_1525),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1575),
.B(n_1530),
.C(n_1535),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1581),
.A2(n_1534),
.B1(n_1525),
.B2(n_1547),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_SL g1598 ( 
.A(n_1579),
.B(n_1533),
.C(n_1536),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1583),
.A2(n_1541),
.B(n_1513),
.Y(n_1599)
);

AOI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1573),
.A2(n_1533),
.B1(n_1571),
.B2(n_1536),
.C(n_1531),
.Y(n_1600)
);

AOI221x1_ASAP7_75t_L g1601 ( 
.A1(n_1582),
.A2(n_1538),
.B1(n_1540),
.B2(n_1524),
.C(n_1531),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1585),
.A2(n_1530),
.B1(n_1402),
.B2(n_1539),
.Y(n_1602)
);

AOI222xp33_ASAP7_75t_L g1603 ( 
.A1(n_1590),
.A2(n_1398),
.B1(n_1403),
.B2(n_1413),
.C1(n_1418),
.C2(n_1503),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_SL g1604 ( 
.A(n_1593),
.B(n_1579),
.C(n_1577),
.Y(n_1604)
);

NAND4xp25_ASAP7_75t_L g1605 ( 
.A(n_1598),
.B(n_1587),
.C(n_1589),
.D(n_1580),
.Y(n_1605)
);

NAND3xp33_ASAP7_75t_L g1606 ( 
.A(n_1592),
.B(n_1580),
.C(n_1576),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_L g1607 ( 
.A(n_1594),
.B(n_1576),
.Y(n_1607)
);

AND4x1_ASAP7_75t_L g1608 ( 
.A(n_1595),
.B(n_1588),
.C(n_1584),
.D(n_1586),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_L g1609 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1596),
.B(n_1586),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1597),
.B(n_1539),
.C(n_1484),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1602),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1600),
.Y(n_1613)
);

OAI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1607),
.A2(n_1603),
.B(n_1601),
.C(n_1178),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1604),
.A2(n_1484),
.B1(n_1503),
.B2(n_1502),
.C(n_1478),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1609),
.Y(n_1616)
);

NOR4xp25_ASAP7_75t_L g1617 ( 
.A(n_1606),
.B(n_1478),
.C(n_1502),
.D(n_1191),
.Y(n_1617)
);

OAI211xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1613),
.A2(n_1191),
.B(n_1510),
.C(n_1448),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1616),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1618),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1614),
.Y(n_1621)
);

NOR2x1_ASAP7_75t_L g1622 ( 
.A(n_1617),
.B(n_1605),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1615),
.Y(n_1623)
);

NOR2x1_ASAP7_75t_L g1624 ( 
.A(n_1616),
.B(n_1610),
.Y(n_1624)
);

NAND4xp75_ASAP7_75t_L g1625 ( 
.A(n_1624),
.B(n_1612),
.C(n_1608),
.D(n_1611),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1619),
.B(n_1467),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1621),
.B(n_1622),
.Y(n_1627)
);

NAND2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1620),
.B(n_1179),
.Y(n_1628)
);

NAND4xp75_ASAP7_75t_L g1629 ( 
.A(n_1623),
.B(n_1230),
.C(n_1180),
.D(n_1238),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1627),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1628),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1629),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1630),
.Y(n_1633)
);

XOR2xp5_ASAP7_75t_L g1634 ( 
.A(n_1633),
.B(n_1625),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1634),
.Y(n_1635)
);

AOI311xp33_ASAP7_75t_L g1636 ( 
.A1(n_1634),
.A2(n_1626),
.A3(n_1632),
.B(n_1631),
.C(n_1439),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1635),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1636),
.A2(n_1180),
.B1(n_1230),
.B2(n_1463),
.Y(n_1638)
);

AO221x1_ASAP7_75t_L g1639 ( 
.A1(n_1638),
.A2(n_1463),
.B1(n_1448),
.B2(n_1452),
.C(n_1443),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1637),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1640),
.A2(n_1258),
.B(n_1248),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1641),
.A2(n_1639),
.B1(n_1258),
.B2(n_1227),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1463),
.B1(n_1443),
.B2(n_1448),
.C(n_1452),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1643),
.A2(n_1452),
.B1(n_1433),
.B2(n_1435),
.Y(n_1644)
);


endmodule