module fake_jpeg_27613_n_260 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_241;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_25),
.CON(n_30),
.SN(n_30)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_34),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_16),
.B1(n_19),
.B2(n_23),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_56),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_59),
.B1(n_61),
.B2(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_19),
.B1(n_26),
.B2(n_16),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_21),
.B1(n_12),
.B2(n_24),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_37),
.B1(n_33),
.B2(n_29),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_12),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_72),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_47),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_38),
.B1(n_46),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_82),
.B1(n_68),
.B2(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_78),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_79),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_35),
.C(n_43),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_88),
.C(n_74),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_13),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_43),
.C(n_45),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_15),
.B(n_17),
.C(n_23),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_15),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_102),
.B(n_103),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_55),
.B1(n_58),
.B2(n_50),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_99),
.B1(n_106),
.B2(n_73),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_61),
.B1(n_45),
.B2(n_49),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_111),
.B1(n_105),
.B2(n_103),
.Y(n_133)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_59),
.B1(n_36),
.B2(n_65),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_89),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_53),
.Y(n_102)
);

NAND2x1_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_20),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_43),
.B1(n_61),
.B2(n_45),
.Y(n_106)
);

NAND5xp2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_32),
.C(n_24),
.D(n_18),
.E(n_25),
.Y(n_107)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_113),
.Y(n_128)
);

OR2x4_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_45),
.B1(n_49),
.B2(n_18),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_43),
.B1(n_51),
.B2(n_23),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_114),
.B1(n_80),
.B2(n_18),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_17),
.B1(n_15),
.B2(n_32),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_123),
.B1(n_137),
.B2(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_71),
.C(n_72),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_121),
.C(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_84),
.C(n_73),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_125),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_13),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_140),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_11),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_10),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_57),
.B1(n_20),
.B2(n_2),
.Y(n_137)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_139),
.Y(n_168)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_0),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_144),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_20),
.C(n_10),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_4),
.C(n_5),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_92),
.B(n_100),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_132),
.B1(n_141),
.B2(n_128),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_108),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_172),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_118),
.B(n_117),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_120),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_110),
.CI(n_103),
.CON(n_155),
.SN(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_163),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_90),
.B(n_102),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_161),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_102),
.B1(n_112),
.B2(n_94),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_164),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_107),
.B(n_114),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_125),
.A2(n_3),
.B(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_170),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_3),
.B(n_4),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_140),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_5),
.B(n_6),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_131),
.C(n_143),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_192),
.C(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_149),
.A2(n_116),
.B1(n_135),
.B2(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_123),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_122),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_137),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_171),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_150),
.C(n_152),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.C(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_168),
.C(n_161),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_176),
.B1(n_193),
.B2(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_169),
.C(n_148),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_155),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_207),
.B1(n_186),
.B2(n_174),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_157),
.B1(n_147),
.B2(n_170),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_183),
.B(n_173),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_220),
.B(n_221),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_189),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_212),
.Y(n_225)
);

FAx1_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_179),
.CI(n_172),
.CON(n_213),
.SN(n_213)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_218),
.B(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_178),
.C(n_191),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_208),
.C(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_202),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_199),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_157),
.B(n_188),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_229),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_198),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_209),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_205),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_220),
.B1(n_218),
.B2(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_238),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_213),
.B(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_147),
.B1(n_213),
.B2(n_154),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_166),
.B1(n_163),
.B2(n_155),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_231),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_229),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_243),
.B(n_244),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_223),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_240),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_245),
.B(n_247),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_9),
.B(n_6),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_9),
.B(n_6),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_234),
.B1(n_145),
.B2(n_8),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_145),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_5),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_254),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_258),
.A2(n_256),
.B(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_259),
.B(n_7),
.Y(n_260)
);


endmodule