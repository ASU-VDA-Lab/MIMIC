module fake_jpeg_25740_n_287 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_18),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_54),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_17),
.B1(n_16),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_58),
.B1(n_41),
.B2(n_44),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_61),
.Y(n_70)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_33),
.B1(n_41),
.B2(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_40),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_44),
.B1(n_41),
.B2(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_86),
.B1(n_48),
.B2(n_44),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_60),
.B1(n_51),
.B2(n_39),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_103),
.B1(n_71),
.B2(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_67),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_93),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_67),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_105),
.B(n_87),
.Y(n_118)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_106),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_39),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_40),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_43),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_112),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_71),
.B1(n_85),
.B2(n_79),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_52),
.B1(n_61),
.B2(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_90),
.B1(n_81),
.B2(n_48),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_19),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_119),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_123),
.B(n_124),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_79),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_96),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_70),
.B(n_56),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_72),
.B(n_86),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_130),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_43),
.B(n_81),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_81),
.C(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_134),
.B1(n_154),
.B2(n_23),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_148),
.B(n_33),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_90),
.B1(n_81),
.B2(n_44),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_147),
.B1(n_122),
.B2(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_58),
.B1(n_82),
.B2(n_80),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_82),
.B(n_22),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_108),
.B(n_130),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_66),
.B1(n_64),
.B2(n_23),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_119),
.C(n_112),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_166),
.C(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_159),
.A2(n_19),
.B1(n_50),
.B2(n_18),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_117),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_142),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_124),
.B1(n_99),
.B2(n_93),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_120),
.B1(n_23),
.B2(n_17),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_106),
.C(n_73),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_120),
.C(n_73),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_73),
.C(n_53),
.Y(n_170)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_178),
.Y(n_198)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_150),
.B(n_154),
.C(n_144),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_10),
.B(n_12),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_53),
.C(n_59),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_27),
.C(n_35),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_14),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_53),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_63),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_155),
.B1(n_19),
.B2(n_18),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_202),
.B1(n_13),
.B2(n_26),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_59),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_7),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_176),
.B1(n_180),
.B2(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_176),
.B1(n_50),
.B2(n_13),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_166),
.C(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_15),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_217),
.C(n_218),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_176),
.CI(n_178),
.CON(n_210),
.SN(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_216),
.B1(n_201),
.B2(n_16),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_25),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_50),
.B1(n_13),
.B2(n_16),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_27),
.C(n_28),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_27),
.C(n_28),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_221),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_27),
.C(n_28),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_190),
.B1(n_198),
.B2(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_228),
.B1(n_229),
.B2(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_190),
.B(n_184),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_233),
.B(n_11),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_221),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_200),
.B(n_10),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_1),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_211),
.B1(n_219),
.B2(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_241),
.B1(n_245),
.B2(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_246),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_207),
.B1(n_218),
.B2(n_212),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_212),
.C(n_215),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_248),
.C(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_205),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_12),
.B(n_7),
.Y(n_257)
);

NAND2x1_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_11),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_255),
.C(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_233),
.C(n_35),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_9),
.CI(n_8),
.CON(n_256),
.SN(n_256)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_2),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_12),
.B(n_24),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_25),
.B(n_3),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_254),
.B1(n_252),
.B2(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_2),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_256),
.C(n_257),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_268),
.B(n_3),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_24),
.B1(n_15),
.B2(n_29),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_24),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_273),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_24),
.C(n_35),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_269),
.B(n_261),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_275),
.B(n_5),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_275),
.C(n_265),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_276),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_24),
.Y(n_282)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_25),
.B(n_14),
.Y(n_283)
);

OAI321xp33_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_25),
.A3(n_14),
.B1(n_6),
.B2(n_5),
.C(n_4),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_25),
.C(n_6),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_4),
.A3(n_6),
.B1(n_14),
.B2(n_281),
.C1(n_258),
.C2(n_266),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_4),
.Y(n_287)
);


endmodule