module fake_ibex_862_n_910 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_910);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_910;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_170;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_741;
wire n_807;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_58),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_38),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_112),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_108),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_59),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_55),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_33),
.B(n_127),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_45),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_87),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_31),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_99),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_34),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_72),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_41),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_11),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_6),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_163),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_70),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_31),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_96),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_134),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_56),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_36),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_116),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_39),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_11),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_1),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_93),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_64),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_123),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_79),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_103),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_100),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_65),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_66),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_25),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_94),
.B(n_40),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_37),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_3),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_27),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_114),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_43),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_61),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_124),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_76),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_133),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_164),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_101),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_81),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_23),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_57),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_48),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_21),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_126),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_115),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_37),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_121),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_23),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_53),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_5),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_12),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_27),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_51),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_91),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_165),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_26),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_102),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_83),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_135),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_63),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_17),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_156),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_47),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_71),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_201),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_190),
.A2(n_67),
.B(n_158),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_193),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_223),
.B(n_0),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_210),
.B(n_2),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_221),
.A2(n_69),
.B(n_157),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_206),
.B(n_265),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_201),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_223),
.B(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_221),
.A2(n_73),
.B(n_154),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_244),
.B(n_44),
.Y(n_305)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_214),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_214),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_187),
.B(n_7),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_250),
.A2(n_75),
.B(n_153),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_177),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_62),
.B(n_152),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_172),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_210),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_214),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_212),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_259),
.A2(n_200),
.B1(n_220),
.B2(n_197),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_199),
.B(n_46),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_214),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_224),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_231),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_175),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_231),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_248),
.B(n_12),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_212),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_176),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_239),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_217),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_217),
.B(n_14),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_231),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_178),
.A2(n_84),
.B(n_150),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_179),
.A2(n_82),
.B(n_144),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_180),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g341 ( 
.A1(n_182),
.A2(n_80),
.B(n_141),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_184),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_186),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_243),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_269),
.B(n_271),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_204),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_207),
.B(n_18),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_251),
.B(n_18),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_207),
.B(n_213),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_278),
.B(n_19),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_191),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_243),
.Y(n_354)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_194),
.A2(n_89),
.B(n_140),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_195),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_213),
.B(n_20),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_231),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_196),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_209),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_219),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_240),
.B(n_202),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_203),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_208),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_211),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_228),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_216),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_226),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_227),
.B(n_21),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_230),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_331),
.A2(n_228),
.B1(n_204),
.B2(n_264),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_358),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_302),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_302),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_300),
.B(n_351),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_335),
.B(n_232),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_335),
.B(n_233),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_345),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_276),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_SL g392 ( 
.A(n_348),
.B(n_237),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_348),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_312),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_350),
.B(n_238),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_350),
.B(n_246),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

AND3x2_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_275),
.C(n_222),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_296),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_261),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_357),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_291),
.B(n_192),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_296),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_283),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_310),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_303),
.B(n_247),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_318),
.B(n_276),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_329),
.Y(n_419)
);

BUFx4f_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_303),
.B(n_183),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_315),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_315),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_314),
.B(n_252),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_317),
.B(n_255),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_329),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_328),
.B(n_256),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_301),
.B(n_237),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_322),
.A2(n_254),
.B1(n_253),
.B2(n_264),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_328),
.B(n_262),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_332),
.B(n_339),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_334),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_339),
.B(n_342),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g434 ( 
.A(n_326),
.B(n_258),
.C(n_229),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_323),
.B(n_185),
.Y(n_435)
);

XNOR2x2_ASAP7_75t_R g436 ( 
.A(n_321),
.B(n_22),
.Y(n_436)
);

NOR2x1p5_ASAP7_75t_L g437 ( 
.A(n_346),
.B(n_241),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_366),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

AND3x2_ASAP7_75t_L g440 ( 
.A(n_305),
.B(n_268),
.C(n_279),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_342),
.B(n_185),
.Y(n_441)
);

AO21x2_ASAP7_75t_L g442 ( 
.A1(n_293),
.A2(n_287),
.B(n_286),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_344),
.B(n_286),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_308),
.B(n_253),
.Y(n_446)
);

AO21x2_ASAP7_75t_L g447 ( 
.A1(n_299),
.A2(n_287),
.B(n_174),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_338),
.B(n_254),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_299),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_297),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_344),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_L g452 ( 
.A1(n_321),
.A2(n_280),
.B1(n_242),
.B2(n_284),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_343),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_347),
.A2(n_270),
.B1(n_263),
.B2(n_267),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_306),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_330),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_288),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g459 ( 
.A1(n_349),
.A2(n_245),
.B1(n_257),
.B2(n_270),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_349),
.B(n_170),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_288),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_356),
.B(n_173),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_306),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_356),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_294),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_306),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_294),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_304),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_368),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_370),
.B(n_181),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_306),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_295),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_304),
.Y(n_473)
);

INVx8_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_309),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_372),
.Y(n_477)
);

INVx6_ASAP7_75t_L g478 ( 
.A(n_368),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_353),
.B(n_188),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

OAI22x1_ASAP7_75t_L g481 ( 
.A1(n_429),
.A2(n_371),
.B1(n_353),
.B2(n_363),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_380),
.B1(n_446),
.B2(n_454),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_439),
.B(n_359),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_477),
.B(n_198),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_420),
.B(n_205),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_363),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_414),
.B(n_364),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_376),
.A2(n_367),
.B1(n_365),
.B2(n_364),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_441),
.B(n_367),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_381),
.B(n_290),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_290),
.Y(n_491)
);

OAI221xp5_ASAP7_75t_L g492 ( 
.A1(n_379),
.A2(n_289),
.B1(n_292),
.B2(n_298),
.C(n_311),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_407),
.B(n_289),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_391),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_421),
.B(n_340),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_438),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_384),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_406),
.A2(n_311),
.B1(n_298),
.B2(n_369),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_437),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_L g501 ( 
.A(n_435),
.B(n_304),
.C(n_316),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_412),
.B(n_410),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_225),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

OAI22xp33_ASAP7_75t_L g505 ( 
.A1(n_428),
.A2(n_369),
.B1(n_316),
.B2(n_313),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_422),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_377),
.B(n_235),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_450),
.B(n_236),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_423),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_431),
.B(n_369),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_448),
.A2(n_369),
.B1(n_313),
.B2(n_341),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_393),
.B(n_277),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_388),
.B(n_281),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_478),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_408),
.B(n_260),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_388),
.B(n_285),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_431),
.B(n_355),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_390),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_453),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_396),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_474),
.Y(n_525)
);

INVx8_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_385),
.B(n_355),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_385),
.B(n_355),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_435),
.A2(n_341),
.B(n_337),
.Y(n_531)
);

NOR3xp33_ASAP7_75t_L g532 ( 
.A(n_452),
.B(n_373),
.C(n_392),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_458),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_380),
.B(n_249),
.Y(n_534)
);

O2A1O1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_433),
.A2(n_337),
.B(n_338),
.C(n_26),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_394),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_460),
.B(n_337),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_394),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_397),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_462),
.B(n_24),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_443),
.B(n_98),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_446),
.B(n_28),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_443),
.B(n_106),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_470),
.B(n_107),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_467),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_470),
.B(n_90),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_434),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_479),
.B(n_119),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_459),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_382),
.B(n_34),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_424),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_472),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_383),
.B(n_122),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_424),
.B(n_35),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_400),
.B(n_128),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_425),
.B(n_36),
.Y(n_561)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_409),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_409),
.B(n_400),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_401),
.B(n_129),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_425),
.B(n_38),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_475),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_415),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_415),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_528),
.A2(n_473),
.B(n_449),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_555),
.B(n_427),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_495),
.B(n_403),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_403),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_532),
.A2(n_430),
.B1(n_427),
.B2(n_442),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_525),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_500),
.B(n_430),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_526),
.A2(n_473),
.B1(n_432),
.B2(n_440),
.Y(n_577)
);

NAND2x1_ASAP7_75t_L g578 ( 
.A(n_536),
.B(n_456),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_SL g579 ( 
.A(n_497),
.B(n_482),
.C(n_498),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_530),
.A2(n_442),
.B(n_447),
.Y(n_580)
);

AO21x1_ASAP7_75t_L g581 ( 
.A1(n_505),
.A2(n_480),
.B(n_476),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_483),
.B(n_447),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_526),
.A2(n_469),
.B1(n_471),
.B2(n_466),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_527),
.Y(n_585)
);

O2A1O1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_540),
.A2(n_378),
.B(n_375),
.C(n_374),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_512),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_490),
.B(n_455),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_546),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_491),
.B(n_49),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_516),
.B(n_52),
.Y(n_591)
);

AO21x1_ASAP7_75t_L g592 ( 
.A1(n_537),
.A2(n_389),
.B(n_445),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_554),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_54),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_554),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_504),
.Y(n_598)
);

AO21x1_ASAP7_75t_L g599 ( 
.A1(n_519),
.A2(n_387),
.B(n_426),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_487),
.B(n_60),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_513),
.B(n_489),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_501),
.A2(n_531),
.B(n_511),
.Y(n_602)
);

NOR2x1p5_ASAP7_75t_SL g603 ( 
.A(n_506),
.B(n_509),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_539),
.B(n_88),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_539),
.B(n_130),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_496),
.A2(n_387),
.B(n_417),
.Y(n_606)
);

O2A1O1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_553),
.A2(n_419),
.B(n_417),
.C(n_416),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_535),
.A2(n_568),
.B(n_567),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_481),
.B(n_132),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_507),
.A2(n_419),
.B(n_411),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_518),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_544),
.A2(n_553),
.B1(n_492),
.B2(n_565),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_524),
.B(n_405),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_484),
.B(n_137),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_521),
.A2(n_386),
.B(n_395),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_518),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_545),
.A2(n_559),
.B(n_561),
.C(n_547),
.Y(n_618)
);

CKINVDCx10_ASAP7_75t_R g619 ( 
.A(n_562),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_529),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_508),
.B(n_138),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_557),
.A2(n_399),
.B(n_160),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_488),
.B(n_503),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_518),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_520),
.B(n_522),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_560),
.A2(n_517),
.B(n_514),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_523),
.B(n_533),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_543),
.B(n_556),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_549),
.B(n_541),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_562),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_499),
.A2(n_510),
.B(n_534),
.C(n_550),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g633 ( 
.A(n_551),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_493),
.B(n_485),
.Y(n_634)
);

AO32x2_ASAP7_75t_L g635 ( 
.A1(n_552),
.A2(n_538),
.A3(n_542),
.B1(n_564),
.B2(n_562),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_593),
.B(n_515),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_620),
.Y(n_637)
);

OAI21xp33_ASAP7_75t_SL g638 ( 
.A1(n_595),
.A2(n_630),
.B(n_601),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_631),
.B(n_617),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_623),
.B(n_624),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_618),
.B(n_612),
.C(n_607),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_575),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_616),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_609),
.B(n_574),
.C(n_632),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_626),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_628),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_629),
.A2(n_582),
.B1(n_571),
.B2(n_583),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_579),
.B(n_633),
.C(n_573),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_603),
.A2(n_586),
.B(n_614),
.C(n_591),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_572),
.B(n_576),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_619),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_575),
.B(n_597),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_585),
.B(n_597),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_621),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_613),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_616),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_611),
.B(n_588),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_634),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_594),
.B(n_590),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_589),
.B(n_600),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_625),
.Y(n_661)
);

AO31x2_ASAP7_75t_L g662 ( 
.A1(n_577),
.A2(n_622),
.A3(n_606),
.B(n_584),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_615),
.A2(n_610),
.A3(n_605),
.B(n_604),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_635),
.B(n_578),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_570),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_570),
.B(n_596),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_587),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_570),
.B(n_451),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_570),
.B(n_596),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_612),
.A2(n_595),
.B1(n_593),
.B2(n_570),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_570),
.B(n_596),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_601),
.A2(n_574),
.B(n_502),
.C(n_632),
.Y(n_672)
);

AO31x2_ASAP7_75t_L g673 ( 
.A1(n_581),
.A2(n_599),
.A3(n_592),
.B(n_602),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_581),
.A2(n_599),
.A3(n_592),
.B(n_602),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_617),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_570),
.B(n_439),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_570),
.B(n_596),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_570),
.B(n_596),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_598),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_570),
.B(n_439),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_439),
.Y(n_681)
);

NOR2x1_ASAP7_75t_R g682 ( 
.A(n_617),
.B(n_438),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_570),
.B(n_446),
.Y(n_683)
);

NOR2x1_ASAP7_75t_SL g684 ( 
.A(n_631),
.B(n_448),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_570),
.B(n_451),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_R g686 ( 
.A(n_617),
.B(n_345),
.Y(n_686)
);

NOR2x1_ASAP7_75t_R g687 ( 
.A(n_617),
.B(n_438),
.Y(n_687)
);

OAI21x1_ASAP7_75t_SL g688 ( 
.A1(n_607),
.A2(n_627),
.B(n_608),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_612),
.A2(n_595),
.B1(n_593),
.B2(n_570),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_612),
.A2(n_595),
.B1(n_593),
.B2(n_570),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_587),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_569),
.A2(n_530),
.B(n_528),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_569),
.A2(n_530),
.B(n_528),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_623),
.A2(n_540),
.B(n_553),
.C(n_601),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_598),
.Y(n_695)
);

NOR4xp25_ASAP7_75t_L g696 ( 
.A(n_579),
.B(n_553),
.C(n_607),
.D(n_301),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_601),
.A2(n_574),
.B(n_502),
.C(n_632),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_581),
.A2(n_599),
.A3(n_592),
.B(n_602),
.Y(n_698)
);

BUFx4_ASAP7_75t_SL g699 ( 
.A(n_617),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_570),
.B(n_596),
.Y(n_700)
);

OAI22x1_ASAP7_75t_L g701 ( 
.A1(n_570),
.A2(n_429),
.B1(n_540),
.B2(n_321),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_617),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_598),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_570),
.B(n_446),
.Y(n_704)
);

BUFx8_ASAP7_75t_L g705 ( 
.A(n_587),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_570),
.B(n_596),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_601),
.A2(n_574),
.B(n_502),
.C(n_632),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_570),
.B(n_439),
.Y(n_708)
);

AO31x2_ASAP7_75t_L g709 ( 
.A1(n_581),
.A2(n_599),
.A3(n_592),
.B(n_602),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g710 ( 
.A1(n_602),
.A2(n_581),
.B(n_580),
.Y(n_710)
);

AO32x2_ASAP7_75t_L g711 ( 
.A1(n_577),
.A2(n_553),
.A3(n_499),
.B1(n_468),
.B2(n_581),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_570),
.B(n_596),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_570),
.B(n_596),
.Y(n_713)
);

AO31x2_ASAP7_75t_L g714 ( 
.A1(n_581),
.A2(n_599),
.A3(n_592),
.B(n_602),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_570),
.B(n_596),
.Y(n_715)
);

AO31x2_ASAP7_75t_L g716 ( 
.A1(n_581),
.A2(n_599),
.A3(n_592),
.B(n_602),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_705),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_645),
.B(n_646),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_637),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_701),
.A2(n_648),
.B1(n_654),
.B2(n_641),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_666),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_669),
.B(n_671),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_SL g723 ( 
.A1(n_647),
.A2(n_684),
.B(n_649),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_SL g724 ( 
.A1(n_672),
.A2(n_707),
.B(n_697),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_657),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_677),
.B(n_678),
.Y(n_726)
);

NAND2x1p5_ASAP7_75t_L g727 ( 
.A(n_656),
.B(n_639),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_688),
.A2(n_644),
.B(n_710),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_680),
.B(n_681),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_642),
.Y(n_730)
);

AO21x2_ASAP7_75t_L g731 ( 
.A1(n_692),
.A2(n_693),
.B(n_664),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_643),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_638),
.A2(n_640),
.B(n_694),
.Y(n_733)
);

NOR2x1_ASAP7_75t_R g734 ( 
.A(n_651),
.B(n_702),
.Y(n_734)
);

CKINVDCx14_ASAP7_75t_R g735 ( 
.A(n_665),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_708),
.A2(n_683),
.B1(n_704),
.B2(n_700),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_705),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_661),
.Y(n_738)
);

AO21x2_ASAP7_75t_L g739 ( 
.A1(n_696),
.A2(n_660),
.B(n_659),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_667),
.Y(n_740)
);

OA21x2_ASAP7_75t_L g741 ( 
.A1(n_673),
.A2(n_716),
.B(n_698),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_706),
.B(n_715),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_652),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_679),
.B(n_703),
.Y(n_744)
);

BUFx12f_ASAP7_75t_L g745 ( 
.A(n_691),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_712),
.B(n_713),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_673),
.A2(n_674),
.B(n_714),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_670),
.A2(n_690),
.B(n_689),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_658),
.A2(n_650),
.B(n_695),
.Y(n_749)
);

OA21x2_ASAP7_75t_L g750 ( 
.A1(n_673),
.A2(n_716),
.B(n_709),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_653),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_676),
.B(n_685),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_655),
.B(n_668),
.Y(n_753)
);

BUFx2_ASAP7_75t_R g754 ( 
.A(n_675),
.Y(n_754)
);

INVx6_ASAP7_75t_L g755 ( 
.A(n_636),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_711),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_636),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_663),
.A2(n_662),
.B(n_686),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_682),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_687),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_665),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_641),
.A2(n_697),
.B(n_672),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_637),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_699),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_665),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_641),
.A2(n_697),
.B(n_672),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_683),
.B(n_704),
.Y(n_768)
);

NOR2x1_ASAP7_75t_SL g769 ( 
.A(n_645),
.B(n_646),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_651),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_656),
.B(n_654),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_665),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_746),
.B(n_735),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_723),
.B(n_755),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_758),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_719),
.B(n_764),
.Y(n_776)
);

INVx3_ASAP7_75t_SL g777 ( 
.A(n_765),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_735),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_730),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_725),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_SL g781 ( 
.A(n_758),
.B(n_765),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_725),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_732),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_732),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_718),
.B(n_739),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_739),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_718),
.B(n_742),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_763),
.B(n_767),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_731),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_756),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_751),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_762),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_738),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_744),
.B(n_749),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_780),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_785),
.B(n_759),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_788),
.B(n_748),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_785),
.B(n_757),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_776),
.B(n_741),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_790),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_788),
.B(n_795),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_774),
.B(n_728),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_779),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_792),
.A2(n_720),
.B1(n_733),
.B2(n_736),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_795),
.B(n_750),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_782),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_774),
.B(n_724),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_779),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_783),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_776),
.B(n_747),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_787),
.B(n_747),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_783),
.B(n_750),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_775),
.A2(n_727),
.B1(n_761),
.B2(n_766),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_784),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_787),
.B(n_741),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_810),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_812),
.B(n_789),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_801),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_801),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_812),
.B(n_789),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_802),
.B(n_784),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_810),
.Y(n_823)
);

INVx3_ASAP7_75t_R g824 ( 
.A(n_804),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_802),
.B(n_792),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_816),
.B(n_791),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_816),
.B(n_800),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_803),
.B(n_797),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_809),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_827),
.B(n_797),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_827),
.B(n_806),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_818),
.B(n_800),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_825),
.B(n_806),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_822),
.B(n_815),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_819),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_819),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_818),
.B(n_811),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_821),
.B(n_813),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_817),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_826),
.B(n_799),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_820),
.B(n_796),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_829),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_826),
.B(n_799),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_828),
.B(n_799),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_834),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_839),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_842),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_830),
.B(n_828),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_835),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_830),
.B(n_828),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_836),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_831),
.B(n_823),
.Y(n_852)
);

OAI211xp5_ASAP7_75t_L g853 ( 
.A1(n_841),
.A2(n_720),
.B(n_778),
.C(n_773),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_833),
.B(n_815),
.Y(n_854)
);

NAND2x1_ASAP7_75t_SL g855 ( 
.A(n_844),
.B(n_777),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_833),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_831),
.B(n_838),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_857),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_SL g859 ( 
.A1(n_847),
.A2(n_775),
.B1(n_717),
.B2(n_737),
.Y(n_859)
);

CKINVDCx14_ASAP7_75t_R g860 ( 
.A(n_857),
.Y(n_860)
);

AOI222xp33_ASAP7_75t_L g861 ( 
.A1(n_846),
.A2(n_853),
.B1(n_845),
.B2(n_805),
.C1(n_856),
.C2(n_854),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_852),
.B(n_838),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_855),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_852),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_848),
.A2(n_844),
.B1(n_828),
.B2(n_840),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_848),
.A2(n_843),
.B1(n_840),
.B2(n_837),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_851),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_849),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_850),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_860),
.A2(n_814),
.B(n_850),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_860),
.A2(n_805),
.B1(n_843),
.B2(n_808),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_859),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_862),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_861),
.B(n_832),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_SL g875 ( 
.A1(n_863),
.A2(n_793),
.B(n_824),
.C(n_760),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_873),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_875),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_872),
.A2(n_865),
.B(n_866),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_874),
.A2(n_858),
.B1(n_864),
.B2(n_867),
.Y(n_879)
);

AOI222xp33_ASAP7_75t_L g880 ( 
.A1(n_871),
.A2(n_864),
.B1(n_868),
.B2(n_869),
.C1(n_781),
.C2(n_772),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_870),
.B(n_832),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_874),
.B(n_786),
.C(n_794),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_877),
.B(n_882),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_878),
.A2(n_734),
.B(n_769),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_879),
.B(n_876),
.Y(n_885)
);

AOI211xp5_ASAP7_75t_L g886 ( 
.A1(n_881),
.A2(n_777),
.B(n_880),
.C(n_807),
.Y(n_886)
);

AND3x1_ASAP7_75t_L g887 ( 
.A(n_877),
.B(n_777),
.C(n_770),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_882),
.B(n_740),
.C(n_786),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_883),
.B(n_885),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_886),
.B(n_746),
.C(n_752),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_753),
.C(n_729),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_884),
.B(n_726),
.C(n_722),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_887),
.B(n_743),
.Y(n_893)
);

NOR3xp33_ASAP7_75t_L g894 ( 
.A(n_889),
.B(n_892),
.C(n_891),
.Y(n_894)
);

NAND4xp75_ASAP7_75t_L g895 ( 
.A(n_893),
.B(n_754),
.C(n_770),
.D(n_768),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_890),
.Y(n_896)
);

AO221x1_ASAP7_75t_L g897 ( 
.A1(n_893),
.A2(n_829),
.B1(n_804),
.B2(n_824),
.C(n_721),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_889),
.A2(n_808),
.B1(n_774),
.B2(n_798),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_896),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_895),
.Y(n_900)
);

XNOR2xp5_ASAP7_75t_L g901 ( 
.A(n_900),
.B(n_894),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_899),
.Y(n_902)
);

OAI22x1_ASAP7_75t_L g903 ( 
.A1(n_901),
.A2(n_900),
.B1(n_897),
.B2(n_753),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_902),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_904),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_905),
.A2(n_903),
.B1(n_898),
.B2(n_745),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_905),
.B(n_745),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_907),
.Y(n_908)
);

AO21x2_ASAP7_75t_L g909 ( 
.A1(n_908),
.A2(n_906),
.B(n_753),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_909),
.A2(n_743),
.B1(n_730),
.B2(n_771),
.Y(n_910)
);


endmodule