module fake_jpeg_22453_n_230 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_45),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_48),
.B1(n_27),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_13),
.Y(n_63)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_36),
.B1(n_34),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_56),
.B1(n_51),
.B2(n_23),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_64),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_44),
.C(n_50),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_13),
.C(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_18),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_35),
.B1(n_14),
.B2(n_0),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_46),
.B(n_42),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_68),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_43),
.B1(n_42),
.B2(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_67),
.B1(n_66),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_52),
.B1(n_51),
.B2(n_54),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_85),
.B1(n_93),
.B2(n_73),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_63),
.B(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_89),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_73),
.B1(n_72),
.B2(n_65),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_110),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_104),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_58),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_76),
.C(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_62),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_72),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_90),
.B(n_77),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_120),
.B1(n_7),
.B2(n_1),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_121),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_128),
.C(n_135),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_76),
.B1(n_86),
.B2(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_81),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_129),
.B(n_112),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_93),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_90),
.B(n_77),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_101),
.B(n_17),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_60),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_112),
.C(n_97),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_141),
.B(n_152),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_106),
.B1(n_103),
.B2(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_102),
.B1(n_115),
.B2(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_147),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_110),
.B(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_110),
.B1(n_107),
.B2(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_107),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_101),
.C(n_94),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_149),
.C(n_151),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_101),
.C(n_60),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_14),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_126),
.B(n_130),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_151),
.Y(n_182)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_125),
.B(n_122),
.C(n_133),
.D(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_168),
.C(n_169),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_122),
.C(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_144),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_131),
.C(n_134),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_132),
.C(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_142),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_148),
.C(n_149),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_182),
.C(n_163),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_181),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_153),
.B1(n_125),
.B2(n_118),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_117),
.B1(n_174),
.B2(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_162),
.B1(n_138),
.B2(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_169),
.B1(n_164),
.B2(n_120),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_189),
.A2(n_196),
.B(n_0),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_192),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_158),
.B(n_136),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_3),
.B(n_4),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_8),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_178),
.C(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_198),
.C(n_201),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_158),
.B(n_156),
.C(n_182),
.D(n_146),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_3),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_194),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_186),
.C(n_198),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_6),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_197),
.C(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_217),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_208),
.B1(n_185),
.B2(n_5),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_6),
.B(n_9),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_215),
.C(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_213),
.B(n_219),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_6),
.B(n_9),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_225),
.C(n_11),
.Y(n_228)
);

AOI32xp33_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_12),
.Y(n_230)
);


endmodule