module real_aes_17049_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_0), .A2(n_59), .B1(n_637), .B2(n_971), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_0), .A2(n_260), .B1(n_434), .B2(n_488), .Y(n_982) );
INVx1_ASAP7_75t_L g383 ( .A(n_1), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_1), .A2(n_91), .B1(n_431), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g978 ( .A(n_2), .Y(n_978) );
XNOR2x2_ASAP7_75t_L g848 ( .A(n_3), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g296 ( .A(n_4), .Y(n_296) );
AND2x2_ASAP7_75t_L g334 ( .A(n_4), .B(n_237), .Y(n_334) );
AND2x2_ASAP7_75t_L g418 ( .A(n_4), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_4), .B(n_306), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_5), .A2(n_152), .B1(n_518), .B2(n_968), .C(n_973), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_5), .A2(n_49), .B1(n_434), .B2(n_565), .Y(n_984) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_6), .A2(n_195), .B1(n_385), .B2(n_387), .Y(n_551) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_6), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_7), .A2(n_34), .B1(n_866), .B2(n_871), .Y(n_865) );
INVx1_ASAP7_75t_L g890 ( .A(n_7), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_8), .A2(n_62), .B1(n_434), .B2(n_462), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_8), .A2(n_141), .B1(n_366), .B2(n_385), .Y(n_635) );
INVx1_ASAP7_75t_L g912 ( .A(n_9), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_9), .A2(n_165), .B1(n_494), .B2(n_892), .C(n_931), .Y(n_930) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_10), .B(n_1214), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_10), .B(n_93), .Y(n_1216) );
INVx2_ASAP7_75t_L g1220 ( .A(n_10), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_11), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_12), .A2(n_254), .B1(n_545), .B2(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g577 ( .A(n_12), .Y(n_577) );
XNOR2xp5_ASAP7_75t_L g478 ( .A(n_13), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g440 ( .A(n_14), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_15), .A2(n_60), .B1(n_385), .B2(n_387), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_15), .A2(n_277), .B1(n_422), .B2(n_425), .C(n_428), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g1231 ( .A1(n_16), .A2(n_182), .B1(n_1215), .B2(n_1221), .Y(n_1231) );
INVx1_ASAP7_75t_L g1173 ( .A(n_17), .Y(n_1173) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_17), .A2(n_181), .B1(n_1040), .B2(n_1191), .Y(n_1190) );
OAI221xp5_ASAP7_75t_L g1179 ( .A1(n_18), .A2(n_43), .B1(n_444), .B2(n_1180), .C(n_1181), .Y(n_1179) );
INVx1_ASAP7_75t_L g1201 ( .A(n_18), .Y(n_1201) );
INVx1_ASAP7_75t_L g437 ( .A(n_19), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_20), .A2(n_162), .B1(n_806), .B2(n_808), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_20), .A2(n_235), .B1(n_501), .B2(n_834), .C(n_837), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_21), .A2(n_212), .B1(n_1211), .B2(n_1218), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_22), .A2(n_277), .B1(n_385), .B2(n_387), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_22), .A2(n_60), .B1(n_462), .B2(n_464), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_23), .A2(n_269), .B1(n_1113), .B2(n_1117), .Y(n_1112) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_23), .A2(n_269), .B1(n_1152), .B2(n_1155), .Y(n_1151) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_24), .A2(n_164), .B1(n_385), .B2(n_702), .Y(n_856) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_24), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_25), .A2(n_79), .B1(n_702), .B2(n_917), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_25), .A2(n_172), .B1(n_428), .B2(n_834), .C(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g823 ( .A(n_26), .Y(n_823) );
INVx1_ASAP7_75t_L g596 ( .A(n_27), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g1238 ( .A1(n_28), .A2(n_216), .B1(n_1211), .B2(n_1221), .Y(n_1238) );
AOI22xp5_ASAP7_75t_L g1254 ( .A1(n_29), .A2(n_103), .B1(n_1211), .B2(n_1218), .Y(n_1254) );
XOR2x2_ASAP7_75t_L g989 ( .A(n_30), .B(n_990), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_31), .A2(n_86), .B1(n_1211), .B2(n_1218), .Y(n_1230) );
INVx1_ASAP7_75t_L g740 ( .A(n_32), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_33), .A2(n_422), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g511 ( .A(n_33), .Y(n_511) );
INVx1_ASAP7_75t_L g887 ( .A(n_34), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_35), .A2(n_235), .B1(n_806), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_35), .A2(n_162), .B1(n_488), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g323 ( .A(n_36), .Y(n_323) );
INVx1_ASAP7_75t_L g357 ( .A(n_36), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_37), .A2(n_133), .B1(n_422), .B2(n_612), .C(n_615), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_37), .A2(n_205), .B1(n_476), .B2(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g338 ( .A(n_38), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_39), .A2(n_210), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g512 ( .A(n_39), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_40), .A2(n_128), .B1(n_385), .B2(n_702), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_40), .A2(n_57), .B1(n_428), .B2(n_827), .C(n_828), .Y(n_826) );
INVxp67_ASAP7_75t_SL g1164 ( .A(n_41), .Y(n_1164) );
AND4x1_ASAP7_75t_L g1204 ( .A(n_41), .B(n_1166), .C(n_1169), .D(n_1188), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_42), .A2(n_65), .B1(n_1482), .B2(n_1485), .Y(n_1484) );
AOI221xp5_ASAP7_75t_L g1489 ( .A1(n_42), .A2(n_256), .B1(n_940), .B2(n_1001), .C(n_1186), .Y(n_1489) );
INVx1_ASAP7_75t_L g1203 ( .A(n_43), .Y(n_1203) );
INVx1_ASAP7_75t_L g289 ( .A(n_44), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_45), .A2(n_242), .B1(n_428), .B2(n_484), .C(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_45), .A2(n_276), .B1(n_366), .B2(n_385), .Y(n_513) );
INVx2_ASAP7_75t_L g329 ( .A(n_46), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_47), .A2(n_70), .B1(n_1218), .B2(n_1225), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_48), .A2(n_230), .B1(n_810), .B2(n_1435), .Y(n_1434) );
AOI221xp5_ASAP7_75t_L g1450 ( .A1(n_48), .A2(n_168), .B1(n_484), .B2(n_501), .C(n_1451), .Y(n_1450) );
AOI221xp5_ASAP7_75t_L g967 ( .A1(n_49), .A2(n_56), .B1(n_804), .B2(n_968), .C(n_969), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_50), .A2(n_123), .B1(n_997), .B2(n_999), .C(n_1001), .Y(n_996) );
INVx1_ASAP7_75t_L g1039 ( .A(n_50), .Y(n_1039) );
INVx1_ASAP7_75t_L g534 ( .A(n_51), .Y(n_534) );
OAI222xp33_ASAP7_75t_L g571 ( .A1(n_51), .A2(n_251), .B1(n_448), .B2(n_494), .C1(n_572), .C2(n_579), .Y(n_571) );
INVx1_ASAP7_75t_L g961 ( .A(n_52), .Y(n_961) );
INVx1_ASAP7_75t_L g960 ( .A(n_53), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_54), .A2(n_145), .B1(n_637), .B2(n_1480), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_54), .A2(n_146), .B1(n_1491), .B2(n_1493), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_55), .A2(n_136), .B1(n_488), .B2(n_882), .Y(n_1005) );
INVx1_ASAP7_75t_L g1026 ( .A(n_55), .Y(n_1026) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_56), .A2(n_152), .B1(n_425), .B2(n_563), .C(n_622), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_57), .A2(n_229), .B1(n_385), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g1440 ( .A1(n_58), .A2(n_114), .B1(n_473), .B2(n_804), .Y(n_1440) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_58), .A2(n_148), .B1(n_434), .B2(n_462), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_59), .A2(n_67), .B1(n_459), .B2(n_484), .C(n_622), .Y(n_985) );
INVx1_ASAP7_75t_L g595 ( .A(n_61), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_62), .A2(n_272), .B1(n_385), .B2(n_640), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_63), .A2(n_127), .B1(n_1211), .B2(n_1218), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_64), .Y(n_1426) );
INVx1_ASAP7_75t_L g1508 ( .A(n_65), .Y(n_1508) );
INVx1_ASAP7_75t_L g766 ( .A(n_66), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_66), .A2(n_130), .B1(n_422), .B2(n_484), .C(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_SL g970 ( .A1(n_67), .A2(n_260), .B1(n_637), .B2(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_68), .A2(n_184), .B1(n_706), .B2(n_810), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_68), .A2(n_76), .B1(n_944), .B2(n_945), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_69), .A2(n_217), .B1(n_351), .B2(n_842), .Y(n_1168) );
OAI211xp5_ASAP7_75t_L g1170 ( .A1(n_69), .A2(n_878), .B(n_1171), .C(n_1174), .Y(n_1170) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_71), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_72), .Y(n_1445) );
INVx1_ASAP7_75t_L g1475 ( .A(n_73), .Y(n_1475) );
OAI211xp5_ASAP7_75t_L g1487 ( .A1(n_73), .A2(n_413), .B(n_1488), .C(n_1495), .Y(n_1487) );
INVx1_ASAP7_75t_L g1008 ( .A(n_74), .Y(n_1008) );
INVx1_ASAP7_75t_L g797 ( .A(n_75), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_76), .A2(n_97), .B1(n_810), .B2(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g536 ( .A(n_77), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g1431 ( .A(n_78), .Y(n_1431) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_79), .Y(n_938) );
AOI22xp5_ASAP7_75t_L g1243 ( .A1(n_80), .A2(n_126), .B1(n_1211), .B2(n_1218), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_81), .A2(n_134), .B1(n_351), .B2(n_842), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_82), .A2(n_273), .B1(n_464), .B2(n_1178), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_82), .A2(n_108), .B1(n_810), .B2(n_1196), .Y(n_1197) );
AOI22xp5_ASAP7_75t_SL g1242 ( .A1(n_83), .A2(n_266), .B1(n_1221), .B2(n_1225), .Y(n_1242) );
INVx1_ASAP7_75t_L g675 ( .A(n_84), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_84), .A2(n_225), .B1(n_518), .B2(n_704), .C(n_707), .Y(n_703) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_85), .Y(n_291) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_85), .B(n_289), .Y(n_1212) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_87), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_88), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_89), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_90), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_91), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_92), .A2(n_129), .B1(n_637), .B2(n_858), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_92), .A2(n_180), .B1(n_459), .B2(n_899), .C(n_903), .Y(n_898) );
INVx1_ASAP7_75t_L g1214 ( .A(n_93), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_93), .B(n_1220), .Y(n_1222) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_94), .A2(n_240), .B1(n_730), .B2(n_733), .Y(n_729) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_94), .Y(n_737) );
INVxp67_ASAP7_75t_SL g1184 ( .A(n_95), .Y(n_1184) );
AOI22xp33_ASAP7_75t_SL g1199 ( .A1(n_95), .A2(n_218), .B1(n_543), .B2(n_709), .Y(n_1199) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_96), .A2(n_107), .B1(n_1215), .B2(n_1221), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_97), .A2(n_184), .B1(n_459), .B2(n_884), .C(n_940), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g924 ( .A1(n_98), .A2(n_176), .B1(n_866), .B2(n_871), .Y(n_924) );
INVx1_ASAP7_75t_L g951 ( .A(n_98), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_99), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_100), .A2(n_274), .B1(n_1211), .B2(n_1215), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_101), .A2(n_205), .B1(n_462), .B2(n_489), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_101), .A2(n_133), .B1(n_545), .B2(n_637), .Y(n_638) );
INVx1_ASAP7_75t_L g1011 ( .A(n_102), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g1433 ( .A1(n_104), .A2(n_148), .B1(n_804), .B2(n_915), .Y(n_1433) );
AOI221xp5_ASAP7_75t_L g1447 ( .A1(n_104), .A2(n_114), .B1(n_428), .B2(n_828), .C(n_834), .Y(n_1447) );
INVx1_ASAP7_75t_L g620 ( .A(n_105), .Y(n_620) );
INVx1_ASAP7_75t_L g627 ( .A(n_106), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_108), .A2(n_227), .B1(n_459), .B2(n_999), .C(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g378 ( .A(n_109), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_109), .A2(n_422), .B(n_459), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g1079 ( .A(n_110), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_111), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g361 ( .A(n_111), .Y(n_361) );
INVx1_ASAP7_75t_L g392 ( .A(n_111), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g1427 ( .A(n_112), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_113), .A2(n_160), .B1(n_548), .B2(n_710), .Y(n_770) );
INVx1_ASAP7_75t_L g780 ( .A(n_113), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_115), .A2(n_256), .B1(n_1480), .B2(n_1482), .Y(n_1479) );
INVx1_ASAP7_75t_L g1505 ( .A(n_115), .Y(n_1505) );
OAI22xp33_ASAP7_75t_L g1122 ( .A1(n_116), .A2(n_186), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
OAI22xp33_ASAP7_75t_L g1130 ( .A1(n_116), .A2(n_186), .B1(n_1131), .B2(n_1134), .Y(n_1130) );
AOI22xp5_ASAP7_75t_L g1226 ( .A1(n_117), .A2(n_244), .B1(n_1211), .B2(n_1218), .Y(n_1226) );
INVx1_ASAP7_75t_L g854 ( .A(n_118), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_118), .A2(n_203), .B1(n_444), .B2(n_892), .C(n_893), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g1496 ( .A(n_119), .Y(n_1496) );
INVx1_ASAP7_75t_L g686 ( .A(n_120), .Y(n_686) );
INVx1_ASAP7_75t_L g568 ( .A(n_121), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_122), .A2(n_155), .B1(n_649), .B2(n_652), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_122), .A2(n_215), .B1(n_637), .B2(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g1027 ( .A(n_123), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1046 ( .A(n_124), .B(n_317), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_125), .A2(n_238), .B1(n_340), .B2(n_351), .Y(n_339) );
OAI211xp5_ASAP7_75t_L g412 ( .A1(n_125), .A2(n_413), .B(n_420), .C(n_436), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_128), .A2(n_229), .B1(n_462), .B2(n_830), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_129), .A2(n_183), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_130), .A2(n_255), .B1(n_367), .B2(n_760), .C(n_761), .Y(n_759) );
XNOR2xp5_ASAP7_75t_L g741 ( .A(n_131), .B(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_132), .A2(n_163), .B1(n_395), .B2(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g574 ( .A(n_132), .Y(n_574) );
OAI211xp5_ASAP7_75t_L g877 ( .A1(n_134), .A2(n_878), .B(n_879), .C(n_886), .Y(n_877) );
XOR2x2_ASAP7_75t_L g906 ( .A(n_135), .B(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g1035 ( .A(n_136), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_137), .A2(n_214), .B1(n_385), .B2(n_543), .Y(n_542) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_137), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_138), .Y(n_1065) );
OAI211xp5_ASAP7_75t_SL g1100 ( .A1(n_139), .A2(n_1095), .B(n_1101), .C(n_1104), .Y(n_1100) );
INVx1_ASAP7_75t_L g1150 ( .A(n_139), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_140), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_141), .A2(n_272), .B1(n_484), .B2(n_563), .C(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_142), .Y(n_626) );
INVx1_ASAP7_75t_L g492 ( .A(n_143), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_144), .A2(n_340), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g1501 ( .A(n_145), .Y(n_1501) );
AOI22xp33_ASAP7_75t_SL g1477 ( .A1(n_146), .A2(n_149), .B1(n_637), .B2(n_1478), .Y(n_1477) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_147), .A2(n_271), .B1(n_730), .B2(n_733), .Y(n_749) );
INVxp33_ASAP7_75t_SL g789 ( .A(n_147), .Y(n_789) );
INVx1_ASAP7_75t_L g1507 ( .A(n_149), .Y(n_1507) );
AOI22xp5_ASAP7_75t_L g1233 ( .A1(n_150), .A2(n_258), .B1(n_1221), .B2(n_1234), .Y(n_1233) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_151), .A2(n_276), .B1(n_415), .B2(n_462), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_151), .A2(n_242), .B1(n_385), .B2(n_518), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_153), .A2(n_340), .B(n_589), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_154), .Y(n_1444) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_155), .A2(n_264), .B1(n_699), .B2(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g491 ( .A(n_156), .Y(n_491) );
INVx1_ASAP7_75t_L g567 ( .A(n_157), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_158), .Y(n_1077) );
BUFx3_ASAP7_75t_L g322 ( .A(n_159), .Y(n_322) );
INVx1_ASAP7_75t_L g775 ( .A(n_160), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_161), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_163), .A2(n_254), .B1(n_434), .B2(n_565), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_164), .A2(n_248), .B1(n_563), .B2(n_827), .C(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g911 ( .A(n_165), .Y(n_911) );
INVx1_ASAP7_75t_L g756 ( .A(n_166), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_166), .A2(n_209), .B1(n_422), .B2(n_484), .C(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_167), .A2(n_168), .B1(n_476), .B2(n_1438), .Y(n_1437) );
AOI22xp33_ASAP7_75t_SL g1448 ( .A1(n_167), .A2(n_230), .B1(n_434), .B2(n_462), .Y(n_1448) );
INVx1_ASAP7_75t_L g1016 ( .A(n_169), .Y(n_1016) );
OAI21xp5_ASAP7_75t_SL g1454 ( .A1(n_170), .A2(n_842), .B(n_1455), .Y(n_1454) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_171), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_172), .A2(n_241), .B1(n_804), .B2(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g744 ( .A(n_173), .Y(n_744) );
INVx1_ASAP7_75t_L g979 ( .A(n_174), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_175), .Y(n_814) );
INVx1_ASAP7_75t_L g950 ( .A(n_176), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_177), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_178), .Y(n_1108) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_179), .A2(n_215), .B1(n_652), .B2(n_671), .C(n_673), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_179), .A2(n_220), .B1(n_385), .B2(n_554), .C(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_180), .A2(n_183), .B1(n_546), .B2(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g1172 ( .A(n_181), .Y(n_1172) );
OAI21xp5_ASAP7_75t_SL g986 ( .A1(n_185), .A2(n_340), .B(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g601 ( .A(n_187), .Y(n_601) );
INVx1_ASAP7_75t_L g764 ( .A(n_188), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_189), .Y(n_1060) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_190), .Y(n_874) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_191), .A2(n_245), .B1(n_448), .B2(n_494), .C(n_495), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_191), .A2(n_245), .B1(n_402), .B2(n_405), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g1224 ( .A1(n_192), .A2(n_279), .B1(n_1221), .B2(n_1225), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_193), .A2(n_197), .B1(n_1215), .B2(n_1221), .Y(n_1264) );
INVx1_ASAP7_75t_L g1472 ( .A(n_194), .Y(n_1472) );
OAI222xp33_ASAP7_75t_L g1499 ( .A1(n_194), .A2(n_275), .B1(n_494), .B2(n_1180), .C1(n_1500), .C2(n_1506), .Y(n_1499) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_195), .Y(n_583) );
INVx1_ASAP7_75t_L g1109 ( .A(n_196), .Y(n_1109) );
OAI211xp5_ASAP7_75t_L g1137 ( .A1(n_196), .A2(n_1138), .B(n_1140), .C(n_1142), .Y(n_1137) );
XOR2x2_ASAP7_75t_L g1051 ( .A(n_197), .B(n_1052), .Y(n_1051) );
OAI211xp5_ASAP7_75t_L g993 ( .A1(n_198), .A2(n_570), .B(n_994), .C(n_995), .Y(n_993) );
INVx1_ASAP7_75t_L g1043 ( .A(n_198), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_199), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_200), .A2(n_263), .B1(n_425), .B2(n_485), .C(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1019 ( .A(n_200), .Y(n_1019) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_201), .Y(n_1182) );
AOI22xp33_ASAP7_75t_SL g1193 ( .A1(n_201), .A2(n_226), .B1(n_917), .B2(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1013 ( .A(n_202), .Y(n_1013) );
OAI332xp33_ASAP7_75t_SL g1017 ( .A1(n_202), .A2(n_508), .A3(n_553), .B1(n_1018), .B2(n_1024), .B3(n_1030), .C1(n_1034), .C2(n_1040), .Y(n_1017) );
INVx1_ASAP7_75t_L g853 ( .A(n_203), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g1498 ( .A(n_204), .Y(n_1498) );
INVx1_ASAP7_75t_L g821 ( .A(n_206), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_207), .Y(n_927) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_208), .Y(n_302) );
AOI21xp33_ASAP7_75t_L g769 ( .A1(n_209), .A2(n_706), .B(n_707), .Y(n_769) );
INVx1_ASAP7_75t_L g516 ( .A(n_210), .Y(n_516) );
INVx1_ASAP7_75t_L g816 ( .A(n_211), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_213), .Y(n_1430) );
AOI21xp33_ASAP7_75t_L g561 ( .A1(n_214), .A2(n_562), .B(n_563), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_218), .A2(n_226), .B1(n_899), .B2(n_1001), .C(n_1176), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_219), .A2(n_598), .B1(n_599), .B2(n_642), .Y(n_597) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_219), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_220), .A2(n_225), .B1(n_656), .B2(n_657), .C(n_659), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_221), .A2(n_239), .B1(n_351), .B2(n_842), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_222), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_223), .A2(n_246), .B1(n_488), .B2(n_882), .Y(n_1002) );
INVx1_ASAP7_75t_L g1033 ( .A(n_223), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_224), .A2(n_278), .B1(n_340), .B2(n_351), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_227), .A2(n_273), .B1(n_810), .B2(n_1196), .Y(n_1195) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_228), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_228), .A2(n_233), .B1(n_722), .B2(n_724), .C(n_726), .Y(n_721) );
INVx1_ASAP7_75t_L g522 ( .A(n_231), .Y(n_522) );
OAI211xp5_ASAP7_75t_SL g750 ( .A1(n_232), .A2(n_719), .B(n_726), .C(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g785 ( .A(n_232), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_233), .A2(n_243), .B1(n_662), .B2(n_667), .C(n_668), .Y(n_661) );
INVx1_ASAP7_75t_L g1010 ( .A(n_234), .Y(n_1010) );
INVx1_ASAP7_75t_L g608 ( .A(n_236), .Y(n_608) );
BUFx3_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
INVx1_ASAP7_75t_L g419 ( .A(n_237), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_239), .A2(n_413), .B(n_942), .C(n_949), .Y(n_941) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_240), .Y(n_682) );
INVxp67_ASAP7_75t_SL g935 ( .A(n_241), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_243), .A2(n_247), .B1(n_712), .B2(n_715), .Y(n_711) );
XOR2xp5_ASAP7_75t_L g1423 ( .A(n_244), .B(n_1424), .Y(n_1423) );
AOI22xp33_ASAP7_75t_L g1459 ( .A1(n_244), .A2(n_1460), .B1(n_1465), .B2(n_1515), .Y(n_1459) );
INVx1_ASAP7_75t_L g1021 ( .A(n_246), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_247), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_248), .A2(n_262), .B1(n_385), .B2(n_862), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g1071 ( .A(n_249), .Y(n_1071) );
INVx1_ASAP7_75t_L g327 ( .A(n_250), .Y(n_327) );
INVx1_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
INVx2_ASAP7_75t_L g470 ( .A(n_250), .Y(n_470) );
INVx1_ASAP7_75t_L g532 ( .A(n_251), .Y(n_532) );
XNOR2x1_ASAP7_75t_L g957 ( .A(n_252), .B(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g610 ( .A(n_253), .Y(n_610) );
INVx1_ASAP7_75t_L g776 ( .A(n_255), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_257), .A2(n_259), .B1(n_1218), .B2(n_1221), .Y(n_1217) );
INVx1_ASAP7_75t_L g845 ( .A(n_259), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_261), .A2(n_842), .B(n_843), .Y(n_841) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_262), .Y(n_897) );
INVxp67_ASAP7_75t_SL g1031 ( .A(n_263), .Y(n_1031) );
INVx1_ASAP7_75t_L g674 ( .A(n_264), .Y(n_674) );
OAI22xp33_ASAP7_75t_SL g401 ( .A1(n_265), .A2(n_270), .B1(n_402), .B2(n_405), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_265), .A2(n_270), .B1(n_444), .B2(n_448), .C(n_453), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g313 ( .A(n_266), .B(n_314), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_267), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g1466 ( .A1(n_268), .A2(n_1467), .B1(n_1468), .B2(n_1514), .Y(n_1466) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_268), .Y(n_1514) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_271), .Y(n_747) );
INVx1_ASAP7_75t_L g1471 ( .A(n_275), .Y(n_1471) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_278), .A2(n_413), .B(n_482), .C(n_490), .Y(n_481) );
OAI21xp33_ASAP7_75t_L g1509 ( .A1(n_280), .A2(n_1510), .B(n_1511), .Y(n_1509) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_307), .B(n_1205), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx4f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_292), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g1458 ( .A(n_286), .B(n_295), .Y(n_1458) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g1464 ( .A(n_288), .B(n_291), .Y(n_1464) );
INVx1_ASAP7_75t_L g1519 ( .A(n_288), .Y(n_1519) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_291), .B(n_1519), .Y(n_1521) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g1127 ( .A(n_295), .B(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g429 ( .A(n_296), .B(n_306), .Y(n_429) );
AND2x4_ASAP7_75t_L g460 ( .A(n_296), .B(n_305), .Y(n_460) );
INVx1_ASAP7_75t_L g1123 ( .A(n_297), .Y(n_1123) );
AND2x4_ASAP7_75t_SL g1457 ( .A(n_297), .B(n_1458), .Y(n_1457) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_299), .B(n_304), .Y(n_298) );
INVxp67_ASAP7_75t_L g582 ( .A(n_299), .Y(n_582) );
OR2x6_ASAP7_75t_L g1115 ( .A(n_299), .B(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g654 ( .A(n_300), .Y(n_654) );
BUFx4f_ASAP7_75t_L g934 ( .A(n_300), .Y(n_934) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
INVx1_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
INVx2_ASAP7_75t_L g417 ( .A(n_302), .Y(n_417) );
AND2x2_ASAP7_75t_L g423 ( .A(n_302), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g427 ( .A(n_302), .B(n_303), .Y(n_427) );
NAND2x1_ASAP7_75t_L g457 ( .A(n_302), .B(n_303), .Y(n_457) );
INVx1_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
AND2x2_ASAP7_75t_L g416 ( .A(n_303), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g424 ( .A(n_303), .Y(n_424) );
BUFx2_ASAP7_75t_L g451 ( .A(n_303), .Y(n_451) );
OR2x2_ASAP7_75t_L g576 ( .A(n_303), .B(n_336), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_303), .B(n_417), .Y(n_587) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g1103 ( .A(n_305), .Y(n_1103) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g1107 ( .A(n_306), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_306), .B(n_348), .Y(n_1111) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_791), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
XNOR2x1_ASAP7_75t_L g310 ( .A(n_311), .B(n_526), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_477), .B1(n_478), .B2(n_525), .Y(n_312) );
INVx1_ASAP7_75t_L g525 ( .A(n_313), .Y(n_525) );
AND4x1_ASAP7_75t_L g314 ( .A(n_315), .B(n_363), .C(n_411), .D(n_471), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_338), .B(n_339), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_316), .A2(n_522), .B(n_523), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_316), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_316), .B(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_316), .A2(n_631), .B1(n_797), .B2(n_798), .C(n_799), .Y(n_796) );
AOI21xp33_ASAP7_75t_SL g873 ( .A1(n_316), .A2(n_874), .B(n_875), .Y(n_873) );
AOI21xp33_ASAP7_75t_SL g926 ( .A1(n_316), .A2(n_927), .B(n_928), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_316), .A2(n_631), .B1(n_960), .B2(n_961), .C(n_962), .Y(n_959) );
AOI21xp33_ASAP7_75t_L g1166 ( .A1(n_316), .A2(n_1167), .B(n_1168), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1425 ( .A1(n_316), .A2(n_631), .B1(n_1426), .B2(n_1427), .C(n_1428), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_316), .B(n_1513), .Y(n_1512) );
INVx8_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_330), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_324), .Y(n_318) );
BUFx3_ASAP7_75t_L g757 ( .A(n_319), .Y(n_757) );
INVx1_ASAP7_75t_L g1023 ( .A(n_319), .Y(n_1023) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_320), .Y(n_398) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g382 ( .A(n_321), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_322), .Y(n_345) );
INVx2_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
AND2x4_ASAP7_75t_L g367 ( .A(n_322), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g869 ( .A(n_322), .B(n_356), .Y(n_869) );
INVx1_ASAP7_75t_L g344 ( .A(n_323), .Y(n_344) );
INVx2_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
OR2x2_ASAP7_75t_L g341 ( .A(n_324), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g474 ( .A(n_324), .Y(n_474) );
INVx1_ASAP7_75t_L g593 ( .A(n_324), .Y(n_593) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
OR2x2_ASAP7_75t_L g372 ( .A(n_325), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_SL g660 ( .A(n_325), .B(n_429), .Y(n_660) );
INVx1_ASAP7_75t_L g783 ( .A(n_325), .Y(n_783) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_325), .Y(n_1161) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g350 ( .A(n_326), .Y(n_350) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g714 ( .A(n_328), .Y(n_714) );
INVx1_ASAP7_75t_L g732 ( .A(n_328), .Y(n_732) );
INVx3_ASAP7_75t_L g359 ( .A(n_329), .Y(n_359) );
NAND2xp33_ASAP7_75t_SL g373 ( .A(n_329), .B(n_361), .Y(n_373) );
BUFx3_ASAP7_75t_L g541 ( .A(n_329), .Y(n_541) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
AND2x4_ASAP7_75t_L g369 ( .A(n_331), .B(n_358), .Y(n_369) );
INVx1_ASAP7_75t_L g680 ( .A(n_331), .Y(n_680) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_332), .B(n_418), .Y(n_685) );
INVx1_ASAP7_75t_L g681 ( .A(n_333), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_334), .B(n_348), .Y(n_347) );
AND2x6_ASAP7_75t_L g435 ( .A(n_334), .B(n_426), .Y(n_435) );
INVx1_ASAP7_75t_L g452 ( .A(n_334), .Y(n_452) );
AND2x2_ASAP7_75t_L g606 ( .A(n_334), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_334), .B(n_470), .Y(n_664) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_335), .Y(n_433) );
AND2x2_ASAP7_75t_L g439 ( .A(n_335), .B(n_418), .Y(n_439) );
INVx3_ASAP7_75t_L g463 ( .A(n_335), .Y(n_463) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_346), .Y(n_340) );
AND2x4_ASAP7_75t_L g842 ( .A(n_341), .B(n_346), .Y(n_842) );
INVx3_ASAP7_75t_L g768 ( .A(n_342), .Y(n_768) );
INVx4_ASAP7_75t_L g1029 ( .A(n_342), .Y(n_1029) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g727 ( .A(n_343), .Y(n_727) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_343), .Y(n_1073) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
BUFx2_ASAP7_75t_L g1149 ( .A(n_344), .Y(n_1149) );
INVx2_ASAP7_75t_L g404 ( .A(n_345), .Y(n_404) );
AND2x4_ASAP7_75t_L g548 ( .A(n_345), .B(n_410), .Y(n_548) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_345), .Y(n_1146) );
INVx2_ASAP7_75t_SL g787 ( .A(n_346), .Y(n_787) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_350), .Y(n_346) );
OR2x2_ASAP7_75t_L g667 ( .A(n_347), .B(n_350), .Y(n_667) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVxp67_ASAP7_75t_L g362 ( .A(n_350), .Y(n_362) );
INVx1_ASAP7_75t_L g695 ( .A(n_350), .Y(n_695) );
INVx1_ASAP7_75t_L g1128 ( .A(n_350), .Y(n_1128) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_362), .Y(n_351) );
OR2x6_ASAP7_75t_L g538 ( .A(n_352), .B(n_362), .Y(n_538) );
INVx2_ASAP7_75t_L g720 ( .A(n_352), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_353), .B(n_358), .Y(n_352) );
INVx8_ASAP7_75t_L g386 ( .A(n_353), .Y(n_386) );
BUFx3_ASAP7_75t_L g710 ( .A(n_353), .Y(n_710) );
AND2x2_ASAP7_75t_L g713 ( .A(n_353), .B(n_714), .Y(n_713) );
BUFx3_ASAP7_75t_L g917 ( .A(n_353), .Y(n_917) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
AND2x4_ASAP7_75t_L g376 ( .A(n_354), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVxp67_ASAP7_75t_L g377 ( .A(n_357), .Y(n_377) );
AND2x6_ASAP7_75t_L g723 ( .A(n_358), .B(n_403), .Y(n_723) );
AND2x2_ASAP7_75t_L g725 ( .A(n_358), .B(n_409), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_358), .Y(n_728) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND3x1_ASAP7_75t_L g390 ( .A(n_359), .B(n_391), .C(n_392), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_359), .B(n_392), .Y(n_554) );
OR2x4_ASAP7_75t_L g1133 ( .A(n_359), .B(n_869), .Y(n_1133) );
INVx1_ASAP7_75t_L g1136 ( .A(n_359), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_359), .B(n_367), .Y(n_1141) );
OR2x6_ASAP7_75t_L g1156 ( .A(n_359), .B(n_382), .Y(n_1156) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND3x4_ASAP7_75t_L g540 ( .A(n_361), .B(n_505), .C(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g1159 ( .A(n_361), .Y(n_1159) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_370), .C(n_401), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_365), .B(n_507), .C(n_520), .Y(n_506) );
INVx3_ASAP7_75t_L g555 ( .A(n_365), .Y(n_555) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_365), .A2(n_620), .B(n_631), .C(n_632), .Y(n_630) );
INVx3_ASAP7_75t_L g800 ( .A(n_365), .Y(n_800) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g387 ( .A(n_367), .Y(n_387) );
INVx2_ASAP7_75t_L g519 ( .A(n_367), .Y(n_519) );
BUFx3_ASAP7_75t_L g702 ( .A(n_367), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_367), .B(n_714), .Y(n_716) );
BUFx2_ASAP7_75t_L g804 ( .A(n_367), .Y(n_804) );
BUFx2_ASAP7_75t_L g862 ( .A(n_367), .Y(n_862) );
BUFx2_ASAP7_75t_L g1194 ( .A(n_367), .Y(n_1194) );
INVx1_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
NAND2x1_ASAP7_75t_L g402 ( .A(n_369), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_SL g406 ( .A(n_369), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_SL g533 ( .A(n_369), .B(n_403), .Y(n_533) );
AND2x4_ASAP7_75t_L g817 ( .A(n_369), .B(n_407), .Y(n_817) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_369), .B(n_403), .Y(n_1202) );
OAI22xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_374), .B1(n_388), .B2(n_393), .Y(n_370) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_371), .Y(n_1055) );
BUFx4f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx8_ASAP7_75t_L g508 ( .A(n_372), .Y(n_508) );
BUFx2_ASAP7_75t_L g707 ( .A(n_373), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_379), .B2(n_383), .C(n_384), .Y(n_374) );
INVx3_ASAP7_75t_L g592 ( .A(n_375), .Y(n_592) );
INVx1_ASAP7_75t_L g699 ( .A(n_375), .Y(n_699) );
OR2x6_ASAP7_75t_SL g730 ( .A(n_375), .B(n_731), .Y(n_730) );
BUFx2_ASAP7_75t_L g920 ( .A(n_375), .Y(n_920) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_376), .Y(n_395) );
BUFx8_ASAP7_75t_L g476 ( .A(n_376), .Y(n_476) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_376), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_379), .A2(n_510), .B1(n_511), .B2(n_512), .C(n_513), .Y(n_509) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g1485 ( .A(n_385), .Y(n_1485) );
INVx8_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g473 ( .A(n_386), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_386), .Y(n_760) );
INVx2_ASAP7_75t_L g968 ( .A(n_386), .Y(n_968) );
INVx3_ASAP7_75t_L g1478 ( .A(n_386), .Y(n_1478) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_389), .Y(n_514) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g864 ( .A(n_390), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B1(n_397), .B2(n_399), .C(n_400), .Y(n_393) );
INVx1_ASAP7_75t_L g545 ( .A(n_394), .Y(n_545) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g859 ( .A(n_395), .Y(n_859) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_395), .Y(n_971) );
INVx2_ASAP7_75t_L g1064 ( .A(n_395), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_395), .B(n_1136), .Y(n_1135) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_396), .A2(n_454), .B(n_458), .C(n_461), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_397), .A2(n_496), .B1(n_510), .B2(n_516), .C(n_517), .Y(n_515) );
CKINVDCx8_ASAP7_75t_R g397 ( .A(n_398), .Y(n_397) );
INVx3_ASAP7_75t_L g1066 ( .A(n_398), .Y(n_1066) );
INVx3_ASAP7_75t_L g1078 ( .A(n_398), .Y(n_1078) );
INVx2_ASAP7_75t_L g815 ( .A(n_402), .Y(n_815) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_406), .A2(n_532), .B1(n_533), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_406), .A2(n_533), .B1(n_608), .B2(n_610), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_406), .A2(n_533), .B1(n_964), .B2(n_965), .Y(n_963) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_443), .B(n_466), .Y(n_411) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_414), .B(n_536), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g825 ( .A1(n_414), .A2(n_435), .B1(n_797), .B2(n_826), .C(n_829), .Y(n_825) );
INVx3_ASAP7_75t_L g878 ( .A(n_414), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g1446 ( .A1(n_414), .A2(n_435), .B1(n_1426), .B2(n_1447), .C(n_1448), .Y(n_1446) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
BUFx2_ASAP7_75t_L g882 ( .A(n_415), .Y(n_882) );
INVx1_ASAP7_75t_L g1494 ( .A(n_415), .Y(n_1494) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
INVx2_ASAP7_75t_L g465 ( .A(n_416), .Y(n_465) );
BUFx3_ASAP7_75t_L g489 ( .A(n_416), .Y(n_489) );
AND2x4_ASAP7_75t_L g441 ( .A(n_418), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_SL g447 ( .A(n_418), .B(n_426), .Y(n_447) );
AND2x2_ASAP7_75t_L g618 ( .A(n_418), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g739 ( .A(n_418), .B(n_442), .Y(n_739) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_419), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_430), .B(n_435), .Y(n_420) );
BUFx2_ASAP7_75t_L g828 ( .A(n_422), .Y(n_828) );
INVx1_ASAP7_75t_L g998 ( .A(n_422), .Y(n_998) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_423), .Y(n_442) );
INVx2_ASAP7_75t_L g902 ( .A(n_423), .Y(n_902) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_423), .B(n_1116), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g484 ( .A(n_426), .Y(n_484) );
BUFx3_ASAP7_75t_L g827 ( .A(n_426), .Y(n_827) );
BUFx3_ASAP7_75t_L g903 ( .A(n_426), .Y(n_903) );
BUFx3_ASAP7_75t_L g940 ( .A(n_426), .Y(n_940) );
INVx1_ASAP7_75t_L g1000 ( .A(n_426), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_426), .B(n_1103), .Y(n_1102) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g614 ( .A(n_427), .Y(n_614) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_L g563 ( .A(n_429), .Y(n_563) );
AND2x4_ASAP7_75t_L g781 ( .A(n_429), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g1001 ( .A(n_429), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_429), .B(n_782), .Y(n_1098) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g1492 ( .A(n_433), .Y(n_1492) );
BUFx3_ASAP7_75t_L g830 ( .A(n_434), .Y(n_830) );
INVx1_ASAP7_75t_SL g946 ( .A(n_434), .Y(n_946) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_435), .A2(n_483), .B(n_487), .Y(n_482) );
INVx1_ASAP7_75t_L g570 ( .A(n_435), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_435), .A2(n_618), .B1(n_620), .B2(n_621), .C(n_624), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_435), .A2(n_880), .B(n_883), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_435), .A2(n_943), .B(n_947), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_435), .A2(n_618), .B1(n_960), .B2(n_981), .C(n_982), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g1174 ( .A1(n_435), .A2(n_1175), .B(n_1177), .Y(n_1174) );
AOI21xp5_ASAP7_75t_L g1488 ( .A1(n_435), .A2(n_1489), .B(n_1490), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_437), .A2(n_440), .B1(n_472), .B2(n_475), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_438), .A2(n_441), .B1(n_567), .B2(n_568), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_438), .A2(n_441), .B1(n_626), .B2(n_627), .Y(n_625) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_438), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_438), .A2(n_441), .B1(n_978), .B2(n_979), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_438), .B(n_1013), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_438), .A2(n_824), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_438), .A2(n_824), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_439), .A2(n_441), .B1(n_491), .B2(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g694 ( .A(n_439), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g889 ( .A(n_439), .Y(n_889) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_441), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_441), .A2(n_618), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1497 ( .A(n_441), .Y(n_1497) );
INVx1_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_442), .Y(n_562) );
INVx2_ASAP7_75t_L g623 ( .A(n_442), .Y(n_623) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
INVx1_ASAP7_75t_L g994 ( .A(n_445), .Y(n_994) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g609 ( .A(n_447), .Y(n_609) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_448), .Y(n_1180) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g892 ( .A(n_449), .Y(n_892) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g607 ( .A(n_451), .Y(n_607) );
INVx1_ASAP7_75t_L g666 ( .A(n_451), .Y(n_666) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_451), .B(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g573 ( .A(n_455), .Y(n_573) );
INVx4_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx4f_ASAP7_75t_L g560 ( .A(n_456), .Y(n_560) );
BUFx4f_ASAP7_75t_L g658 ( .A(n_456), .Y(n_658) );
OR2x6_ASAP7_75t_L g668 ( .A(n_456), .B(n_669), .Y(n_668) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g499 ( .A(n_457), .Y(n_499) );
INVx1_ASAP7_75t_L g578 ( .A(n_459), .Y(n_578) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
INVx3_ASAP7_75t_L g615 ( .A(n_460), .Y(n_615) );
INVx2_ASAP7_75t_L g1007 ( .A(n_460), .Y(n_1007) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g488 ( .A(n_463), .Y(n_488) );
INVx1_ASAP7_75t_L g565 ( .A(n_463), .Y(n_565) );
INVx2_ASAP7_75t_L g881 ( .A(n_463), .Y(n_881) );
INVx1_ASAP7_75t_L g944 ( .A(n_463), .Y(n_944) );
INVx2_ASAP7_75t_L g1178 ( .A(n_463), .Y(n_1178) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g619 ( .A(n_465), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_466), .A2(n_819), .B(n_841), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g975 ( .A1(n_466), .A2(n_976), .B(n_986), .Y(n_975) );
OAI21xp5_ASAP7_75t_L g992 ( .A1(n_466), .A2(n_993), .B(n_1003), .Y(n_992) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g603 ( .A(n_467), .Y(n_603) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g1187 ( .A(n_468), .Y(n_1187) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x6_ASAP7_75t_L g553 ( .A(n_469), .B(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g676 ( .A(n_469), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g969 ( .A(n_469), .B(n_554), .Y(n_969) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g505 ( .A(n_470), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_472), .A2(n_475), .B1(n_491), .B2(n_492), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_472), .A2(n_591), .B1(n_626), .B2(n_627), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_472), .A2(n_475), .B1(n_821), .B2(n_823), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_472), .A2(n_475), .B1(n_1444), .B2(n_1445), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_472), .A2(n_475), .B1(n_1496), .B2(n_1498), .Y(n_1511) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x4_ASAP7_75t_L g590 ( .A(n_473), .B(n_474), .Y(n_590) );
AND2x4_ASAP7_75t_L g475 ( .A(n_474), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g871 ( .A(n_475), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_475), .B(n_1010), .Y(n_1045) );
INVx2_ASAP7_75t_L g1191 ( .A(n_475), .Y(n_1191) );
INVx2_ASAP7_75t_SL g510 ( .A(n_476), .Y(n_510) );
INVx2_ASAP7_75t_SL g807 ( .A(n_476), .Y(n_807) );
INVx3_ASAP7_75t_L g1020 ( .A(n_476), .Y(n_1020) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND4x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_506), .C(n_521), .D(n_524), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_493), .B(n_503), .Y(n_480) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OAI211xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_500), .C(n_502), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_497), .A2(n_1063), .B1(n_1071), .B2(n_1090), .Y(n_1089) );
INVx5_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g688 ( .A(n_499), .B(n_685), .Y(n_688) );
BUFx2_ASAP7_75t_SL g1095 ( .A(n_499), .Y(n_1095) );
O2A1O1Ixp5_ASAP7_75t_SL g556 ( .A1(n_503), .A2(n_557), .B(n_571), .C(n_588), .Y(n_556) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g735 ( .A(n_504), .Y(n_735) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI31xp33_ASAP7_75t_SL g748 ( .A1(n_505), .A2(n_749), .A3(n_750), .B(n_754), .Y(n_748) );
INVx2_ASAP7_75t_SL g904 ( .A(n_505), .Y(n_904) );
OAI22xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_509), .B1(n_514), .B2(n_515), .Y(n_507) );
INVx1_ASAP7_75t_L g811 ( .A(n_514), .Y(n_811) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g543 ( .A(n_519), .Y(n_543) );
INVx2_ASAP7_75t_L g640 ( .A(n_519), .Y(n_640) );
INVx1_ASAP7_75t_L g1482 ( .A(n_519), .Y(n_1482) );
XOR2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_643), .Y(n_526) );
XNOR2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_597), .Y(n_527) );
XOR2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_596), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_556), .C(n_594), .Y(n_529) );
AND4x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .C(n_539), .D(n_555), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_537), .B(n_1011), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_537), .B(n_1475), .Y(n_1474) );
INVx5_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g631 ( .A(n_538), .Y(n_631) );
AOI33xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .A3(n_544), .B1(n_549), .B2(n_551), .B3(n_552), .Y(n_539) );
AOI33xp33_ASAP7_75t_L g634 ( .A1(n_540), .A2(n_635), .A3(n_636), .B1(n_638), .B2(n_639), .B3(n_641), .Y(n_634) );
BUFx3_ASAP7_75t_L g802 ( .A(n_540), .Y(n_802) );
AOI33xp33_ASAP7_75t_L g855 ( .A1(n_540), .A2(n_856), .A3(n_857), .B1(n_860), .B2(n_861), .B3(n_863), .Y(n_855) );
AOI33xp33_ASAP7_75t_L g913 ( .A1(n_540), .A2(n_914), .A3(n_918), .B1(n_921), .B2(n_922), .B3(n_923), .Y(n_913) );
INVx1_ASAP7_75t_L g973 ( .A(n_540), .Y(n_973) );
AOI33xp33_ASAP7_75t_L g1192 ( .A1(n_540), .A2(n_1193), .A3(n_1195), .B1(n_1197), .B2(n_1198), .B3(n_1199), .Y(n_1192) );
INVx3_ASAP7_75t_L g1145 ( .A(n_541), .Y(n_1145) );
INVx2_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g550 ( .A(n_547), .Y(n_550) );
INVx1_ASAP7_75t_L g808 ( .A(n_547), .Y(n_808) );
INVx5_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx12f_ASAP7_75t_L g637 ( .A(n_548), .Y(n_637) );
BUFx2_ASAP7_75t_L g700 ( .A(n_548), .Y(n_700) );
AND2x4_ASAP7_75t_L g734 ( .A(n_548), .B(n_732), .Y(n_734) );
BUFx3_ASAP7_75t_L g810 ( .A(n_548), .Y(n_810) );
BUFx3_ASAP7_75t_L g1438 ( .A(n_548), .Y(n_1438) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g641 ( .A(n_553), .Y(n_641) );
INVx3_ASAP7_75t_L g762 ( .A(n_554), .Y(n_762) );
INVx1_ASAP7_75t_L g872 ( .A(n_555), .Y(n_872) );
NAND4xp25_ASAP7_75t_L g1041 ( .A(n_555), .B(n_1042), .C(n_1044), .D(n_1045), .Y(n_1041) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_558), .B(n_566), .C(n_569), .D(n_570), .Y(n_557) );
OAI211xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_561), .C(n_564), .Y(n_558) );
BUFx3_ASAP7_75t_L g948 ( .A(n_562), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_567), .A2(n_568), .B1(n_590), .B2(n_591), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_577), .C(n_578), .Y(n_572) );
INVx2_ASAP7_75t_L g656 ( .A(n_575), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_575), .A2(n_658), .B1(n_674), .B2(n_675), .C(n_676), .Y(n_673) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_576), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1504 ( .A(n_576), .Y(n_1504) );
OAI221xp5_ASAP7_75t_L g1500 ( .A1(n_578), .A2(n_1095), .B1(n_1501), .B2(n_1502), .C(n_1505), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_583), .B2(n_584), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_584), .A2(n_654), .B1(n_775), .B2(n_776), .Y(n_774) );
OAI22x1_ASAP7_75t_SL g779 ( .A1(n_584), .A2(n_654), .B1(n_758), .B2(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g651 ( .A(n_585), .Y(n_651) );
INVx2_ASAP7_75t_SL g896 ( .A(n_585), .Y(n_896) );
BUFx6f_ASAP7_75t_L g937 ( .A(n_585), .Y(n_937) );
INVx4_ASAP7_75t_L g1088 ( .A(n_585), .Y(n_1088) );
INVx8_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g672 ( .A(n_586), .Y(n_672) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_586), .B(n_1107), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_590), .A2(n_591), .B1(n_978), .B2(n_979), .Y(n_987) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVxp67_ASAP7_75t_L g870 ( .A(n_593), .Y(n_870) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .C(n_630), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_628), .Y(n_602) );
AOI21xp5_ASAP7_75t_SL g1441 ( .A1(n_603), .A2(n_1442), .B(n_1454), .Y(n_1441) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_617), .C(n_625), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B1(n_609), .B2(n_610), .C1(n_611), .C2(n_616), .Y(n_605) );
INVx1_ASAP7_75t_L g840 ( .A(n_606), .Y(n_840) );
AOI222xp33_ASAP7_75t_L g983 ( .A1(n_606), .A2(n_609), .B1(n_964), .B2(n_965), .C1(n_984), .C2(n_985), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_606), .A2(n_1005), .B1(n_1006), .B2(n_1008), .Y(n_1004) );
AOI222xp33_ASAP7_75t_L g831 ( .A1(n_609), .A2(n_814), .B1(n_816), .B2(n_832), .C1(n_833), .C2(n_839), .Y(n_831) );
AOI222xp33_ASAP7_75t_L g1449 ( .A1(n_609), .A2(n_839), .B1(n_1430), .B2(n_1431), .C1(n_1450), .C2(n_1453), .Y(n_1449) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g836 ( .A(n_614), .Y(n_836) );
AND2x4_ASAP7_75t_L g683 ( .A(n_619), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g838 ( .A(n_622), .Y(n_838) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g885 ( .A(n_623), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_741), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_740), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_696), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g646 ( .A(n_647), .B(n_678), .C(n_690), .Y(n_646) );
AOI211xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_655), .B(n_661), .C(n_670), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_650), .Y(n_1183) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g893 ( .A1(n_653), .A2(n_894), .B1(n_895), .B2(n_897), .C(n_898), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g1506 ( .A1(n_653), .A2(n_1183), .B1(n_1507), .B2(n_1508), .Y(n_1506) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_654), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g786 ( .A(n_662), .Y(n_786) );
NAND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g669 ( .A(n_663), .Y(n_669) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_668), .Y(n_790) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_676), .Y(n_777) );
INVx4_ASAP7_75t_L g1081 ( .A(n_676), .Y(n_1081) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B1(n_683), .B2(n_686), .C1(n_687), .C2(n_689), .Y(n_678) );
AOI21xp33_ASAP7_75t_SL g788 ( .A1(n_679), .A2(n_789), .B(n_790), .Y(n_788) );
AND2x4_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g784 ( .A1(n_683), .A2(n_752), .B1(n_764), .B2(n_785), .C1(n_786), .C2(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_686), .A2(n_718), .B(n_721), .C(n_729), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g772 ( .A1(n_687), .A2(n_753), .B1(n_773), .B2(n_777), .C1(n_778), .C2(n_781), .Y(n_772) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_694), .Y(n_743) );
AND2x4_ASAP7_75t_L g738 ( .A(n_695), .B(n_739), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_717), .B(n_735), .C(n_736), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B1(n_703), .B2(n_708), .C(n_711), .Y(n_697) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_705), .A2(n_756), .B1(n_757), .B2(n_758), .C(n_759), .Y(n_755) );
INVx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx5_ASAP7_75t_L g1070 ( .A(n_706), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1436 ( .A(n_706), .Y(n_1436) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_713), .A2(n_716), .B1(n_744), .B2(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx4_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_723), .A2(n_725), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OR2x6_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g1038 ( .A(n_727), .Y(n_1038) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_738), .B(n_747), .Y(n_746) );
AOI211x1_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B(n_745), .C(n_771), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_763), .C(n_765), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_757), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B(n_769), .C(n_770), .Y(n_765) );
INVx3_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g1061 ( .A(n_768), .Y(n_1061) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_784), .C(n_788), .Y(n_771) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
XOR2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_953), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_905), .B1(n_906), .B2(n_952), .Y(n_792) );
INVx1_ASAP7_75t_L g952 ( .A(n_793), .Y(n_952) );
XNOR2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_847), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_794) );
INVx1_ASAP7_75t_L g846 ( .A(n_795), .Y(n_846) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_818), .Y(n_795) );
NAND3xp33_ASAP7_75t_SL g799 ( .A(n_800), .B(n_801), .C(n_813), .Y(n_799) );
INVx2_ASAP7_75t_SL g925 ( .A(n_800), .Y(n_925) );
NAND3xp33_ASAP7_75t_SL g962 ( .A(n_800), .B(n_963), .C(n_966), .Y(n_962) );
AND4x1_ASAP7_75t_L g1188 ( .A(n_800), .B(n_1189), .C(n_1192), .D(n_1200), .Y(n_1188) );
NAND3xp33_ASAP7_75t_SL g1428 ( .A(n_800), .B(n_1429), .C(n_1432), .Y(n_1428) );
AND4x1_ASAP7_75t_L g1469 ( .A(n_800), .B(n_1470), .C(n_1474), .D(n_1476), .Y(n_1469) );
AOI33xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .A3(n_805), .B1(n_809), .B2(n_811), .B3(n_812), .Y(n_801) );
AOI33xp33_ASAP7_75t_L g1432 ( .A1(n_802), .A2(n_1433), .A3(n_1434), .B1(n_1437), .B2(n_1439), .B3(n_1440), .Y(n_1432) );
AOI33xp33_ASAP7_75t_L g1476 ( .A1(n_802), .A2(n_922), .A3(n_1477), .B1(n_1479), .B2(n_1483), .B3(n_1484), .Y(n_1476) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_815), .A2(n_817), .B1(n_853), .B2(n_854), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_815), .A2(n_817), .B1(n_911), .B2(n_912), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_815), .A2(n_817), .B1(n_1008), .B2(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_815), .A2(n_817), .B1(n_1430), .B2(n_1431), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_815), .A2(n_1471), .B1(n_1472), .B2(n_1473), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_817), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1473 ( .A(n_817), .Y(n_1473) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_825), .C(n_831), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_824), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_824), .A2(n_887), .B1(n_888), .B2(n_890), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_824), .A2(n_888), .B1(n_950), .B2(n_951), .Y(n_949) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g1015 ( .A(n_842), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1510 ( .A(n_842), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND3xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_873), .C(n_876), .Y(n_849) );
NOR3xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_865), .C(n_872), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_855), .Y(n_851) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
BUFx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
BUFx2_ASAP7_75t_L g922 ( .A(n_864), .Y(n_922) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_864), .Y(n_1198) );
BUFx2_ASAP7_75t_L g1439 ( .A(n_864), .Y(n_1439) );
OR2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_870), .Y(n_866) );
OR2x6_ASAP7_75t_L g1040 ( .A(n_867), .B(n_870), .Y(n_1040) );
INVx2_ASAP7_75t_SL g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
BUFx3_ASAP7_75t_L g1025 ( .A(n_869), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_869), .Y(n_1036) );
BUFx4f_ASAP7_75t_L g1059 ( .A(n_869), .Y(n_1059) );
OR2x4_ASAP7_75t_L g1154 ( .A(n_869), .B(n_1136), .Y(n_1154) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_891), .B(n_904), .Y(n_876) );
BUFx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_888), .A2(n_1496), .B1(n_1497), .B2(n_1498), .Y(n_1495) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx2_ASAP7_75t_L g1452 ( .A(n_901), .Y(n_1452) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g1186 ( .A(n_902), .Y(n_1186) );
OAI21xp5_ASAP7_75t_L g929 ( .A1(n_904), .A2(n_930), .B(n_941), .Y(n_929) );
O2A1O1Ixp5_ASAP7_75t_L g1486 ( .A1(n_904), .A2(n_1487), .B(n_1499), .C(n_1509), .Y(n_1486) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_926), .C(n_929), .Y(n_907) );
NOR3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_924), .C(n_925), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_913), .Y(n_909) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g1075 ( .A(n_922), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_935), .B1(n_936), .B2(n_938), .C(n_939), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx6f_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx3_ASAP7_75t_L g1085 ( .A(n_934), .Y(n_1085) );
INVx5_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_SL g945 ( .A(n_946), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_1048), .B2(n_1049), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_988), .B1(n_989), .B2(n_1047), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_957), .Y(n_1047) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_975), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_970), .B1(n_972), .B2(n_974), .Y(n_966) );
INVx2_ASAP7_75t_L g1032 ( .A(n_971), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_980), .C(n_983), .Y(n_976) );
INVxp67_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NOR3xp33_ASAP7_75t_L g990 ( .A(n_991), .B(n_1041), .C(n_1046), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_1014), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_1002), .Y(n_995) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1000), .Y(n_1176) );
NAND3xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1009), .C(n_1012), .Y(n_1003) );
AOI21xp5_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1016), .B(n_1017), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1020), .B1(n_1021), .B2(n_1022), .Y(n_1018) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1026), .B1(n_1027), .B2(n_1028), .Y(n_1024) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B1(n_1037), .B2(n_1039), .Y(n_1034) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
OA22x2_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1051), .B1(n_1162), .B2(n_1163), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
NAND3xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1099), .C(n_1129), .Y(n_1052) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1080), .Y(n_1053) );
OAI33xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .A3(n_1062), .B1(n_1067), .B2(n_1075), .B3(n_1076), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1060), .B2(n_1061), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_1057), .A2(n_1077), .B1(n_1083), .B2(n_1086), .Y(n_1082) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_1058), .A2(n_1077), .B1(n_1078), .B2(n_1079), .Y(n_1076) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_1060), .A2(n_1079), .B1(n_1086), .B2(n_1090), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1065), .B2(n_1066), .Y(n_1062) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1064), .Y(n_1196) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_1065), .A2(n_1074), .B1(n_1093), .B2(n_1095), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1071), .B1(n_1072), .B2(n_1074), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx8_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
BUFx3_ASAP7_75t_L g1481 ( .A(n_1070), .Y(n_1481) );
BUFx6f_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1073), .Y(n_1139) );
OAI33xp33_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .A3(n_1089), .B1(n_1091), .B2(n_1092), .B3(n_1096), .Y(n_1080) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx2_ASAP7_75t_SL g1084 ( .A(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_1093), .A2(n_1182), .B1(n_1183), .B2(n_1184), .C(n_1185), .Y(n_1181) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
OAI31xp33_ASAP7_75t_SL g1099 ( .A1(n_1100), .A2(n_1112), .A3(n_1122), .B(n_1126), .Y(n_1099) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1108), .B1(n_1109), .B2(n_1110), .Y(n_1104) );
BUFx3_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1108), .A2(n_1143), .B1(n_1147), .B2(n_1150), .Y(n_1142) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx3_ASAP7_75t_SL g1124 ( .A(n_1125), .Y(n_1124) );
BUFx3_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
OAI31xp33_ASAP7_75t_SL g1129 ( .A1(n_1130), .A2(n_1137), .A3(n_1151), .B(n_1157), .Y(n_1129) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
CKINVDCx8_ASAP7_75t_R g1140 ( .A(n_1141), .Y(n_1140) );
BUFx3_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1146), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_1145), .B(n_1149), .Y(n_1148) );
BUFx6f_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx2_ASAP7_75t_SL g1153 ( .A(n_1154), .Y(n_1153) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
INVx1_ASAP7_75t_SL g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
AO21x2_ASAP7_75t_L g1163 ( .A1(n_1164), .A2(n_1165), .B(n_1204), .Y(n_1163) );
NAND3xp33_ASAP7_75t_SL g1165 ( .A(n_1166), .B(n_1169), .C(n_1188), .Y(n_1165) );
OAI21xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1179), .B(n_1187), .Y(n_1169) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1419), .B1(n_1422), .B2(n_1456), .C(n_1459), .Y(n_1205) );
AOI21xp5_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1310), .B(n_1331), .Y(n_1206) );
OAI211xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1227), .B(n_1258), .C(n_1296), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1223), .Y(n_1208) );
INVx3_ASAP7_75t_L g1267 ( .A(n_1209), .Y(n_1267) );
INVx3_ASAP7_75t_L g1307 ( .A(n_1209), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1209), .B(n_1284), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1209), .B(n_1330), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1209), .B(n_1352), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1209), .B(n_1223), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1209), .B(n_1276), .Y(n_1376) );
AND2x4_ASAP7_75t_SL g1209 ( .A(n_1210), .B(n_1217), .Y(n_1209) );
INVx2_ASAP7_75t_L g1421 ( .A(n_1211), .Y(n_1421) );
AND2x6_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1213), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1212), .B(n_1216), .Y(n_1215) );
AND2x4_ASAP7_75t_L g1218 ( .A(n_1212), .B(n_1219), .Y(n_1218) );
AND2x6_ASAP7_75t_L g1221 ( .A(n_1212), .B(n_1222), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1212), .B(n_1216), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1212), .B(n_1216), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1518 ( .A(n_1213), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1214), .B(n_1220), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1223), .B(n_1252), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1223), .B(n_1307), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1223), .B(n_1251), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1223), .B(n_1252), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1223), .B(n_1338), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1226), .Y(n_1223) );
AND2x4_ASAP7_75t_L g1271 ( .A(n_1224), .B(n_1226), .Y(n_1271) );
AOI211xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1236), .B(n_1244), .C(n_1249), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1228), .B(n_1288), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1228), .B(n_1283), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1228), .B(n_1248), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1232), .Y(n_1228) );
INVx3_ASAP7_75t_L g1247 ( .A(n_1229), .Y(n_1247) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1229), .Y(n_1280) );
NOR2xp33_ASAP7_75t_L g1314 ( .A(n_1229), .B(n_1232), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1229), .B(n_1364), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1229), .B(n_1251), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1229), .B(n_1400), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1231), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1232), .B(n_1275), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1232), .B(n_1257), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g1292 ( .A(n_1232), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1232), .B(n_1291), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1232), .B(n_1298), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1232), .B(n_1288), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1235), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1233), .B(n_1235), .Y(n_1260) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1236), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1383 ( .A(n_1236), .B(n_1247), .Y(n_1383) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1240), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1237), .B(n_1240), .Y(n_1248) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1237), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1237), .B(n_1241), .Y(n_1288) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1237), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1240), .B(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1240), .Y(n_1275) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1241), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1243), .Y(n_1241) );
INVxp67_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1248), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1246), .B(n_1274), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1246), .B(n_1276), .Y(n_1293) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1247), .B(n_1251), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1247), .B(n_1248), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1247), .B(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1247), .B(n_1343), .Y(n_1365) );
OAI21xp33_ASAP7_75t_L g1368 ( .A1(n_1247), .A2(n_1359), .B(n_1369), .Y(n_1368) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_1247), .B(n_1388), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1247), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1248), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1248), .B(n_1314), .Y(n_1350) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1255), .Y(n_1249) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1250), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1251), .B(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1252), .Y(n_1285) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1252), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1254), .Y(n_1252) );
NOR3xp33_ASAP7_75t_L g1378 ( .A(n_1255), .B(n_1307), .C(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1256), .B(n_1292), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1256), .B(n_1376), .Y(n_1375) );
OAI32xp33_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1262), .A3(n_1266), .B1(n_1268), .B2(n_1294), .Y(n_1258) );
AOI332xp33_ASAP7_75t_L g1384 ( .A1(n_1259), .A2(n_1267), .A3(n_1324), .B1(n_1330), .B2(n_1352), .B3(n_1385), .C1(n_1387), .C2(n_1389), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1261), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1260), .B(n_1283), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1260), .B(n_1328), .Y(n_1359) );
AOI22xp5_ASAP7_75t_SL g1269 ( .A1(n_1261), .A2(n_1270), .B1(n_1272), .B2(n_1276), .Y(n_1269) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1262), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1262), .B(n_1267), .Y(n_1319) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_1262), .A2(n_1263), .B1(n_1398), .B2(n_1406), .Y(n_1397) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
AOI211xp5_ASAP7_75t_L g1312 ( .A1(n_1263), .A2(n_1313), .B(n_1315), .C(n_1316), .Y(n_1312) );
O2A1O1Ixp33_ASAP7_75t_SL g1354 ( .A1(n_1263), .A2(n_1355), .B(n_1356), .C(n_1357), .Y(n_1354) );
O2A1O1Ixp33_ASAP7_75t_L g1361 ( .A1(n_1263), .A2(n_1362), .B(n_1372), .C(n_1380), .Y(n_1361) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1263), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1265), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1266), .B(n_1295), .Y(n_1294) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g1310 ( .A1(n_1267), .A2(n_1311), .B1(n_1312), .B2(n_1319), .C(n_1320), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1395 ( .A1(n_1267), .A2(n_1396), .B1(n_1397), .B2(n_1410), .Y(n_1395) );
INVxp67_ASAP7_75t_SL g1311 ( .A(n_1268), .Y(n_1311) );
NAND4xp25_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1277), .C(n_1286), .D(n_1289), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1270), .B(n_1287), .Y(n_1286) );
NAND2xp5_ASAP7_75t_SL g1300 ( .A(n_1270), .B(n_1280), .Y(n_1300) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1270), .Y(n_1355) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1271), .Y(n_1330) );
CKINVDCx6p67_ASAP7_75t_R g1335 ( .A(n_1271), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1271), .B(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
AOI21xp33_ASAP7_75t_L g1404 ( .A1(n_1273), .A2(n_1279), .B(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1274), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1275), .B(n_1292), .Y(n_1303) );
CKINVDCx14_ASAP7_75t_R g1405 ( .A(n_1276), .Y(n_1405) );
OAI21xp5_ASAP7_75t_L g1277 ( .A1(n_1278), .A2(n_1282), .B(n_1284), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_1278), .A2(n_1367), .B1(n_1368), .B2(n_1370), .Y(n_1366) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1281), .Y(n_1279) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1280), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1280), .B(n_1386), .Y(n_1385) );
NAND2xp5_ASAP7_75t_SL g1394 ( .A(n_1280), .B(n_1283), .Y(n_1394) );
CKINVDCx14_ASAP7_75t_R g1344 ( .A(n_1281), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g1374 ( .A(n_1282), .Y(n_1374) );
OAI21xp5_ASAP7_75t_L g1289 ( .A1(n_1283), .A2(n_1290), .B(n_1293), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1283), .B(n_1314), .Y(n_1313) );
OAI21xp5_ASAP7_75t_L g1357 ( .A1(n_1283), .A2(n_1293), .B(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1284), .Y(n_1318) );
OAI21xp33_ASAP7_75t_L g1391 ( .A1(n_1284), .A2(n_1329), .B(n_1392), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1284), .B(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
OAI21xp5_ASAP7_75t_SL g1349 ( .A1(n_1285), .A2(n_1350), .B(n_1351), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1287), .B(n_1318), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1288), .B(n_1292), .Y(n_1343) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1288), .Y(n_1400) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1290), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1292), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1292), .B(n_1328), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1292), .B(n_1383), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1292), .B(n_1394), .Y(n_1393) );
A2O1A1Ixp33_ASAP7_75t_L g1296 ( .A1(n_1297), .A2(n_1299), .B(n_1301), .C(n_1304), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1298), .B(n_1314), .Y(n_1356) );
INVxp67_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1308), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1307), .B(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1347 ( .A(n_1315), .B(n_1348), .Y(n_1347) );
A2O1A1Ixp33_ASAP7_75t_L g1362 ( .A1(n_1315), .A2(n_1363), .B(n_1365), .C(n_1366), .Y(n_1362) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_1315), .Y(n_1403) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
AOI211xp5_ASAP7_75t_L g1332 ( .A1(n_1319), .A2(n_1333), .B(n_1354), .C(n_1360), .Y(n_1332) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1324), .B1(n_1326), .B2(n_1329), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1360 ( .A(n_1322), .B(n_1327), .Y(n_1360) );
OAI211xp5_ASAP7_75t_SL g1380 ( .A1(n_1322), .A2(n_1381), .B(n_1384), .C(n_1391), .Y(n_1380) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1323), .Y(n_1386) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1328), .B(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1329), .Y(n_1373) );
A2O1A1Ixp33_ASAP7_75t_L g1410 ( .A1(n_1330), .A2(n_1353), .B(n_1411), .C(n_1412), .Y(n_1410) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_1330), .A2(n_1403), .B1(n_1413), .B2(n_1414), .C(n_1417), .Y(n_1412) );
NAND3xp33_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1361), .C(n_1395), .Y(n_1331) );
OAI211xp5_ASAP7_75t_L g1333 ( .A1(n_1334), .A2(n_1336), .B(n_1340), .C(n_1349), .Y(n_1333) );
CKINVDCx6p67_ASAP7_75t_R g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
AOI211xp5_ASAP7_75t_L g1406 ( .A1(n_1337), .A2(n_1352), .B(n_1407), .C(n_1408), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_1338), .B(n_1388), .Y(n_1407) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1339), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g1340 ( .A1(n_1341), .A2(n_1345), .B(n_1347), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1344), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1343), .B(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1353), .Y(n_1351) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1365), .Y(n_1413) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B(n_1375), .C(n_1377), .Y(n_1372) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_1378), .Y(n_1377) );
NAND2xp5_ASAP7_75t_SL g1414 ( .A(n_1381), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
AOI211xp5_ASAP7_75t_L g1398 ( .A1(n_1386), .A2(n_1399), .B(n_1401), .C(n_1404), .Y(n_1398) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_1389), .Y(n_1396) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1408), .Y(n_1411) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
CKINVDCx20_ASAP7_75t_R g1419 ( .A(n_1420), .Y(n_1419) );
CKINVDCx20_ASAP7_75t_R g1420 ( .A(n_1421), .Y(n_1420) );
BUFx3_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1441), .Y(n_1424) );
INVx2_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
NAND3xp33_ASAP7_75t_SL g1442 ( .A(n_1443), .B(n_1446), .C(n_1449), .Y(n_1442) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx2_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
HB1xp67_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
BUFx3_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVxp33_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
NAND3x1_ASAP7_75t_SL g1468 ( .A(n_1469), .B(n_1486), .C(n_1512), .Y(n_1468) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
HB1xp67_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx4_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx2_ASAP7_75t_SL g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
OAI21xp5_ASAP7_75t_L g1517 ( .A1(n_1518), .A2(n_1519), .B(n_1520), .Y(n_1517) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
endmodule