module fake_netlist_1_9960_n_730 (n_117, n_44, n_133, n_149, n_81, n_69, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_730);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_730;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_230;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_188), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_98), .Y(n_215) );
INVxp33_ASAP7_75t_SL g216 ( .A(n_85), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_43), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_200), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_59), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_205), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
INVxp67_ASAP7_75t_L g222 ( .A(n_100), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_57), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_58), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_78), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_167), .B(n_159), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_147), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_55), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_30), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_40), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_211), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_148), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_163), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_197), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_113), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_28), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_32), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_52), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_64), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_90), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_7), .B(n_48), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_138), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_177), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_91), .Y(n_244) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_174), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_126), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_201), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_15), .Y(n_248) );
INVxp33_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_166), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_119), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_38), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_111), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_180), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_208), .Y(n_257) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_67), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_51), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_61), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_22), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_192), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_45), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_34), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_191), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_13), .Y(n_266) );
BUFx10_ASAP7_75t_L g267 ( .A(n_153), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_37), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_31), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_120), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_99), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g272 ( .A(n_199), .B(n_20), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_178), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_83), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_50), .B(n_81), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_1), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_189), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_82), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_103), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_3), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_134), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_69), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_106), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_123), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_140), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_170), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_20), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_179), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_196), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_35), .B(n_168), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_6), .B(n_129), .Y(n_293) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_127), .Y(n_294) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_14), .B(n_95), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_115), .Y(n_296) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_173), .B(n_183), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_72), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_203), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_110), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_76), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_194), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_93), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_161), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_114), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_8), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_162), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_71), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_75), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_63), .Y(n_310) );
INVxp33_ASAP7_75t_SL g311 ( .A(n_128), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_77), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_23), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_101), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_73), .Y(n_315) );
XOR2xp5_ASAP7_75t_L g316 ( .A(n_198), .B(n_46), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_107), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_84), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_97), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_87), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_136), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_190), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_185), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_86), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_70), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_158), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_229), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_267), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_267), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_229), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_249), .B(n_0), .Y(n_331) );
BUFx8_ASAP7_75t_L g332 ( .A(n_276), .Y(n_332) );
XOR2x2_ASAP7_75t_L g333 ( .A(n_241), .B(n_2), .Y(n_333) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_263), .B(n_24), .Y(n_334) );
INVx5_ASAP7_75t_L g335 ( .A(n_223), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_277), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_282), .B(n_224), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_275), .B(n_2), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_309), .B(n_3), .Y(n_339) );
CKINVDCx6p67_ASAP7_75t_R g340 ( .A(n_217), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_230), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_231), .Y(n_342) );
OAI22xp5_ASAP7_75t_SL g343 ( .A1(n_261), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_215), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_218), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_222), .B(n_4), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_223), .Y(n_347) );
BUFx12f_ASAP7_75t_L g348 ( .A(n_214), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_246), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_251), .A2(n_26), .B(n_25), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_223), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_280), .B(n_5), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_219), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_220), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_343), .B(n_272), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_352), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_352), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_344), .B(n_310), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_328), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_345), .B(n_221), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_330), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_330), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_328), .B(n_222), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_353), .B(n_225), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_347), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_337), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_245), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_348), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_339), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_347), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_329), .B(n_228), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_337), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
AND2x6_ASAP7_75t_L g379 ( .A(n_338), .B(n_236), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_373), .A2(n_350), .B(n_354), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_365), .B(n_329), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_350), .B(n_338), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_365), .B(n_340), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_355), .A2(n_313), .B1(n_289), .B2(n_331), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_369), .B(n_334), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_360), .B(n_340), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_379), .A2(n_334), .B1(n_338), .B2(n_341), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_364), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_368), .A2(n_331), .B(n_346), .C(n_342), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_362), .B(n_332), .Y(n_392) );
AO22x1_ASAP7_75t_L g393 ( .A1(n_375), .A2(n_311), .B1(n_216), .B2(n_258), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_379), .A2(n_324), .B1(n_258), .B2(n_239), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_379), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_362), .B(n_349), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_376), .B(n_349), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_358), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_376), .B(n_294), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_370), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_371), .B(n_324), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_356), .B(n_232), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_355), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_379), .B(n_233), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_379), .B(n_234), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_377), .B(n_235), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_361), .B(n_237), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_361), .B(n_240), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_366), .B(n_247), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_366), .B(n_252), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_394), .B(n_359), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_382), .A2(n_359), .B(n_363), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_243), .B(n_238), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_394), .B(n_248), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_401), .B(n_388), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_401), .B(n_266), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_388), .B(n_306), .Y(n_419) );
INVx5_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_381), .A2(n_250), .B(n_244), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_397), .A2(n_255), .B(n_253), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_383), .A2(n_259), .B(n_256), .Y(n_423) );
AND2x6_ASAP7_75t_L g424 ( .A(n_395), .B(n_262), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_386), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_399), .A2(n_265), .B(n_264), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_402), .A2(n_274), .B(n_270), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_385), .A2(n_242), .B1(n_271), .B2(n_260), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_386), .B(n_273), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_409), .A2(n_323), .B1(n_296), .B2(n_333), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_409), .A2(n_333), .B1(n_316), .B2(n_286), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_395), .B(n_254), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_404), .A2(n_287), .B(n_284), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_393), .B(n_247), .Y(n_434) );
OR2x6_ASAP7_75t_L g435 ( .A(n_400), .B(n_293), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_391), .B(n_307), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_406), .B(n_257), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_405), .A2(n_291), .B(n_290), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_407), .B(n_268), .Y(n_441) );
AO22x1_ASAP7_75t_L g442 ( .A1(n_424), .A2(n_403), .B1(n_384), .B2(n_322), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_425), .B(n_410), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_412), .A2(n_408), .B(n_390), .Y(n_444) );
BUFx5_ASAP7_75t_L g445 ( .A(n_424), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_416), .B(n_389), .Y(n_446) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_414), .A2(n_297), .B(n_292), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_438), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_426), .A2(n_300), .B(n_299), .Y(n_449) );
BUFx10_ASAP7_75t_L g450 ( .A(n_424), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_411), .A2(n_314), .B(n_302), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_423), .A2(n_295), .B(n_318), .C(n_326), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_417), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_429), .A2(n_279), .B(n_269), .Y(n_455) );
OAI21x1_ASAP7_75t_L g456 ( .A1(n_433), .A2(n_325), .B(n_317), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_440), .A2(n_374), .B(n_367), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_431), .A2(n_321), .B1(n_281), .B2(n_283), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_418), .B(n_336), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_436), .A2(n_378), .B(n_374), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_438), .B(n_320), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_420), .Y(n_462) );
AO22x2_ASAP7_75t_L g463 ( .A1(n_434), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_9), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_421), .A2(n_226), .B(n_378), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_441), .A2(n_288), .B(n_285), .Y(n_467) );
AO31x2_ASAP7_75t_L g468 ( .A1(n_422), .A2(n_351), .A3(n_305), .B(n_315), .Y(n_468) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_427), .A2(n_303), .B(n_301), .Y(n_469) );
OAI21x1_ASAP7_75t_L g470 ( .A1(n_432), .A2(n_278), .B(n_227), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_428), .Y(n_471) );
AO32x2_ASAP7_75t_L g472 ( .A1(n_437), .A2(n_351), .A3(n_278), .B1(n_298), .B2(n_305), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_439), .A2(n_308), .B(n_304), .Y(n_473) );
OAI21x1_ASAP7_75t_L g474 ( .A1(n_419), .A2(n_278), .B(n_227), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_464), .B(n_435), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_471), .B(n_312), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_462), .Y(n_477) );
AOI21x1_ASAP7_75t_L g478 ( .A1(n_474), .A2(n_351), .B(n_305), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_454), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_446), .B(n_11), .Y(n_481) );
OAI21x1_ASAP7_75t_L g482 ( .A1(n_470), .A2(n_315), .B(n_298), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_444), .A2(n_372), .B(n_335), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_451), .A2(n_335), .B(n_319), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_465), .B(n_11), .Y(n_485) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_447), .A2(n_351), .B(n_315), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_460), .A2(n_372), .B(n_335), .Y(n_488) );
AO31x2_ASAP7_75t_L g489 ( .A1(n_452), .A2(n_298), .A3(n_335), .B(n_372), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_463), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_468), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_449), .B(n_12), .Y(n_492) );
OAI21x1_ASAP7_75t_L g493 ( .A1(n_457), .A2(n_132), .B(n_213), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_450), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_459), .A2(n_131), .B(n_212), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_466), .A2(n_130), .B(n_207), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_461), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_468), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_443), .A2(n_125), .B(n_204), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_458), .B(n_16), .Y(n_500) );
OAI21x1_ASAP7_75t_L g501 ( .A1(n_456), .A2(n_124), .B(n_202), .Y(n_501) );
AO31x2_ASAP7_75t_L g502 ( .A1(n_468), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_445), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_469), .A2(n_467), .B(n_473), .Y(n_504) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_472), .A2(n_122), .B(n_195), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_455), .A2(n_17), .B1(n_18), .B2(n_19), .C(n_21), .Y(n_506) );
OAI21x1_ASAP7_75t_L g507 ( .A1(n_469), .A2(n_135), .B(n_193), .Y(n_507) );
BUFx12f_ASAP7_75t_L g508 ( .A(n_450), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_472), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_472), .B(n_23), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_444), .A2(n_27), .B(n_29), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_454), .B(n_33), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_442), .A2(n_36), .B1(n_39), .B2(n_41), .C(n_42), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_474), .A2(n_44), .B(n_47), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_49), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_479), .B(n_53), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_485), .B(n_54), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_512), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_475), .B(n_56), .Y(n_521) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_509), .A2(n_60), .B(n_62), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_508), .Y(n_523) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_491), .A2(n_65), .B(n_66), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_498), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_511), .Y(n_526) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_483), .A2(n_68), .B(n_74), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_497), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_511), .Y(n_529) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_478), .A2(n_79), .B(n_80), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_481), .Y(n_531) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_490), .B(n_88), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_513), .A2(n_89), .B(n_92), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_492), .Y(n_534) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_516), .A2(n_94), .B(n_96), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_510), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_494), .Y(n_537) );
OR2x6_ASAP7_75t_L g538 ( .A(n_475), .B(n_102), .Y(n_538) );
OR2x6_ASAP7_75t_L g539 ( .A(n_503), .B(n_104), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_514), .Y(n_540) );
OR2x6_ASAP7_75t_L g541 ( .A(n_487), .B(n_105), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_501), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_502), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_489), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_489), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_500), .B(n_108), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_486), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_486), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_504), .B(n_109), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_476), .B(n_112), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_484), .B(n_116), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_515), .B(n_117), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_493), .B(n_118), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_513), .B(n_121), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_507), .Y(n_556) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_482), .A2(n_133), .B(n_137), .Y(n_557) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_488), .A2(n_139), .B(n_141), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_506), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_499), .B(n_142), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_505), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_484), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_495), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_496), .Y(n_564) );
OAI21x1_ASAP7_75t_L g565 ( .A1(n_478), .A2(n_143), .B(n_144), .Y(n_565) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_478), .A2(n_145), .B(n_146), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_477), .Y(n_567) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_478), .A2(n_149), .B(n_150), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_480), .B(n_151), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_479), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_480), .B(n_152), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_491), .Y(n_572) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_478), .A2(n_154), .B(n_155), .Y(n_573) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_509), .A2(n_156), .B(n_157), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_543), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_567), .Y(n_577) );
INVx4_ASAP7_75t_L g578 ( .A(n_541), .Y(n_578) );
INVx4_ASAP7_75t_L g579 ( .A(n_541), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_570), .B(n_160), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_544), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_536), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_526), .B(n_165), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_519), .B(n_169), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_531), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_528), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_537), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_534), .B(n_172), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_532), .B(n_176), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_518), .Y(n_591) );
BUFx2_ASAP7_75t_L g592 ( .A(n_537), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
OR2x6_ASAP7_75t_SL g594 ( .A(n_547), .B(n_181), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_541), .B(n_182), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_538), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_536), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_525), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_571), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_521), .B(n_184), .Y(n_601) );
INVx5_ASAP7_75t_L g602 ( .A(n_539), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_539), .B(n_186), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_539), .B(n_187), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_549), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_571), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_572), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_523), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_517), .B(n_569), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_532), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_559), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_540), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_545), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_551), .B(n_562), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_551), .B(n_562), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_553), .B(n_552), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_555), .A2(n_550), .B1(n_554), .B2(n_552), .Y(n_618) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_546), .Y(n_619) );
AND2x4_ASAP7_75t_SL g620 ( .A(n_554), .B(n_560), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_564), .B(n_563), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_522), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_574), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_560), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_527), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_527), .B(n_564), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_524), .B(n_533), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_542), .B(n_524), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_533), .A2(n_561), .B1(n_535), .B2(n_542), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_548), .B(n_556), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_599), .B(n_548), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_599), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_594), .B(n_535), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_584), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_588), .B(n_558), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_586), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_576), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_598), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_605), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_607), .B(n_557), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_608), .B(n_530), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_575), .Y(n_642) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_608), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_614), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_620), .B(n_565), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_620), .B(n_566), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_624), .B(n_568), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_612), .B(n_573), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_592), .B(n_587), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_617), .A2(n_615), .B1(n_616), .B2(n_578), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_581), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_587), .B(n_582), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_613), .B(n_596), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_597), .B(n_578), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_593), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_610), .B(n_579), .Y(n_656) );
BUFx3_ASAP7_75t_L g657 ( .A(n_609), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_600), .B(n_606), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_621), .Y(n_659) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_595), .B(n_604), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_624), .B(n_591), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_602), .B(n_628), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_618), .B(n_580), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_614), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_590), .A2(n_627), .B(n_602), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_589), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_619), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_602), .B(n_628), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_630), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_626), .B(n_619), .Y(n_671) );
NOR2xp67_ASAP7_75t_L g672 ( .A(n_633), .B(n_611), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_671), .B(n_625), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_660), .A2(n_603), .B1(n_604), .B2(n_577), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_670), .B(n_623), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_663), .B(n_611), .Y(n_676) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_668), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_658), .B(n_622), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_659), .B(n_629), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_657), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_661), .B(n_629), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_632), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_631), .B(n_639), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_638), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_641), .B(n_590), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_649), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_641), .B(n_603), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_642), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_634), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_636), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_651), .B(n_583), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_674), .A2(n_633), .B1(n_650), .B2(n_664), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_686), .B(n_643), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_680), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_682), .B(n_665), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_673), .B(n_653), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_690), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_689), .B(n_656), .Y(n_698) );
AND2x4_ASAP7_75t_SL g699 ( .A(n_689), .B(n_652), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_684), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_679), .B(n_637), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_687), .B(n_662), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_679), .B(n_655), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_681), .B(n_644), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_677), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_694), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_692), .A2(n_672), .B1(n_687), .B2(n_654), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_699), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_704), .B(n_705), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_695), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_693), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_701), .B(n_675), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_709), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_707), .A2(n_703), .B1(n_698), .B2(n_696), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_711), .B(n_702), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_708), .B(n_700), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_706), .A2(n_667), .B(n_697), .Y(n_717) );
AOI211xp5_ASAP7_75t_SL g718 ( .A1(n_710), .A2(n_666), .B(n_676), .C(n_685), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_712), .A2(n_585), .B(n_645), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g720 ( .A1(n_718), .A2(n_714), .B(n_716), .C(n_717), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_713), .A2(n_715), .B(n_719), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_720), .B(n_585), .C(n_601), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_722), .B(n_721), .C(n_648), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_723), .B(n_683), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_724), .A2(n_646), .B1(n_645), .B2(n_663), .Y(n_725) );
OAI22x1_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_647), .B1(n_669), .B2(n_663), .Y(n_726) );
AOI22x1_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_647), .B1(n_669), .B2(n_635), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_727), .B(n_688), .Y(n_728) );
OR2x6_ASAP7_75t_L g729 ( .A(n_728), .B(n_691), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_640), .B(n_678), .Y(n_730) );
endmodule