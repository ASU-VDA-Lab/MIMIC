module real_jpeg_15928_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_0),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_0),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_0),
.B(n_135),
.Y(n_134)
);

NAND2x1p5_ASAP7_75t_L g155 ( 
.A(n_0),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_0),
.B(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_3),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_9),
.B1(n_109),
.B2(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_50),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_4),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_85),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_6),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_7),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_7),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_7),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_7),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_8),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_8),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_8),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_8),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_8),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_8),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_9),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_9),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_9),
.B(n_317),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_11),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_11),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_11),
.B(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_14),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_14),
.B(n_71),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_14),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_14),
.B(n_261),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_14),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_14),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_14),
.B(n_331),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_192),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_191),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_141),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_20),
.B(n_141),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.C(n_118),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_21),
.B(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_61),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_23),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_26),
.B(n_35),
.C(n_36),
.Y(n_190)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_41),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_43),
.A2(n_47),
.B(n_52),
.C(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_46),
.B(n_51),
.Y(n_165)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_49),
.Y(n_327)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.C(n_57),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_53),
.A2(n_57),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_60),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_61),
.B(n_143),
.C(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.C(n_83),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_62),
.B(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_66),
.C(n_70),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_74),
.A2(n_75),
.B1(n_83),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_78),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_79),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_81),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_82),
.Y(n_336)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.C(n_90),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_84),
.A2(n_90),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_84),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_87),
.B(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_90),
.Y(n_207)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_92),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_93),
.B(n_118),
.Y(n_195)
);

XOR2x2_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_108),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_107),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_149),
.C(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_96),
.B(n_100),
.C(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_106),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_103),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_SL g232 ( 
.A(n_106),
.B(n_134),
.Y(n_232)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_124),
.B(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_111),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_132),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_123),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_125),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_132),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_139),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_133),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_230)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_168),
.B2(n_169),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_162),
.B2(n_163),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_162),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_188),
.B(n_240),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_221),
.B(n_347),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_194),
.B(n_196),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_203),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_204),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.C(n_217),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_217),
.Y(n_270)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_248),
.B(n_346),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_245),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_225),
.B(n_245),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_226),
.A2(n_227),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_229),
.B(n_231),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.C(n_239),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_244),
.Y(n_315)
);

AOI21x1_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_274),
.B(n_345),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_271),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_250),
.B(n_271),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_269),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_269),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.C(n_266),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_266),
.Y(n_279)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_293),
.B(n_344),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_291),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_276),
.B(n_291),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_289),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_278),
.B1(n_304),
.B2(n_306),
.Y(n_303)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_289),
.B1(n_290),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_307),
.B(n_343),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_295),
.B(n_303),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.C(n_301),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_301),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_304),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_322),
.B(n_342),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_319),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_309),
.B(n_319),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_316),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_316),
.Y(n_328)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_329),
.B(n_341),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_324),
.B(n_328),
.Y(n_341)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);


endmodule