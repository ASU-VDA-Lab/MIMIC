module fake_jpeg_918_n_510 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_510);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_0),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_57),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_19),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_38),
.B1(n_53),
.B2(n_40),
.Y(n_130)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_76),
.Y(n_122)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_77),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_78),
.Y(n_181)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_36),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_80),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_83),
.Y(n_198)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_91),
.Y(n_193)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_94),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_18),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_97),
.B(n_100),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_33),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_51),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_13),
.Y(n_124)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_117),
.Y(n_165)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_47),
.B(n_16),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_116),
.B(n_5),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_124),
.B(n_132),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_55),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_129),
.B(n_134),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_130),
.A2(n_88),
.B1(n_113),
.B2(n_98),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_55),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_48),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_42),
.B1(n_29),
.B2(n_52),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_136),
.A2(n_151),
.B1(n_154),
.B2(n_175),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_42),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_141),
.B(n_144),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_58),
.B(n_37),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_51),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_145),
.B(n_159),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_66),
.A2(n_38),
.B1(n_37),
.B2(n_41),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_80),
.A2(n_51),
.B1(n_52),
.B2(n_41),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_64),
.B(n_40),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_30),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_161),
.B(n_169),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_71),
.B(n_30),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_81),
.A2(n_82),
.B1(n_69),
.B2(n_56),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_31),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_177),
.B(n_189),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_83),
.A2(n_31),
.B1(n_29),
.B2(n_22),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_180),
.A2(n_190),
.B1(n_197),
.B2(n_154),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_85),
.B(n_16),
.C(n_22),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_11),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_16),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_81),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_121),
.B(n_2),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_191),
.B(n_204),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_91),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_200),
.B(n_140),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_93),
.B(n_6),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_206),
.Y(n_284)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

BUFx2_ASAP7_75t_SL g310 ( 
.A(n_207),
.Y(n_310)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_211),
.A2(n_225),
.B1(n_274),
.B2(n_185),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_122),
.A2(n_119),
.B(n_95),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_260),
.C(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_171),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_213),
.Y(n_319)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_214),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_90),
.B1(n_109),
.B2(n_8),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_215),
.A2(n_152),
.B1(n_158),
.B2(n_202),
.Y(n_301)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_164),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

BUFx6f_ASAP7_75t_SL g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_220),
.Y(n_315)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_7),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_223),
.B(n_243),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_224),
.B(n_228),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_126),
.B(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_226),
.B(n_232),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_231),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_137),
.B(n_10),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_233),
.A2(n_264),
.B(n_266),
.Y(n_322)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_139),
.Y(n_234)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_186),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_238),
.Y(n_320)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_125),
.Y(n_239)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_241),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_242),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_164),
.A2(n_11),
.B1(n_12),
.B2(n_143),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_244),
.A2(n_251),
.B1(n_261),
.B2(n_265),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_246),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_160),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_135),
.B(n_11),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_254),
.Y(n_305)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_153),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_149),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_256),
.Y(n_290)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_149),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_257),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_175),
.A2(n_163),
.B1(n_157),
.B2(n_166),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_258),
.A2(n_230),
.B1(n_209),
.B2(n_261),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_197),
.A2(n_190),
.B(n_167),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_171),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_156),
.Y(n_262)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_146),
.B(n_168),
.CI(n_196),
.CON(n_263),
.SN(n_263)
);

MAJIxp5_ASAP7_75t_SL g306 ( 
.A(n_263),
.B(n_264),
.C(n_259),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_172),
.B(n_179),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_183),
.A2(n_150),
.B1(n_205),
.B2(n_203),
.Y(n_265)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_131),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_267),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_155),
.B(n_185),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_269),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_155),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_156),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_272),
.Y(n_296)
);

AO22x1_ASAP7_75t_SL g271 ( 
.A1(n_183),
.A2(n_198),
.B1(n_199),
.B2(n_158),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_275),
.B1(n_243),
.B2(n_253),
.Y(n_304)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_131),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_127),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_192),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_304),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_211),
.A2(n_192),
.B1(n_127),
.B2(n_133),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_300),
.B1(n_307),
.B2(n_271),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_229),
.A2(n_133),
.B1(n_150),
.B2(n_182),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_316),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_240),
.A2(n_236),
.B1(n_212),
.B2(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_217),
.A2(n_152),
.B1(n_173),
.B2(n_174),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_276),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_226),
.A2(n_232),
.B1(n_260),
.B2(n_233),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_209),
.B(n_227),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_238),
.C(n_210),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_252),
.A2(n_233),
.B(n_263),
.C(n_264),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_323),
.B(n_220),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_285),
.A2(n_323),
.B(n_303),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_326),
.A2(n_337),
.B(n_354),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_284),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_258),
.C(n_206),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_329),
.C(n_331),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_214),
.C(n_239),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_275),
.C(n_213),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_332),
.Y(n_369)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_279),
.A2(n_263),
.B1(n_267),
.B2(n_272),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_334),
.A2(n_335),
.B1(n_340),
.B2(n_355),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_336),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_237),
.B(n_255),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_325),
.A2(n_231),
.B1(n_234),
.B2(n_257),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_344),
.B1(n_347),
.B2(n_360),
.Y(n_370)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_341),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_279),
.A2(n_271),
.B1(n_219),
.B2(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_352),
.B(n_353),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_346),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_321),
.A2(n_316),
.B1(n_304),
.B2(n_306),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_247),
.B1(n_250),
.B2(n_262),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_345),
.A2(n_291),
.B1(n_278),
.B2(n_293),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_270),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_304),
.A2(n_322),
.B1(n_298),
.B2(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_357),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_277),
.B(n_286),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_319),
.B(n_304),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_290),
.A2(n_305),
.B1(n_281),
.B2(n_296),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_294),
.A2(n_296),
.B(n_278),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_356),
.B(n_289),
.CI(n_347),
.CON(n_389),
.SN(n_389)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_313),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_318),
.B(n_291),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_277),
.A2(n_295),
.B1(n_286),
.B2(n_318),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_292),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_363),
.Y(n_386)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_324),
.A3(n_320),
.B1(n_315),
.B2(n_314),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_367),
.A2(n_375),
.B1(n_380),
.B2(n_381),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_324),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_378),
.C(n_379),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_330),
.A2(n_310),
.B1(n_317),
.B2(n_320),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_359),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_392),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_314),
.C(n_284),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_341),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_288),
.B1(n_287),
.B2(n_309),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_343),
.A2(n_293),
.B1(n_288),
.B2(n_287),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_330),
.A2(n_289),
.B1(n_309),
.B2(n_328),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_390),
.B1(n_391),
.B2(n_372),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_389),
.A2(n_357),
.B1(n_351),
.B2(n_362),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_326),
.A2(n_337),
.B1(n_346),
.B2(n_344),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_348),
.B1(n_345),
.B2(n_327),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_356),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_332),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_358),
.B1(n_363),
.B2(n_350),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_394),
.A2(n_349),
.B1(n_339),
.B2(n_336),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_395),
.A2(n_413),
.B(n_420),
.Y(n_423)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_396),
.Y(n_428)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_385),
.Y(n_397)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_378),
.C(n_390),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_399),
.B(n_411),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_404),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_371),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_405),
.Y(n_424)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_407),
.B(n_409),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_332),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_410),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_335),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_386),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_386),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_412),
.A2(n_415),
.B1(n_418),
.B2(n_383),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_376),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_394),
.B1(n_393),
.B2(n_375),
.Y(n_430)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_335),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_419),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_369),
.B(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_387),
.A2(n_392),
.B(n_377),
.Y(n_420)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_364),
.B1(n_370),
.B2(n_383),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_422),
.A2(n_425),
.B1(n_409),
.B2(n_406),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_402),
.A2(n_364),
.B1(n_370),
.B2(n_391),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_368),
.B(n_388),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_439),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_430),
.A2(n_433),
.B1(n_441),
.B2(n_422),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_373),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_432),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_414),
.A2(n_380),
.B1(n_389),
.B2(n_382),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_389),
.C(n_381),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_419),
.C(n_398),
.Y(n_446)
);

FAx1_ASAP7_75t_SL g436 ( 
.A(n_420),
.B(n_366),
.CI(n_367),
.CON(n_436),
.SN(n_436)
);

MAJx2_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_439),
.C(n_438),
.Y(n_459)
);

NAND2xp67_ASAP7_75t_SL g444 ( 
.A(n_438),
.B(n_413),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_401),
.A2(n_369),
.B(n_403),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_401),
.A2(n_405),
.B1(n_415),
.B2(n_418),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_427),
.A2(n_396),
.B1(n_407),
.B2(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_443),
.B(n_447),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_446),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_445),
.A2(n_442),
.B1(n_434),
.B2(n_437),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_431),
.B(n_440),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_400),
.C(n_397),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_450),
.C(n_455),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_404),
.C(n_429),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_429),
.B(n_423),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_451),
.B(n_453),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_441),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_424),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_454),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_425),
.C(n_421),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_456),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_428),
.C(n_423),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_426),
.C(n_434),
.Y(n_464)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_459),
.Y(n_472)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_457),
.Y(n_461)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_465),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_428),
.C(n_434),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_467),
.A2(n_436),
.B1(n_437),
.B2(n_446),
.Y(n_481)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_444),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_449),
.C(n_455),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_473),
.B(n_474),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_472),
.A2(n_452),
.B(n_442),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_453),
.B(n_459),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_477),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_447),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_463),
.Y(n_480)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_480),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_466),
.B(n_448),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_448),
.C(n_460),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_475),
.A2(n_470),
.B1(n_471),
.B2(n_467),
.Y(n_485)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_477),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_482),
.A2(n_471),
.B1(n_468),
.B2(n_464),
.Y(n_490)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_490),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_466),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_476),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_481),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_492),
.B(n_495),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_473),
.C(n_462),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_496),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_496),
.B(n_491),
.Y(n_499)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_497),
.B(n_486),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_488),
.B(n_492),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_498),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_504),
.A2(n_505),
.B(n_500),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_503),
.Y(n_505)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_493),
.B(n_489),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_484),
.B(n_480),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_508),
.A2(n_479),
.B(n_483),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_509),
.B(n_436),
.Y(n_510)
);


endmodule