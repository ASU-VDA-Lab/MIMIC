module real_jpeg_27335_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_299;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_293;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_0),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_0),
.A2(n_115),
.B(n_173),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_77),
.B1(n_78),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_1),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_156),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_156),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_1),
.A2(n_48),
.B1(n_51),
.B2(n_156),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_3),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_3),
.B(n_27),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_27),
.B(n_196),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_154),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_11),
.B(n_48),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_121),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_3),
.A2(n_89),
.B1(n_143),
.B2(n_244),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_5),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_77),
.B1(n_78),
.B2(n_150),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_150),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_5),
.A2(n_48),
.B1(n_51),
.B2(n_150),
.Y(n_236)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_41),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_7),
.A2(n_41),
.B1(n_48),
.B2(n_51),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_45),
.B1(n_77),
.B2(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_9),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_48),
.B1(n_51),
.B2(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_39),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_39),
.B1(n_48),
.B2(n_51),
.Y(n_173)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_56)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_14),
.A2(n_77),
.B1(n_78),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_14),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_127),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_14),
.A2(n_48),
.B1(n_51),
.B2(n_127),
.Y(n_231)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_60),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_24),
.B(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_37),
.B2(n_40),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_25),
.A2(n_31),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_25),
.A2(n_31),
.B1(n_149),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_25),
.A2(n_31),
.B1(n_182),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_27),
.A2(n_28),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_27),
.B(n_74),
.Y(n_170)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_28),
.A2(n_81),
.B1(n_153),
.B2(n_170),
.Y(n_169)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_28),
.A2(n_32),
.A3(n_35),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_31),
.B(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_33),
.B(n_36),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_33),
.A2(n_50),
.B(n_154),
.C(n_223),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_38),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_43),
.A2(n_55),
.B(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_46),
.B(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_55),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_47),
.A2(n_55),
.B1(n_99),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_47),
.A2(n_53),
.B(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_47),
.A2(n_55),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_47),
.A2(n_55),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_47),
.A2(n_55),
.B1(n_203),
.B2(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_47),
.B(n_154),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_51),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_64),
.B(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_67),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_67),
.A2(n_69),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_72),
.A2(n_125),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_72),
.B(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_72),
.A2(n_125),
.B1(n_126),
.B2(n_162),
.Y(n_279)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.C(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_73),
.B(n_102),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_73),
.A2(n_80),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_78),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_78),
.B(n_154),
.CON(n_153),
.SN(n_153)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B(n_101),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_88),
.A2(n_98),
.B1(n_108),
.B2(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_95),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_89),
.A2(n_140),
.B1(n_143),
.B2(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_89),
.A2(n_117),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_89),
.A2(n_94),
.B1(n_236),
.B2(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_90),
.B(n_154),
.Y(n_248)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_96),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_93),
.A2(n_194),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_96),
.A2(n_142),
.B(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_98),
.Y(n_296)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_110),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_105),
.B(n_109),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_110),
.A2(n_111),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.C(n_123),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_112),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_113),
.B(n_118),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_299),
.B(n_304),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_286),
.B(n_298),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_186),
.B(n_267),
.C(n_285),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_174),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_135),
.B(n_174),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_157),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_137),
.B(n_144),
.C(n_157),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_138),
.B(n_139),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_152),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_168),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_159),
.B(n_164),
.C(n_168),
.Y(n_283)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_167),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_171),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_175),
.A2(n_176),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_266),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_259),
.B(n_265),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_214),
.B(n_258),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_205),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_190),
.B(n_205),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_198),
.C(n_201),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_191),
.A2(n_192),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_212),
.C(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_252),
.B(n_257),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_232),
.B(n_251),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_240),
.B(n_250),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_283),
.B2(n_284),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.C(n_284),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_278),
.C(n_281),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.C(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);


endmodule