module fake_jpeg_1489_n_440 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_51),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_59),
.A2(n_21),
.B1(n_29),
.B2(n_15),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_21),
.B(n_1),
.CON(n_70),
.SN(n_70)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_63),
.Y(n_113)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_19),
.B(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_100),
.A2(n_130),
.B1(n_105),
.B2(n_122),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_29),
.B1(n_44),
.B2(n_76),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_105),
.A2(n_120),
.B1(n_122),
.B2(n_23),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_113),
.Y(n_171)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_45),
.A2(n_34),
.B1(n_19),
.B2(n_42),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_36),
.B1(n_35),
.B2(n_22),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_121),
.B1(n_22),
.B2(n_16),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_49),
.A2(n_29),
.B1(n_44),
.B2(n_40),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_37),
.B1(n_34),
.B2(n_24),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_60),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_64),
.A2(n_37),
.B1(n_24),
.B2(n_40),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_52),
.B(n_43),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_67),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_140),
.Y(n_182)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_80),
.B1(n_79),
.B2(n_74),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_144),
.B1(n_148),
.B2(n_170),
.Y(n_184)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_64),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_70),
.B(n_36),
.C(n_35),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_141),
.B(n_145),
.Y(n_206)
);

OR2x2_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_48),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_142),
.B(n_150),
.C(n_156),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_143),
.A2(n_132),
.B1(n_88),
.B2(n_90),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_158),
.Y(n_186)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_91),
.A2(n_69),
.B1(n_62),
.B2(n_58),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_60),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_71),
.B1(n_56),
.B2(n_50),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_161),
.B1(n_119),
.B2(n_131),
.Y(n_183)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_47),
.C(n_46),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_16),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_174),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_98),
.A2(n_129),
.B(n_112),
.C(n_95),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g214 ( 
.A(n_162),
.B(n_2),
.C(n_4),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_8),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_28),
.B1(n_23),
.B2(n_27),
.Y(n_165)
);

OAI22x1_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_1),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_109),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_89),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_97),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_175),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_7),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_176),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_109),
.A2(n_28),
.B1(n_8),
.B2(n_10),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_1),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_97),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_101),
.B1(n_89),
.B2(n_104),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_181),
.A2(n_196),
.B1(n_208),
.B2(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_183),
.A2(n_199),
.B1(n_205),
.B2(n_215),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_101),
.B1(n_131),
.B2(n_133),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_133),
.B1(n_132),
.B2(n_116),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_140),
.B(n_116),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_214),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_162),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_90),
.B1(n_8),
.B2(n_11),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_144),
.A2(n_90),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_219),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_141),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_11),
.B1(n_13),
.B2(n_6),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_5),
.B1(n_6),
.B2(n_184),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_150),
.A2(n_142),
.B1(n_167),
.B2(n_158),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_221),
.B1(n_156),
.B2(n_168),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_6),
.B1(n_2),
.B2(n_5),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_165),
.B(n_160),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_150),
.A2(n_5),
.B1(n_6),
.B2(n_136),
.Y(n_221)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_222),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_150),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_226),
.C(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_155),
.C(n_145),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_146),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_228),
.B(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_186),
.B(n_173),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_206),
.B1(n_184),
.B2(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_163),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_233),
.A2(n_236),
.B(n_242),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_187),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_166),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_147),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_168),
.B1(n_178),
.B2(n_151),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g287 ( 
.A1(n_237),
.A2(n_197),
.B(n_207),
.Y(n_287)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_249),
.Y(n_266)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_139),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_172),
.C(n_153),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_164),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_185),
.B(n_177),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_247),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_187),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_187),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_248),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_203),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_179),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_196),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_183),
.A2(n_178),
.B1(n_154),
.B2(n_175),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_253),
.B1(n_193),
.B2(n_198),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_192),
.B(n_149),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_256),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_199),
.A2(n_154),
.B1(n_157),
.B2(n_169),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_180),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_219),
.B(n_211),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_192),
.B(n_180),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_221),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_137),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_216),
.B1(n_211),
.B2(n_190),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_259),
.B(n_264),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_229),
.A2(n_201),
.B1(n_205),
.B2(n_204),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_293)
);

OAI22x1_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_238),
.B1(n_229),
.B2(n_240),
.Y(n_263)
);

OAI22x1_ASAP7_75t_L g319 ( 
.A1(n_263),
.A2(n_258),
.B1(n_241),
.B2(n_222),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_224),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_191),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_281),
.C(n_289),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_274),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_255),
.B(n_181),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_250),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_232),
.A2(n_231),
.B1(n_244),
.B2(n_235),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_220),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_246),
.A2(n_200),
.B1(n_190),
.B2(n_220),
.Y(n_282)
);

OA21x2_ASAP7_75t_SL g285 ( 
.A1(n_228),
.A2(n_203),
.B(n_195),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_254),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_246),
.A2(n_200),
.B1(n_195),
.B2(n_213),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_286),
.A2(n_251),
.B1(n_253),
.B2(n_234),
.Y(n_313)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_202),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_231),
.A2(n_197),
.B1(n_202),
.B2(n_207),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_237),
.B1(n_248),
.B2(n_247),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_245),
.B(n_242),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_296),
.A2(n_299),
.B(n_303),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_260),
.B(n_230),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_306),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_280),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_309),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_233),
.C(n_223),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_308),
.C(n_315),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_223),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_287),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_249),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_310),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_256),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_312),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_313),
.A2(n_319),
.B1(n_271),
.B2(n_267),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_227),
.B(n_222),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_274),
.B(n_263),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_237),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_282),
.B1(n_287),
.B2(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_241),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_266),
.A2(n_258),
.B1(n_188),
.B2(n_5),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_320),
.A2(n_279),
.B1(n_267),
.B2(n_288),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_285),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_321),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_339),
.B1(n_294),
.B2(n_307),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_340),
.Y(n_368)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_266),
.B(n_289),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_341),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_284),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_317),
.Y(n_334)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_281),
.C(n_259),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_344),
.C(n_345),
.Y(n_351)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_307),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_294),
.B1(n_309),
.B2(n_313),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_308),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_278),
.C(n_270),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_270),
.C(n_264),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_290),
.C(n_272),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_299),
.C(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_349),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_300),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_354),
.A2(n_357),
.B1(n_340),
.B2(n_329),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_358),
.C(n_362),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_326),
.A2(n_293),
.B1(n_307),
.B2(n_299),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_301),
.C(n_304),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_296),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_365),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_297),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_324),
.B(n_306),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_366),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_336),
.B(n_324),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_SL g386 ( 
.A1(n_367),
.A2(n_331),
.A3(n_343),
.B1(n_272),
.B2(n_347),
.C1(n_302),
.C2(n_327),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_331),
.Y(n_374)
);

OAI321xp33_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_333),
.A3(n_325),
.B1(n_336),
.B2(n_338),
.C(n_326),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_374),
.B1(n_383),
.B2(n_387),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_SL g376 ( 
.A(n_361),
.B(n_338),
.C(n_325),
.Y(n_376)
);

OAI221xp5_ASAP7_75t_L g391 ( 
.A1(n_376),
.A2(n_386),
.B1(n_364),
.B2(n_356),
.C(n_352),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_368),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_377),
.B(n_349),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

NAND2xp67_ASAP7_75t_SL g379 ( 
.A(n_359),
.B(n_341),
.Y(n_379)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_330),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_354),
.A2(n_293),
.B1(n_327),
.B2(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_334),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_337),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_322),
.B1(n_332),
.B2(n_342),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_350),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_394),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_384),
.A2(n_368),
.B(n_363),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_381),
.B(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_400),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_365),
.C(n_358),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_393),
.B(n_395),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_348),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_351),
.C(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_397),
.B(n_380),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_399),
.A2(n_401),
.B1(n_387),
.B2(n_339),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_351),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_319),
.B1(n_286),
.B2(n_262),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_375),
.C(n_370),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_405),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_370),
.C(n_383),
.Y(n_405)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_406),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_378),
.C(n_374),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_409),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_355),
.C(n_381),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_382),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_292),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_188),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_413),
.B(n_292),
.Y(n_421)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g416 ( 
.A1(n_410),
.A2(n_376),
.B(n_390),
.C(n_388),
.D(n_398),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_417),
.B(n_420),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_404),
.A2(n_398),
.B(n_411),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_419),
.B(n_408),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_405),
.A2(n_316),
.B1(n_320),
.B2(n_389),
.Y(n_418)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_418),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_407),
.A2(n_409),
.B(n_402),
.Y(n_419)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_420),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_421),
.B(n_403),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_188),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_403),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_425),
.A2(n_426),
.B(n_428),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_430),
.A2(n_419),
.B(n_423),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_433),
.A2(n_434),
.B(n_429),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_425),
.A2(n_414),
.B(n_422),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_436),
.B(n_432),
.Y(n_437)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_431),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_437),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_438),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_439),
.B(n_427),
.Y(n_440)
);


endmodule