module real_aes_7571_n_383 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_383);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_383;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_742;
wire n_766;
wire n_555;
wire n_852;
wire n_974;
wire n_1113;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_889;
wire n_955;
wire n_696;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_1046;
wire n_677;
wire n_948;
wire n_958;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_1140;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_918;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_1098;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_976;
wire n_872;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_780;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_1148;
wire n_409;
wire n_748;
wire n_860;
wire n_909;
wire n_523;
wire n_781;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_504;
wire n_973;
wire n_455;
wire n_725;
wire n_671;
wire n_960;
wire n_1081;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1013;
wire n_1017;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1157;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_385;
wire n_749;
wire n_1056;
wire n_663;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_1155;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_1136;
wire n_720;
wire n_1127;
wire n_968;
wire n_435;
wire n_972;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_1045;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_1156;
wire n_474;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_1097;
wire n_703;
wire n_500;
wire n_601;
wire n_1101;
wire n_1076;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_0), .A2(n_172), .B1(n_665), .B2(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_1), .B(n_454), .Y(n_491) );
XOR2x2_ASAP7_75t_L g397 ( .A(n_2), .B(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_3), .A2(n_299), .B1(n_766), .B2(n_870), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_4), .A2(n_162), .B1(n_453), .B2(n_627), .C(n_1019), .Y(n_1018) );
OA22x2_ASAP7_75t_L g852 ( .A1(n_5), .A2(n_853), .B1(n_854), .B2(n_876), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_5), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_6), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_7), .A2(n_88), .B1(n_700), .B2(n_873), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g1098 ( .A1(n_8), .A2(n_288), .B1(n_528), .B2(n_800), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_9), .A2(n_349), .B1(n_693), .B2(n_702), .Y(n_1000) );
AOI22xp5_ASAP7_75t_SL g664 ( .A1(n_10), .A2(n_379), .B1(n_563), .B2(n_665), .Y(n_664) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_11), .A2(n_217), .B1(n_407), .B2(n_412), .Y(n_416) );
INVx1_ASAP7_75t_L g1123 ( .A(n_11), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_12), .Y(n_894) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_13), .A2(n_61), .B1(n_322), .B2(n_586), .C1(n_588), .C2(n_589), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_14), .A2(n_301), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_15), .A2(n_66), .B1(n_717), .B2(n_1076), .Y(n_1075) );
AOI22xp5_ASAP7_75t_SL g657 ( .A1(n_16), .A2(n_243), .B1(n_658), .B2(n_659), .Y(n_657) );
AO22x1_ASAP7_75t_L g812 ( .A1(n_17), .A2(n_813), .B1(n_844), .B2(n_845), .Y(n_812) );
INVx1_ASAP7_75t_L g844 ( .A(n_17), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_18), .A2(n_104), .B1(n_567), .B2(n_898), .Y(n_1084) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_19), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_20), .A2(n_25), .B1(n_720), .B2(n_800), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_21), .A2(n_382), .B1(n_445), .B2(n_706), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_22), .A2(n_375), .B1(n_769), .B2(n_833), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g1106 ( .A(n_23), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_24), .A2(n_370), .B1(n_434), .B2(n_436), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_26), .A2(n_263), .B1(n_497), .B2(n_499), .Y(n_1105) );
INVx1_ASAP7_75t_L g467 ( .A(n_27), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_28), .A2(n_246), .B1(n_453), .B2(n_579), .C(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_29), .A2(n_363), .B1(n_434), .B2(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_30), .A2(n_174), .B1(n_456), .B2(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_31), .A2(n_337), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_32), .A2(n_97), .B1(n_469), .B2(n_473), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_33), .A2(n_598), .B1(n_638), .B2(n_639), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_33), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_34), .A2(n_559), .B1(n_590), .B2(n_591), .Y(n_558) );
INVx1_ASAP7_75t_L g590 ( .A(n_34), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_35), .A2(n_57), .B1(n_732), .B2(n_1087), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_36), .Y(n_865) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_37), .A2(n_109), .B1(n_407), .B2(n_408), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_38), .A2(n_256), .B1(n_543), .B2(n_727), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_39), .A2(n_101), .B1(n_588), .B2(n_717), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_40), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_41), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_42), .A2(n_250), .B1(n_628), .B2(n_794), .Y(n_1137) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_43), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g1136 ( .A1(n_44), .A2(n_331), .B1(n_487), .B2(n_1036), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_45), .A2(n_326), .B1(n_548), .B2(n_697), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g1133 ( .A(n_46), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_47), .B(n_794), .Y(n_1079) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_48), .A2(n_275), .B1(n_403), .B2(n_662), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_49), .A2(n_227), .B1(n_702), .B2(n_843), .Y(n_842) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_50), .A2(n_144), .B1(n_295), .B2(n_589), .C1(n_635), .C2(n_637), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_51), .B(n_527), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_52), .A2(n_268), .B1(n_526), .B2(n_527), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_53), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_54), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_55), .A2(n_193), .B1(n_527), .B2(n_648), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_56), .A2(n_140), .B1(n_427), .B2(n_659), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_58), .B(n_465), .Y(n_892) );
AOI222xp33_ASAP7_75t_L g1022 ( .A1(n_59), .A2(n_208), .B1(n_315), .B2(n_586), .C1(n_648), .C2(n_716), .Y(n_1022) );
CKINVDCx20_ASAP7_75t_R g977 ( .A(n_60), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_62), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_63), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_64), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_65), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_67), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_68), .A2(n_364), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_69), .A2(n_297), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_70), .A2(n_201), .B1(n_616), .B2(n_705), .Y(n_991) );
INVx1_ASAP7_75t_L g668 ( .A(n_71), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_72), .A2(n_106), .B1(n_836), .B2(n_837), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_73), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_74), .A2(n_202), .B1(n_460), .B2(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_75), .A2(n_269), .B1(n_436), .B2(n_667), .Y(n_809) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_76), .A2(n_77), .B1(n_611), .B2(n_1142), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_78), .A2(n_143), .B1(n_401), .B2(n_496), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_79), .A2(n_251), .B1(n_457), .B2(n_470), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_80), .A2(n_231), .B1(n_840), .B2(n_898), .Y(n_927) );
AOI22xp33_ASAP7_75t_SL g1139 ( .A1(n_81), .A2(n_238), .B1(n_904), .B2(n_1140), .Y(n_1139) );
AOI22xp5_ASAP7_75t_SL g660 ( .A1(n_82), .A2(n_249), .B1(n_427), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g1080 ( .A1(n_83), .A2(n_223), .B1(n_469), .B2(n_957), .Y(n_1080) );
CKINVDCx20_ASAP7_75t_R g976 ( .A(n_84), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g1156 ( .A(n_85), .Y(n_1156) );
OA22x2_ASAP7_75t_L g1157 ( .A1(n_85), .A2(n_1129), .B1(n_1156), .B2(n_1158), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_86), .A2(n_247), .B1(n_436), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_87), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_89), .A2(n_281), .B1(n_496), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_90), .A2(n_213), .B1(n_548), .B2(n_550), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_91), .Y(n_1097) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_92), .A2(n_255), .B1(n_407), .B2(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g1120 ( .A(n_92), .Y(n_1120) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_93), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_94), .A2(n_99), .B1(n_543), .B2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_95), .A2(n_182), .B1(n_800), .B2(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_96), .A2(n_316), .B1(n_553), .B2(n_603), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_98), .Y(n_614) );
AOI22xp5_ASAP7_75t_SL g666 ( .A1(n_100), .A2(n_206), .B1(n_616), .B2(n_667), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g1041 ( .A1(n_102), .A2(n_658), .B(n_1042), .C(n_1045), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_103), .A2(n_285), .B1(n_487), .B2(n_1036), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_105), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_107), .A2(n_114), .B1(n_919), .B2(n_920), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_108), .A2(n_176), .B1(n_457), .B2(n_637), .Y(n_1060) );
INVx1_ASAP7_75t_L g1124 ( .A(n_109), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_110), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_111), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_112), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_113), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_115), .A2(n_196), .B1(n_807), .B2(n_808), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_116), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_117), .A2(n_354), .B1(n_693), .B2(n_904), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_118), .B(n_628), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_119), .A2(n_329), .B1(n_496), .B2(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_120), .A2(n_204), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_121), .A2(n_360), .B1(n_543), .B2(n_705), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_122), .A2(n_239), .B1(n_616), .B2(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_123), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g1145 ( .A1(n_124), .A2(n_272), .B1(n_497), .B2(n_1146), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_125), .A2(n_137), .B1(n_486), .B2(n_526), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_126), .A2(n_185), .B1(n_417), .B2(n_727), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_127), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_128), .A2(n_333), .B1(n_732), .B2(n_766), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_129), .A2(n_240), .B1(n_457), .B2(n_469), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_130), .A2(n_367), .B1(n_771), .B2(n_773), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_131), .A2(n_343), .B1(n_486), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_132), .A2(n_151), .B1(n_603), .B2(n_898), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_133), .A2(n_188), .B1(n_628), .B2(n_629), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_134), .A2(n_361), .B1(n_702), .B2(n_705), .Y(n_701) );
XNOR2x2_ASAP7_75t_L g994 ( .A(n_135), .B(n_995), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_136), .A2(n_149), .B1(n_603), .B2(n_840), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_138), .A2(n_209), .B1(n_543), .B2(n_561), .C(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g510 ( .A(n_139), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_141), .B(n_454), .Y(n_1101) );
AND2x6_ASAP7_75t_L g386 ( .A(n_142), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_142), .Y(n_1117) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_145), .A2(n_369), .B1(n_445), .B2(n_563), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_146), .A2(n_186), .B1(n_504), .B2(n_808), .Y(n_992) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_147), .B(n_627), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_148), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_150), .A2(n_350), .B1(n_436), .B2(n_904), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_152), .A2(n_190), .B1(n_401), .B2(n_417), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_153), .B(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_154), .A2(n_267), .B1(n_715), .B2(n_716), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_155), .Y(n_601) );
AO22x1_ASAP7_75t_L g1006 ( .A1(n_156), .A2(n_1007), .B1(n_1023), .B2(n_1024), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_156), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_157), .A2(n_177), .B1(n_504), .B2(n_1063), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_158), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_159), .B(n_490), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_160), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g1005 ( .A1(n_161), .A2(n_203), .B1(n_338), .B2(n_465), .C1(n_589), .C2(n_715), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_163), .A2(n_304), .B1(n_840), .B2(n_841), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_164), .A2(n_232), .B1(n_628), .B2(n_794), .Y(n_1037) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_165), .A2(n_248), .B1(n_407), .B2(n_408), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_165), .B(n_1122), .Y(n_1121) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_166), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g1046 ( .A(n_167), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_168), .A2(n_291), .B1(n_438), .B2(n_704), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_169), .A2(n_195), .B1(n_401), .B2(n_545), .C(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_170), .A2(n_180), .B1(n_556), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g1039 ( .A1(n_171), .A2(n_266), .B1(n_773), .B2(n_904), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_173), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_175), .A2(n_199), .B1(n_436), .B2(n_504), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_178), .A2(n_257), .B1(n_499), .B2(n_732), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_179), .A2(n_187), .B1(n_629), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_181), .A2(n_325), .B1(n_695), .B2(n_697), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_183), .A2(n_314), .B1(n_705), .B2(n_769), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_184), .A2(n_198), .B1(n_434), .B2(n_545), .C(n_1009), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_189), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_191), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_192), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_194), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_197), .A2(n_300), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g1126 ( .A1(n_200), .A2(n_1127), .B1(n_1128), .B2(n_1148), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_200), .Y(n_1148) );
XNOR2xp5_ASAP7_75t_L g1028 ( .A(n_205), .B(n_1029), .Y(n_1028) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_207), .A2(n_237), .B1(n_659), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_210), .A2(n_230), .B1(n_427), .B2(n_505), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_211), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_212), .A2(n_235), .B1(n_445), .B2(n_1013), .C(n_1014), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_214), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_215), .A2(n_334), .B1(n_697), .B2(n_946), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_216), .A2(n_236), .B1(n_442), .B2(n_445), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_218), .B(n_627), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g942 ( .A(n_219), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_220), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_221), .A2(n_262), .B1(n_507), .B2(n_508), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_222), .A2(n_274), .B1(n_748), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_224), .A2(n_306), .B1(n_766), .B2(n_836), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_225), .B(n_697), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_226), .Y(n_980) );
OA22x2_ASAP7_75t_L g882 ( .A1(n_228), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_228), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_229), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_233), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_234), .A2(n_327), .B1(n_545), .B2(n_843), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_241), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_242), .Y(n_646) );
INVx2_ASAP7_75t_L g391 ( .A(n_244), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_245), .A2(n_296), .B1(n_496), .B2(n_508), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_252), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_253), .Y(n_752) );
XNOR2x1_ASAP7_75t_L g1070 ( .A(n_254), .B(n_1071), .Y(n_1070) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_258), .A2(n_939), .B1(n_964), .B2(n_965), .Y(n_938) );
INVx1_ASAP7_75t_L g964 ( .A(n_258), .Y(n_964) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_259), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_260), .Y(n_888) );
AOI211xp5_ASAP7_75t_L g383 ( .A1(n_261), .A2(n_384), .B(n_392), .C(n_1125), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_264), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_265), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_270), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g955 ( .A(n_271), .Y(n_955) );
OA22x2_ASAP7_75t_L g707 ( .A1(n_273), .A2(n_708), .B1(n_709), .B2(n_733), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_273), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_276), .A2(n_294), .B1(n_500), .B2(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_277), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_278), .Y(n_914) );
AOI22x1_ASAP7_75t_L g742 ( .A1(n_279), .A2(n_743), .B1(n_774), .B2(n_775), .Y(n_742) );
INVx1_ASAP7_75t_L g774 ( .A(n_279), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_280), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g983 ( .A(n_282), .Y(n_983) );
OA22x2_ASAP7_75t_L g906 ( .A1(n_283), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_906) );
CKINVDCx16_ASAP7_75t_R g907 ( .A(n_283), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_284), .A2(n_351), .B1(n_424), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g407 ( .A(n_286), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_286), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_287), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_289), .A2(n_335), .B1(n_836), .B2(n_929), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g1132 ( .A(n_290), .Y(n_1132) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_292), .A2(n_380), .B1(n_627), .B2(n_629), .C(n_631), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_293), .A2(n_328), .B1(n_504), .B2(n_505), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g935 ( .A(n_298), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_302), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_303), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_305), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_307), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_308), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_309), .A2(n_784), .B1(n_785), .B2(n_810), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_309), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_310), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g1134 ( .A(n_311), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_312), .A2(n_358), .B1(n_456), .B2(n_460), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g1065 ( .A(n_313), .Y(n_1065) );
AND2x2_ASAP7_75t_L g390 ( .A(n_317), .B(n_391), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_318), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_319), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_320), .Y(n_979) );
INVx1_ASAP7_75t_L g387 ( .A(n_321), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_323), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_324), .Y(n_515) );
XOR2x2_ASAP7_75t_L g972 ( .A(n_330), .B(n_973), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_332), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_336), .B(n_450), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_339), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_340), .A2(n_374), .B1(n_528), .B2(n_800), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_341), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_342), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g1074 ( .A(n_344), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_345), .B(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_346), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_347), .A2(n_381), .B1(n_450), .B2(n_453), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_348), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_352), .A2(n_362), .B1(n_567), .B2(n_667), .Y(n_1001) );
XNOR2x1_ASAP7_75t_L g511 ( .A(n_353), .B(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_355), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_356), .A2(n_376), .B1(n_697), .B2(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_357), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_359), .B(n_454), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_365), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_366), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_368), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_371), .B(n_526), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_372), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_373), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_377), .B(n_652), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_378), .Y(n_828) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_387), .Y(n_1116) );
OAI21xp5_ASAP7_75t_L g1154 ( .A1(n_388), .A2(n_1115), .B(n_1155), .Y(n_1154) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_848), .B1(n_1110), .B2(n_1111), .C(n_1112), .Y(n_392) );
INVx1_ASAP7_75t_L g1111 ( .A(n_393), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_593), .B1(n_846), .B2(n_847), .Y(n_393) );
INVx1_ASAP7_75t_L g847 ( .A(n_394), .Y(n_847) );
OAI22xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_557), .B1(n_558), .B2(n_592), .Y(n_394) );
INVx1_ASAP7_75t_L g592 ( .A(n_395), .Y(n_592) );
AO22x1_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_475), .B2(n_476), .Y(n_395) );
AO22x1_ASAP7_75t_L g781 ( .A1(n_396), .A2(n_397), .B1(n_782), .B2(n_783), .Y(n_781) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
NOR4xp75_ASAP7_75t_L g398 ( .A(n_399), .B(n_432), .C(n_448), .D(n_463), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_400), .B(n_423), .Y(n_399) );
INVx2_ASAP7_75t_L g618 ( .A(n_401), .Y(n_618) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g667 ( .A(n_402), .Y(n_667) );
INVx2_ASAP7_75t_L g841 ( .A(n_402), .Y(n_841) );
INVx3_ASAP7_75t_L g1087 ( .A(n_402), .Y(n_1087) );
INVx6_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx3_ASAP7_75t_L g504 ( .A(n_403), .Y(n_504) );
BUFx3_ASAP7_75t_L g556 ( .A(n_403), .Y(n_556) );
BUFx3_ASAP7_75t_L g904 ( .A(n_403), .Y(n_904) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_413), .Y(n_403) );
AND2x2_ASAP7_75t_L g435 ( .A(n_404), .B(n_421), .Y(n_435) );
AND2x6_ASAP7_75t_L g438 ( .A(n_404), .B(n_439), .Y(n_438) );
AND2x6_ASAP7_75t_L g466 ( .A(n_404), .B(n_462), .Y(n_466) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_410), .Y(n_404) );
AND2x2_ASAP7_75t_L g444 ( .A(n_405), .B(n_411), .Y(n_444) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g419 ( .A(n_406), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_406), .B(n_411), .Y(n_431) );
AND2x2_ASAP7_75t_L g459 ( .A(n_406), .B(n_416), .Y(n_459) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_409), .Y(n_412) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g420 ( .A(n_411), .Y(n_420) );
INVx1_ASAP7_75t_L g472 ( .A(n_411), .Y(n_472) );
AND2x2_ASAP7_75t_L g426 ( .A(n_413), .B(n_419), .Y(n_426) );
AND2x6_ASAP7_75t_L g454 ( .A(n_413), .B(n_444), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_413), .B(n_444), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_413), .B(n_419), .Y(n_574) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g422 ( .A(n_414), .Y(n_422) );
INVx1_ASAP7_75t_L g430 ( .A(n_414), .Y(n_430) );
OR2x2_ASAP7_75t_L g440 ( .A(n_414), .B(n_415), .Y(n_440) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_416), .Y(n_462) );
AND2x2_ASAP7_75t_L g421 ( .A(n_415), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g1140 ( .A(n_417), .Y(n_1140) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
BUFx3_ASAP7_75t_L g563 ( .A(n_418), .Y(n_563) );
BUFx3_ASAP7_75t_L g704 ( .A(n_418), .Y(n_704) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_419), .B(n_421), .Y(n_625) );
INVx1_ASAP7_75t_L g461 ( .A(n_420), .Y(n_461) );
AND2x4_ASAP7_75t_L g443 ( .A(n_421), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g446 ( .A(n_421), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g471 ( .A(n_422), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g509 ( .A(n_422), .Y(n_509) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_424), .Y(n_946) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx5_ASAP7_75t_L g505 ( .A(n_425), .Y(n_505) );
BUFx3_ASAP7_75t_L g549 ( .A(n_425), .Y(n_549) );
INVx4_ASAP7_75t_L g662 ( .A(n_425), .Y(n_662) );
INVx3_ASAP7_75t_L g732 ( .A(n_425), .Y(n_732) );
INVx1_ASAP7_75t_L g1143 ( .A(n_425), .Y(n_1143) );
INVx8_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g577 ( .A(n_428), .Y(n_577) );
BUFx2_ASAP7_75t_L g611 ( .A(n_428), .Y(n_611) );
BUFx4f_ASAP7_75t_SL g837 ( .A(n_428), .Y(n_837) );
BUFx2_ASAP7_75t_L g929 ( .A(n_428), .Y(n_929) );
INVx6_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g550 ( .A(n_429), .Y(n_550) );
INVx1_ASAP7_75t_SL g697 ( .A(n_429), .Y(n_697) );
INVx1_ASAP7_75t_L g766 ( .A(n_429), .Y(n_766) );
OR2x6_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
INVx1_ASAP7_75t_L g447 ( .A(n_431), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_433), .B(n_441), .Y(n_432) );
INVx1_ASAP7_75t_L g621 ( .A(n_434), .Y(n_621) );
BUFx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_435), .Y(n_499) );
BUFx2_ASAP7_75t_SL g658 ( .A(n_435), .Y(n_658) );
INVx2_ASAP7_75t_L g899 ( .A(n_435), .Y(n_899) );
INVx4_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g616 ( .A(n_437), .Y(n_616) );
INVx4_ASAP7_75t_L g873 ( .A(n_437), .Y(n_873) );
INVx3_ASAP7_75t_L g1013 ( .A(n_437), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_437), .B(n_1046), .Y(n_1045) );
INVx11_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx11_ASAP7_75t_L g501 ( .A(n_438), .Y(n_501) );
AND2x4_ASAP7_75t_L g452 ( .A(n_439), .B(n_444), .Y(n_452) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g517 ( .A(n_440), .B(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g603 ( .A(n_442), .Y(n_603) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_443), .Y(n_507) );
BUFx3_ASAP7_75t_L g659 ( .A(n_443), .Y(n_659) );
BUFx3_ASAP7_75t_L g706 ( .A(n_443), .Y(n_706) );
INVx2_ASAP7_75t_L g834 ( .A(n_443), .Y(n_834) );
INVx1_ASAP7_75t_L g518 ( .A(n_444), .Y(n_518) );
INVx1_ASAP7_75t_L g569 ( .A(n_445), .Y(n_569) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
INVx1_ASAP7_75t_L g554 ( .A(n_446), .Y(n_554) );
BUFx3_ASAP7_75t_L g606 ( .A(n_446), .Y(n_606) );
BUFx2_ASAP7_75t_L g665 ( .A(n_446), .Y(n_665) );
BUFx2_ASAP7_75t_SL g700 ( .A(n_446), .Y(n_700) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_446), .Y(n_727) );
BUFx3_ASAP7_75t_L g843 ( .A(n_446), .Y(n_843) );
AND2x2_ASAP7_75t_L g508 ( .A(n_447), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_449), .B(n_455), .Y(n_448) );
BUFx2_ASAP7_75t_L g579 ( .A(n_450), .Y(n_579) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
INVx5_ASAP7_75t_L g628 ( .A(n_451), .Y(n_628) );
INVx2_ASAP7_75t_L g723 ( .A(n_451), .Y(n_723) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx4f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g630 ( .A(n_454), .Y(n_630) );
BUFx2_ASAP7_75t_L g794 ( .A(n_454), .Y(n_794) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g721 ( .A(n_457), .Y(n_721) );
BUFx2_ASAP7_75t_L g957 ( .A(n_457), .Y(n_957) );
BUFx2_ASAP7_75t_L g1036 ( .A(n_457), .Y(n_1036) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AND2x4_ASAP7_75t_L g470 ( .A(n_459), .B(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g473 ( .A(n_459), .B(n_474), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_459), .B(n_509), .Y(n_533) );
BUFx3_ASAP7_75t_L g487 ( .A(n_460), .Y(n_487) );
BUFx2_ASAP7_75t_SL g655 ( .A(n_460), .Y(n_655) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_460), .Y(n_800) );
BUFx2_ASAP7_75t_SL g1076 ( .A(n_460), .Y(n_1076) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
INVx1_ASAP7_75t_L g538 ( .A(n_462), .Y(n_538) );
OAI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_467), .B(n_468), .Y(n_463) );
OAI21xp33_ASAP7_75t_SL g916 ( .A1(n_464), .A2(n_917), .B(n_918), .Y(n_916) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g484 ( .A(n_466), .Y(n_484) );
INVx4_ASAP7_75t_L g587 ( .A(n_466), .Y(n_587) );
INVx2_ASAP7_75t_SL g681 ( .A(n_466), .Y(n_681) );
INVx2_ASAP7_75t_L g712 ( .A(n_466), .Y(n_712) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_466), .Y(n_789) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_469), .Y(n_588) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_470), .Y(n_526) );
BUFx4f_ASAP7_75t_SL g637 ( .A(n_470), .Y(n_637) );
BUFx2_ASAP7_75t_L g715 ( .A(n_470), .Y(n_715) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_470), .Y(n_748) );
INVx1_ASAP7_75t_L g474 ( .A(n_472), .Y(n_474) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_473), .Y(n_486) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_473), .Y(n_528) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_473), .Y(n_717) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
XNOR2x1_ASAP7_75t_SL g476 ( .A(n_477), .B(n_511), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_477), .A2(n_742), .B1(n_776), .B2(n_777), .Y(n_741) );
INVx1_ASAP7_75t_L g776 ( .A(n_477), .Y(n_776) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
XOR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_510), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_481), .B(n_493), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_488), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_485), .Y(n_482) );
OAI21xp33_ASAP7_75t_SL g523 ( .A1(n_484), .A2(n_524), .B(n_525), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_484), .A2(n_746), .B1(n_747), .B2(n_749), .C(n_750), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g859 ( .A1(n_484), .A2(n_860), .B(n_861), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g978 ( .A1(n_484), .A2(n_825), .B1(n_979), .B2(n_980), .C(n_981), .Y(n_978) );
BUFx4f_ASAP7_75t_SL g589 ( .A(n_486), .Y(n_589) );
INVx2_ASAP7_75t_L g921 ( .A(n_486), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .C(n_492), .Y(n_488) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx2_ASAP7_75t_L g763 ( .A(n_497), .Y(n_763) );
INVx3_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
BUFx3_ASAP7_75t_L g693 ( .A(n_499), .Y(n_693) );
BUFx3_ASAP7_75t_L g769 ( .A(n_499), .Y(n_769) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_499), .Y(n_807) );
INVx5_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g567 ( .A(n_501), .Y(n_567) );
INVx2_ASAP7_75t_L g840 ( .A(n_501), .Y(n_840) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_501), .Y(n_1063) );
INVx1_ASAP7_75t_L g1146 ( .A(n_501), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_505), .Y(n_765) );
BUFx2_ASAP7_75t_L g870 ( .A(n_505), .Y(n_870) );
INVx4_ASAP7_75t_L g546 ( .A(n_507), .Y(n_546) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_540), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .C(n_529), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_519), .B2(n_520), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_516), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_516), .A2(n_521), .B1(n_888), .B2(n_889), .Y(n_887) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_517), .Y(n_675) );
INVx2_ASAP7_75t_L g818 ( .A(n_517), .Y(n_818) );
OAI22xp5_ASAP7_75t_SL g911 ( .A1(n_520), .A2(n_912), .B1(n_914), .B2(n_915), .Y(n_911) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g674 ( .A1(n_521), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g954 ( .A(n_521), .Y(n_954) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g755 ( .A(n_522), .Y(n_755) );
INVx4_ASAP7_75t_L g649 ( .A(n_526), .Y(n_649) );
BUFx2_ASAP7_75t_L g919 ( .A(n_526), .Y(n_919) );
INVx1_ASAP7_75t_L g683 ( .A(n_527), .Y(n_683) );
BUFx4f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_534), .B2(n_535), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_531), .A2(n_535), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx3_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g582 ( .A(n_532), .Y(n_582) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g686 ( .A(n_533), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_533), .A2(n_535), .B1(n_857), .B2(n_858), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_533), .A2(n_537), .B1(n_894), .B2(n_895), .Y(n_893) );
OAI22xp33_ASAP7_75t_SL g922 ( .A1(n_533), .A2(n_688), .B1(n_923), .B2(n_924), .Y(n_922) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_533), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_535), .A2(n_686), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g688 ( .A(n_536), .Y(n_688) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g584 ( .A(n_537), .Y(n_584) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_551), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_547), .Y(n_541) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g803 ( .A(n_546), .Y(n_803) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_554), .A2(n_935), .B1(n_936), .B2(n_937), .Y(n_934) );
INVx1_ASAP7_75t_L g772 ( .A(n_556), .Y(n_772) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
AND4x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_570), .C(n_578), .D(n_585), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g773 ( .A(n_563), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_568), .B2(n_569), .Y(n_564) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_575), .B2(n_576), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_573), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_573), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
OAI21xp33_ASAP7_75t_L g1042 ( .A1(n_573), .A2(n_1043), .B(n_1044), .Y(n_1042) );
BUFx2_ASAP7_75t_R g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_583), .B2(n_584), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_582), .A2(n_584), .B1(n_632), .B2(n_633), .Y(n_631) );
INVx4_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g636 ( .A(n_587), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_587), .A2(n_646), .B(n_647), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g1054 ( .A1(n_587), .A2(n_1055), .B(n_1056), .Y(n_1054) );
OAI21xp5_ASAP7_75t_SL g1073 ( .A1(n_587), .A2(n_1074), .B(n_1075), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g1096 ( .A1(n_587), .A2(n_1097), .B(n_1098), .Y(n_1096) );
INVx2_ASAP7_75t_SL g679 ( .A(n_588), .Y(n_679) );
INVx1_ASAP7_75t_L g846 ( .A(n_593), .Y(n_846) );
XNOR2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_738), .Y(n_593) );
XOR2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_640), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g639 ( .A(n_598), .Y(n_639) );
AND4x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_612), .C(n_626), .D(n_634), .Y(n_598) );
NOR2xp33_ASAP7_75t_SL g599 ( .A(n_600), .B(n_607), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_619), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_618), .A2(n_931), .B1(n_932), .B2(n_933), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_618), .A2(n_623), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g941 ( .A1(n_623), .A2(n_942), .B1(n_943), .B2(n_944), .C(n_945), .Y(n_941) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g933 ( .A(n_624), .Y(n_933) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g652 ( .A(n_630), .Y(n_652) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI222xp33_ASAP7_75t_L g1131 ( .A1(n_636), .A2(n_683), .B1(n_747), .B2(n_1132), .C1(n_1133), .C2(n_1134), .Y(n_1131) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_669), .B1(n_736), .B2(n_737), .Y(n_640) );
INVx2_ASAP7_75t_L g737 ( .A(n_641), .Y(n_737) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
XOR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_668), .Y(n_642) );
NAND3x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_656), .C(n_663), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_650), .Y(n_644) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .C(n_654), .Y(n_650) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g936 ( .A(n_659), .Y(n_936) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g696 ( .A(n_662), .Y(n_696) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_662), .Y(n_836) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g736 ( .A(n_669), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_707), .B1(n_734), .B2(n_735), .Y(n_669) );
INVx2_ASAP7_75t_L g734 ( .A(n_670), .Y(n_734) );
XNOR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_690), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_678), .C(n_685), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_675), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g913 ( .A(n_675), .Y(n_913) );
OAI221xp5_ASAP7_75t_SL g951 ( .A1(n_675), .A2(n_952), .B1(n_953), .B2(n_955), .C(n_956), .Y(n_951) );
OAI222xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_681), .B2(n_682), .C1(n_683), .C2(n_684), .Y(n_678) );
OAI22xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_686), .A2(n_688), .B1(n_828), .B2(n_829), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_688), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_698), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx3_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g943 ( .A(n_700), .Y(n_943) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx4f_ASAP7_75t_SL g808 ( .A(n_704), .Y(n_808) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g735 ( .A(n_707), .Y(n_735) );
INVx2_ASAP7_75t_L g733 ( .A(n_709), .Y(n_733) );
NAND2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_724), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_718), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_713), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g821 ( .A(n_715), .Y(n_821) );
INVx2_ASAP7_75t_L g825 ( .A(n_716), .Y(n_825) );
BUFx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g863 ( .A(n_717), .Y(n_863) );
BUFx2_ASAP7_75t_L g962 ( .A(n_717), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g797 ( .A(n_721), .Y(n_797) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_729), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
XNOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_778), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g777 ( .A(n_742), .Y(n_777) );
INVx2_ASAP7_75t_SL g775 ( .A(n_743), .Y(n_775) );
AND2x4_ASAP7_75t_L g743 ( .A(n_744), .B(n_759), .Y(n_743) );
NOR3xp33_ASAP7_75t_SL g744 ( .A(n_745), .B(n_751), .C(n_756), .Y(n_744) );
OAI222xp33_ASAP7_75t_L g958 ( .A1(n_747), .A2(n_823), .B1(n_959), .B2(n_960), .C1(n_961), .C2(n_963), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_754), .A2(n_816), .B1(n_817), .B2(n_819), .Y(n_815) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g867 ( .A(n_755), .Y(n_867) );
NOR2x1_ASAP7_75t_L g759 ( .A(n_760), .B(n_767), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_764), .Y(n_760) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
BUFx3_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_811), .B2(n_812), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g810 ( .A(n_785), .Y(n_810) );
NAND3x1_ASAP7_75t_L g785 ( .A(n_786), .B(n_801), .C(n_805), .Y(n_785) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_787), .B(n_792), .Y(n_786) );
OAI21xp5_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_790), .B(n_791), .Y(n_787) );
OAI21xp5_ASAP7_75t_SL g1031 ( .A1(n_788), .A2(n_1032), .B(n_1033), .Y(n_1031) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_SL g823 ( .A(n_789), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .C(n_796), .Y(n_792) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_804), .Y(n_801) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_SL g845 ( .A(n_813), .Y(n_845) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_830), .Y(n_813) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_820), .C(n_827), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_817), .A2(n_953), .B1(n_976), .B2(n_977), .Y(n_975) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI222xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_824), .C1(n_825), .C2(n_826), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_838), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_L g875 ( .A(n_834), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_837), .Y(n_1017) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_839), .B(n_842), .Y(n_838) );
INVxp67_ASAP7_75t_L g1110 ( .A(n_848), .Y(n_1110) );
XOR2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_1025), .Y(n_848) );
OAI22xp5_ASAP7_75t_SL g849 ( .A1(n_850), .A2(n_851), .B1(n_968), .B2(n_969), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AOI22x1_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_877), .B1(n_878), .B2(n_967), .Y(n_851) );
INVx1_ASAP7_75t_L g967 ( .A(n_852), .Y(n_967) );
INVx2_ASAP7_75t_L g876 ( .A(n_854), .Y(n_876) );
NAND2x1_ASAP7_75t_L g854 ( .A(n_855), .B(n_868), .Y(n_854) );
NOR3xp33_ASAP7_75t_SL g855 ( .A(n_856), .B(n_859), .C(n_864), .Y(n_855) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
AND4x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_871), .C(n_872), .D(n_874), .Y(n_868) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AO22x2_ASAP7_75t_SL g878 ( .A1(n_879), .A2(n_880), .B1(n_938), .B2(n_966), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_905), .B2(n_906), .Y(n_880) );
INVx2_ASAP7_75t_SL g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
AND3x1_ASAP7_75t_L g885 ( .A(n_886), .B(n_896), .C(n_901), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_890), .C(n_893), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .Y(n_896) );
INVx3_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
XNOR2x2_ASAP7_75t_L g1068 ( .A(n_906), .B(n_1069), .Y(n_1068) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_910), .B(n_925), .Y(n_909) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_916), .C(n_922), .Y(n_910) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx3_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NOR3xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_930), .C(n_934), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
INVx2_ASAP7_75t_L g966 ( .A(n_938), .Y(n_966) );
INVx1_ASAP7_75t_L g965 ( .A(n_939), .Y(n_965) );
AND2x2_ASAP7_75t_SL g939 ( .A(n_940), .B(n_950), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_947), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .Y(n_947) );
NOR2xp33_ASAP7_75t_SL g950 ( .A(n_951), .B(n_958), .Y(n_950) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVxp67_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
XOR2x2_ASAP7_75t_L g969 ( .A(n_970), .B(n_1006), .Y(n_969) );
OAI22xp5_ASAP7_75t_SL g970 ( .A1(n_971), .A2(n_972), .B1(n_993), .B2(n_994), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_986), .Y(n_973) );
NOR3xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_978), .C(n_982), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_990), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NAND4xp75_ASAP7_75t_L g995 ( .A(n_996), .B(n_999), .C(n_1002), .D(n_1005), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
AND2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
AND2x2_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1004), .Y(n_1002) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1007), .Y(n_1024) );
AND4x1_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1012), .C(n_1018), .D(n_1022), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1068), .B1(n_1108), .B2(n_1109), .Y(n_1025) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1026), .Y(n_1108) );
INVx1_ASAP7_75t_SL g1026 ( .A(n_1027), .Y(n_1026) );
OAI22x1_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1047), .B1(n_1066), .B2(n_1067), .Y(n_1027) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1028), .Y(n_1066) );
NAND3x1_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1038), .C(n_1041), .Y(n_1029) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1034), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1037), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1047), .Y(n_1067) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
XOR2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1065), .Y(n_1048) );
NAND3x1_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1053), .C(n_1061), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
NOR2x1_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1057), .Y(n_1053) );
NAND3xp33_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1059), .C(n_1060), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1064), .Y(n_1061) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1068), .Y(n_1109) );
OAI22x1_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1089), .B1(n_1090), .B2(n_1107), .Y(n_1069) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1070), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1081), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1077), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1079), .C(n_1080), .Y(n_1077) );
NOR2x1_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1085), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .Y(n_1085) );
INVx3_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
XOR2x2_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1106), .Y(n_1090) );
NAND3x1_ASAP7_75t_SL g1091 ( .A(n_1092), .B(n_1095), .C(n_1103), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .Y(n_1092) );
NOR2x1_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1099), .Y(n_1095) );
NAND3xp33_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1101), .C(n_1102), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
NOR2x1_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1118), .Y(n_1113) );
OR2x2_ASAP7_75t_SL g1161 ( .A(n_1114), .B(n_1119), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1117), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OAI322xp33_ASAP7_75t_L g1125 ( .A1(n_1116), .A2(n_1126), .A3(n_1149), .B1(n_1153), .B2(n_1156), .C1(n_1157), .C2(n_1159), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1116), .B(n_1152), .Y(n_1155) );
CKINVDCx16_ASAP7_75t_R g1152 ( .A(n_1117), .Y(n_1152) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_1119), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1124), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g1127 ( .A(n_1128), .Y(n_1127) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1129), .Y(n_1158) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1138), .C(n_1144), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1135), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1141), .Y(n_1138) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1147), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
CKINVDCx20_ASAP7_75t_R g1153 ( .A(n_1154), .Y(n_1153) );
CKINVDCx20_ASAP7_75t_R g1159 ( .A(n_1160), .Y(n_1159) );
CKINVDCx20_ASAP7_75t_R g1160 ( .A(n_1161), .Y(n_1160) );
endmodule