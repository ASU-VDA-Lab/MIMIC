module real_jpeg_25837_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_288;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx3_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_2),
.B(n_79),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_42),
.C(n_56),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_180),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_153),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_180),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_2),
.B(n_28),
.C(n_47),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_2),
.A2(n_30),
.B(n_241),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g76 ( 
.A(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_68),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_68),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_8),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_8),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_84),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_211)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_10),
.A2(n_29),
.B1(n_41),
.B2(n_42),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_11),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_63),
.B1(n_83),
.B2(n_110),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_63),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_14),
.A2(n_85),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_14),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_133),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_133),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_15),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_95)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_16),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_20),
.B(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_113),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_65),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_25),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_26),
.A2(n_30),
.B1(n_101),
.B2(n_122),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_27),
.B(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_30),
.A2(n_32),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_30),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_30),
.A2(n_31),
.B1(n_158),
.B2(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_30),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_30),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_35),
.A2(n_123),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_36),
.B(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_40),
.A2(n_49),
.B1(n_92),
.B2(n_125),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_42),
.B(n_248),
.Y(n_247)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_50),
.B1(n_52),
.B2(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_45),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_45),
.A2(n_52),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_49),
.A2(n_125),
.B(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_49),
.A2(n_176),
.B(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_49),
.B(n_180),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_52),
.B(n_177),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_53),
.B(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_54),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_54),
.A2(n_152),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_55),
.A2(n_62),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_55),
.A2(n_128),
.B(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_75),
.A3(n_77),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_60),
.B(n_74),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_60),
.B(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B(n_80),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_72),
.B1(n_79),
.B2(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_72),
.A2(n_81),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_78),
.A2(n_111),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_85),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_97),
.B2(n_98),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_96),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_91),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_92),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_92),
.A2(n_229),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_118)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_102),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_118),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_131),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_121),
.B(n_124),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_151),
.B1(n_153),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_165),
.B(n_289),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_163),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_139),
.B(n_163),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_146),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_144),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_146),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_154),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_149),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_156),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_196),
.B(n_283),
.C(n_288),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_190),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_190),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_182),
.C(n_183),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_168),
.A2(n_169),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_174),
.C(n_178),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_182),
.B(n_183),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_277),
.B(n_282),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_230),
.B(n_276),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_219),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_201),
.B(n_219),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_212),
.C(n_216),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_202),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_205),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B(n_210),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_209),
.A2(n_253),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_212),
.A2(n_216),
.B1(n_217),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_226),
.C(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_270),
.B(n_275),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_249),
.B(n_269),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_243),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_247),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_258),
.B(n_268),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_256),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_263),
.B(n_267),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);


endmodule