module fake_netlist_1_10573_n_665 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_665);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_665;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_50), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_17), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_12), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_1), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_24), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_85), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
BUFx10_ASAP7_75t_L g99 ( .A(n_21), .Y(n_99) );
BUFx2_ASAP7_75t_SL g100 ( .A(n_51), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_40), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_38), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_58), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_37), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_86), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_66), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_10), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_63), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_28), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_36), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_6), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_0), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_43), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_9), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_56), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_23), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_9), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_21), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_64), .Y(n_127) );
INVxp33_ASAP7_75t_SL g128 ( .A(n_71), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_62), .Y(n_129) );
INVxp67_ASAP7_75t_SL g130 ( .A(n_34), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_102), .B(n_0), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_102), .B(n_2), .Y(n_133) );
CKINVDCx11_ASAP7_75t_R g134 ( .A(n_119), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
XNOR2xp5_ASAP7_75t_L g137 ( .A(n_121), .B(n_2), .Y(n_137) );
CKINVDCx8_ASAP7_75t_R g138 ( .A(n_89), .Y(n_138) );
INVx6_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_94), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_94), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_95), .B(n_3), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_125), .B(n_3), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_108), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_97), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_97), .A2(n_4), .B(n_5), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_113), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_101), .B(n_45), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_103), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_103), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_104), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_125), .B(n_8), .Y(n_157) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_104), .A2(n_8), .B(n_10), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_139), .B(n_98), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_135), .B(n_106), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_135), .B(n_106), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_131), .B(n_126), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_139), .B(n_113), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_154), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_139), .B(n_140), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_131), .B(n_123), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_131), .A2(n_126), .B1(n_110), .B2(n_90), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_139), .B(n_128), .Y(n_171) );
INVx6_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_140), .B(n_107), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_132), .B(n_124), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_131), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_132), .B(n_124), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_138), .B(n_111), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
AO22x2_ASAP7_75t_L g183 ( .A1(n_152), .A2(n_127), .B1(n_123), .B2(n_100), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_133), .B(n_144), .Y(n_184) );
INVxp33_ASAP7_75t_L g185 ( .A(n_134), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
INVxp67_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_138), .B(n_116), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
XNOR2x2_ASAP7_75t_L g191 ( .A(n_152), .B(n_137), .Y(n_191) );
AND2x6_ASAP7_75t_L g192 ( .A(n_133), .B(n_127), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_187), .B(n_144), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_184), .B(n_133), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_176), .B(n_156), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_162), .B(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_174), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_169), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_181), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_168), .B(n_147), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_162), .B(n_150), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_164), .B(n_145), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_181), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_186), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_191), .Y(n_208) );
OR2x2_ASAP7_75t_SL g209 ( .A(n_191), .B(n_137), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_162), .B(n_146), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_177), .Y(n_212) );
INVx6_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
INVx3_ASAP7_75t_SL g214 ( .A(n_169), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_184), .B(n_146), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_186), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_190), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_169), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_190), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_189), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_164), .B(n_156), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_189), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_182), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_184), .A2(n_153), .B(n_155), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_182), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_169), .A2(n_158), .B1(n_150), .B2(n_149), .Y(n_228) );
NOR2x1p5_ASAP7_75t_L g229 ( .A(n_185), .B(n_137), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_182), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_184), .B(n_157), .Y(n_231) );
BUFx12f_ASAP7_75t_L g232 ( .A(n_164), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_188), .B(n_157), .Y(n_233) );
AOI221xp5_ASAP7_75t_SL g234 ( .A1(n_170), .A2(n_153), .B1(n_155), .B2(n_122), .C(n_151), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_182), .Y(n_235) );
NAND2x1_ASAP7_75t_L g236 ( .A(n_169), .B(n_142), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_232), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_232), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_214), .A2(n_180), .B1(n_177), .B2(n_164), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_217), .Y(n_240) );
OAI22x1_ASAP7_75t_L g241 ( .A1(n_208), .A2(n_229), .B1(n_204), .B2(n_209), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_222), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_203), .B(n_179), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_219), .B(n_180), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_219), .B(n_180), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_195), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_214), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_193), .A2(n_175), .B(n_178), .C(n_163), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_203), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_219), .B(n_159), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_201), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_210), .A2(n_165), .B(n_171), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
NOR2x1_ASAP7_75t_SL g258 ( .A(n_201), .B(n_161), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_229), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_205), .B(n_141), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_205), .B(n_192), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_196), .A2(n_160), .B(n_149), .C(n_143), .Y(n_263) );
AND2x6_ASAP7_75t_L g264 ( .A(n_211), .B(n_192), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_205), .B(n_192), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_205), .A2(n_222), .B1(n_216), .B2(n_211), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_222), .B(n_192), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_211), .B(n_216), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_216), .B(n_161), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_222), .A2(n_192), .B1(n_183), .B2(n_161), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_215), .B(n_192), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_231), .A2(n_189), .B(n_173), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_233), .B(n_141), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_225), .A2(n_173), .B(n_155), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_207), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_194), .B(n_207), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_217), .Y(n_277) );
BUFx10_ASAP7_75t_L g278 ( .A(n_197), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_199), .Y(n_280) );
NOR2x1_ASAP7_75t_SL g281 ( .A(n_252), .B(n_199), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_272), .A2(n_225), .B(n_235), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_256), .A2(n_226), .B(n_204), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_252), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_250), .A2(n_198), .B(n_194), .C(n_109), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_240), .A2(n_204), .B(n_228), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_261), .A2(n_273), .B1(n_270), .B2(n_241), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_252), .B(n_212), .Y(n_288) );
O2A1O1Ixp5_ASAP7_75t_L g289 ( .A1(n_254), .A2(n_236), .B(n_220), .C(n_218), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_247), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_276), .A2(n_227), .B(n_235), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_243), .B(n_234), .C(n_136), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_241), .A2(n_253), .B1(n_242), .B2(n_260), .Y(n_294) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_279), .A2(n_148), .B(n_200), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_252), .B(n_212), .Y(n_296) );
CKINVDCx6p67_ASAP7_75t_R g297 ( .A(n_238), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_280), .A2(n_227), .B(n_230), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_248), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_251), .B(n_200), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_278), .Y(n_301) );
INVx6_ASAP7_75t_L g302 ( .A(n_278), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_275), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_278), .Y(n_304) );
XOR2xp5_ASAP7_75t_L g305 ( .A(n_237), .B(n_183), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_254), .A2(n_230), .B(n_218), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_246), .B(n_212), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_246), .B(n_202), .Y(n_308) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_274), .A2(n_148), .B(n_206), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_240), .A2(n_236), .B(n_202), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_266), .A2(n_183), .B1(n_192), .B2(n_220), .Y(n_311) );
INVx8_ASAP7_75t_L g312 ( .A(n_264), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_238), .A2(n_183), .B1(n_129), .B2(n_120), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_277), .A2(n_206), .B(n_142), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_277), .A2(n_148), .B(n_112), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_299), .B(n_209), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_287), .B(n_237), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_305), .A2(n_134), .B1(n_260), .B2(n_265), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_311), .A2(n_262), .B1(n_239), .B2(n_267), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_314), .A2(n_263), .B1(n_118), .B2(n_245), .C(n_151), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_304), .B(n_259), .Y(n_323) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_305), .A2(n_245), .B1(n_149), .B2(n_142), .C(n_143), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_299), .B(n_217), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_311), .A2(n_246), .B1(n_212), .B2(n_224), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_286), .A2(n_257), .B(n_148), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_282), .A2(n_269), .B(n_268), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_300), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_300), .B(n_217), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_301), .A2(n_264), .B1(n_249), .B2(n_224), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_293), .A2(n_269), .B(n_268), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_301), .A2(n_249), .B1(n_259), .B2(n_217), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_315), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_308), .A2(n_224), .B1(n_264), .B2(n_99), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_302), .A2(n_264), .B1(n_100), .B2(n_99), .Y(n_336) );
AOI211x1_ASAP7_75t_L g337 ( .A1(n_292), .A2(n_117), .B(n_115), .C(n_114), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_297), .A2(n_259), .B1(n_257), .B2(n_255), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
BUFx4f_ASAP7_75t_SL g341 ( .A(n_297), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_290), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_308), .A2(n_224), .B1(n_264), .B2(n_257), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_291), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
OAI33xp33_ASAP7_75t_L g348 ( .A1(n_317), .A2(n_291), .A3(n_303), .B1(n_285), .B2(n_313), .B3(n_293), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_320), .B(n_281), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_318), .B(n_294), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_334), .Y(n_351) );
AO21x2_ASAP7_75t_L g352 ( .A1(n_332), .A2(n_286), .B(n_316), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_317), .B(n_303), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_342), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_342), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_329), .B(n_295), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_343), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_334), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_329), .B(n_313), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_319), .B(n_307), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_343), .B(n_295), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_345), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_346), .B(n_295), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_345), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_346), .B(n_309), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_325), .B(n_309), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_322), .A2(n_312), .B1(n_302), .B2(n_304), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_338), .B(n_309), .Y(n_371) );
OAI222xp33_ASAP7_75t_L g372 ( .A1(n_326), .A2(n_306), .B1(n_307), .B2(n_284), .C1(n_149), .C2(n_151), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_323), .B(n_281), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_327), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_356), .B(n_337), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_351), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_351), .Y(n_379) );
AND3x1_ASAP7_75t_L g380 ( .A(n_350), .B(n_341), .C(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_366), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_358), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_366), .B(n_150), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_360), .A2(n_321), .B1(n_324), .B2(n_323), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_349), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_363), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_373), .A2(n_312), .B(n_323), .C(n_331), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_366), .B(n_150), .Y(n_390) );
AOI331xp33_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_335), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_15), .C1(n_11), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_368), .B(n_328), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_368), .B(n_150), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_368), .B(n_150), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_362), .B(n_158), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_362), .B(n_158), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_371), .B(n_367), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_362), .B(n_158), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_349), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_353), .B(n_307), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_364), .B(n_158), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_364), .B(n_158), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
OAI321xp33_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_339), .A3(n_333), .B1(n_292), .B2(n_344), .C(n_340), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_355), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_316), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_371), .B(n_316), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_356), .B(n_340), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_356), .B(n_283), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_404), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g412 ( .A1(n_385), .A2(n_353), .B(n_355), .C(n_357), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_404), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_381), .B(n_357), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_381), .B(n_369), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_406), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_401), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_376), .B(n_349), .C(n_373), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_410), .B(n_365), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_386), .B(n_387), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_410), .B(n_347), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_377), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_410), .B(n_347), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_377), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_409), .B(n_361), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_376), .B(n_369), .Y(n_430) );
NAND4xp25_ASAP7_75t_L g431 ( .A(n_385), .B(n_359), .C(n_143), .D(n_142), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_401), .B(n_361), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_393), .B(n_373), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_407), .B(n_347), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_378), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_409), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_393), .B(n_349), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_393), .B(n_349), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_407), .B(n_374), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_380), .B(n_370), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_407), .B(n_374), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_383), .B(n_367), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g444 ( .A(n_405), .B(n_348), .C(n_143), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_382), .B(n_367), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_378), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_392), .B(n_352), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_379), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_392), .B(n_352), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_387), .Y(n_450) );
NAND2xp33_ASAP7_75t_SL g451 ( .A(n_386), .B(n_340), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_382), .B(n_352), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_379), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_392), .B(n_352), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_392), .B(n_375), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_392), .B(n_375), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_386), .B(n_375), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_386), .B(n_359), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_397), .B(n_136), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_382), .B(n_136), .Y(n_460) );
INVx6_ASAP7_75t_L g461 ( .A(n_397), .Y(n_461) );
NAND2x2_ASAP7_75t_L g462 ( .A(n_428), .B(n_380), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_423), .B(n_398), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_431), .B(n_388), .C(n_394), .D(n_384), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_420), .B(n_397), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_420), .B(n_397), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_424), .B(n_397), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
AOI321xp33_ASAP7_75t_L g470 ( .A1(n_441), .A2(n_391), .A3(n_405), .B1(n_394), .B2(n_388), .C(n_384), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_412), .B(n_348), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_413), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_421), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_433), .B(n_408), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_430), .B(n_394), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_440), .B(n_395), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_400), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_426), .B(n_400), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_438), .B(n_408), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_439), .B(n_408), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_434), .B(n_400), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_428), .B(n_398), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
OAI31xp33_ASAP7_75t_L g485 ( .A1(n_431), .A2(n_372), .A3(n_402), .B(n_399), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_434), .B(n_389), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_440), .B(n_389), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_442), .B(n_389), .Y(n_489) );
NOR2xp67_ASAP7_75t_L g490 ( .A(n_419), .B(n_389), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_417), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_442), .B(n_395), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_421), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_422), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_444), .B(n_136), .C(n_384), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_422), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_450), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_426), .B(n_447), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_425), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_458), .B(n_379), .Y(n_500) );
OAI211xp5_ASAP7_75t_SL g501 ( .A1(n_432), .A2(n_142), .B(n_143), .C(n_149), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_457), .B(n_390), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_458), .B(n_390), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_416), .B(n_403), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_414), .B(n_403), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_460), .Y(n_506) );
XNOR2x2_ASAP7_75t_L g507 ( .A(n_419), .B(n_390), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_455), .B(n_395), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_437), .B(n_403), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_459), .B(n_396), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_443), .B(n_396), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_443), .B(n_396), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_423), .B(n_340), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_427), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_427), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_457), .B(n_399), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_447), .B(n_449), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_455), .B(n_399), .Y(n_519) );
AND2x4_ASAP7_75t_SL g520 ( .A(n_415), .B(n_456), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_402), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_497), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_463), .A2(n_423), .B1(n_415), .B2(n_418), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_521), .B(n_459), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_521), .B(n_454), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_498), .B(n_456), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_469), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_520), .B(n_415), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_503), .B(n_452), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_463), .A2(n_451), .B(n_391), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_462), .A2(n_461), .B1(n_415), .B2(n_452), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_512), .B(n_445), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_462), .A2(n_454), .B1(n_461), .B2(n_402), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_520), .Y(n_536) );
AOI32xp33_ASAP7_75t_L g537 ( .A1(n_501), .A2(n_436), .A3(n_429), .B1(n_448), .B2(n_336), .Y(n_537) );
NOR3xp33_ASAP7_75t_SL g538 ( .A(n_464), .B(n_372), .C(n_130), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_488), .B(n_429), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_518), .A2(n_436), .B(n_448), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_498), .B(n_461), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_473), .Y(n_543) );
AOI321xp33_ASAP7_75t_L g544 ( .A1(n_471), .A2(n_96), .A3(n_453), .B1(n_435), .B2(n_425), .C(n_446), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_478), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_475), .B(n_435), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_473), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_514), .A2(n_461), .B1(n_445), .B2(n_435), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_471), .A2(n_453), .B1(n_446), .B2(n_338), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_491), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_474), .B(n_11), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_513), .B(n_453), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g556 ( .A(n_470), .B(n_151), .C(n_289), .D(n_16), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_489), .B(n_136), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_494), .Y(n_558) );
BUFx2_ASAP7_75t_SL g559 ( .A(n_502), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_495), .B(n_284), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_480), .B(n_13), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_516), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_500), .Y(n_565) );
OAI221xp5_ASAP7_75t_SL g566 ( .A1(n_485), .A2(n_151), .B1(n_284), .B2(n_17), .C(n_18), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_501), .A2(n_310), .B(n_283), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_509), .B(n_15), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_502), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_519), .B(n_16), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_484), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_502), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_504), .B(n_18), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_517), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_536), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_556), .A2(n_517), .B1(n_490), .B2(n_518), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_523), .A2(n_514), .B1(n_517), .B2(n_476), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_556), .A2(n_479), .B1(n_477), .B2(n_505), .Y(n_578) );
XNOR2xp5_ASAP7_75t_L g579 ( .A(n_559), .B(n_482), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_553), .A2(n_508), .B1(n_506), .B2(n_510), .C1(n_511), .C2(n_492), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_531), .B(n_481), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_562), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_532), .A2(n_507), .B1(n_477), .B2(n_479), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_574), .A2(n_507), .B1(n_467), .B2(n_466), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_535), .A2(n_467), .B1(n_466), .B2(n_468), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g587 ( .A1(n_566), .A2(n_468), .B(n_486), .C(n_484), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_543), .Y(n_588) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_537), .A2(n_499), .B(n_312), .C(n_298), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_534), .B(n_499), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_569), .B(n_19), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_564), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g593 ( .A1(n_544), .A2(n_538), .B(n_570), .C(n_568), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_572), .B(n_19), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_522), .B(n_20), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_524), .B(n_20), .Y(n_597) );
AO22x2_ASAP7_75t_L g598 ( .A1(n_533), .A2(n_307), .B1(n_296), .B2(n_288), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_565), .B(n_310), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_530), .A2(n_312), .B1(n_296), .B2(n_288), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_555), .B(n_526), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_541), .A2(n_296), .B(n_288), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
OAI211xp5_ASAP7_75t_SL g604 ( .A1(n_563), .A2(n_298), .B(n_223), .C(n_221), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_542), .B(n_22), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g606 ( .A1(n_554), .A2(n_296), .B(n_288), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_543), .B(n_26), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_573), .A2(n_27), .B(n_29), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_557), .A2(n_30), .B(n_31), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_587), .A2(n_561), .B(n_548), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_593), .A2(n_548), .B(n_550), .C(n_560), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_577), .A2(n_550), .B(n_547), .Y(n_614) );
OAI211xp5_ASAP7_75t_L g615 ( .A1(n_584), .A2(n_551), .B(n_525), .C(n_567), .Y(n_615) );
NOR2x1_ASAP7_75t_SL g616 ( .A(n_589), .B(n_527), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_576), .A2(n_546), .B1(n_540), .B2(n_558), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_583), .B(n_552), .Y(n_618) );
AOI322xp5_ASAP7_75t_L g619 ( .A1(n_585), .A2(n_539), .A3(n_545), .B1(n_571), .B2(n_567), .C1(n_312), .C2(n_167), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_582), .Y(n_620) );
AOI31xp33_ASAP7_75t_L g621 ( .A1(n_587), .A2(n_578), .A3(n_579), .B(n_581), .Y(n_621) );
OAI31xp33_ASAP7_75t_L g622 ( .A1(n_598), .A2(n_258), .A3(n_264), .B(n_35), .Y(n_622) );
AND3x4_ASAP7_75t_L g623 ( .A(n_581), .B(n_32), .C(n_33), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_255), .B1(n_172), .B2(n_213), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_598), .A2(n_39), .B(n_41), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_588), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_594), .B(n_167), .C(n_217), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_592), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_597), .A2(n_167), .B1(n_255), .B2(n_221), .C(n_223), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_580), .A2(n_42), .B1(n_44), .B2(n_46), .C(n_47), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_580), .A2(n_172), .B1(n_213), .B2(n_167), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g632 ( .A1(n_604), .A2(n_255), .B(n_49), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_621), .B(n_609), .C(n_595), .Y(n_633) );
AOI221x1_ASAP7_75t_L g634 ( .A1(n_611), .A2(n_591), .B1(n_596), .B2(n_607), .C(n_603), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_613), .A2(n_588), .B(n_608), .C(n_602), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_626), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_611), .A2(n_610), .B(n_605), .C(n_606), .Y(n_637) );
AOI211x1_ASAP7_75t_L g638 ( .A1(n_614), .A2(n_600), .B(n_599), .C(n_601), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_612), .B(n_590), .Y(n_639) );
AO221x1_ASAP7_75t_L g640 ( .A1(n_625), .A2(n_48), .B1(n_54), .B2(n_55), .C(n_61), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g641 ( .A(n_623), .B(n_65), .C(n_67), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_616), .A2(n_167), .B1(n_172), .B2(n_213), .C1(n_73), .C2(n_75), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_618), .Y(n_643) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_622), .B(n_68), .C(n_69), .D(n_70), .E(n_76), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_618), .Y(n_645) );
AND4x1_ASAP7_75t_L g646 ( .A(n_633), .B(n_617), .C(n_629), .D(n_624), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_638), .A2(n_620), .B1(n_615), .B2(n_628), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_636), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_641), .B(n_627), .Y(n_649) );
NOR4xp75_ASAP7_75t_SL g650 ( .A(n_634), .B(n_619), .C(n_632), .D(n_630), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_643), .B(n_631), .Y(n_651) );
AOI211x1_ASAP7_75t_SL g652 ( .A1(n_641), .A2(n_77), .B(n_78), .C(n_79), .Y(n_652) );
OAI222xp33_ASAP7_75t_L g653 ( .A1(n_647), .A2(n_635), .B1(n_637), .B2(n_645), .C1(n_639), .C2(n_642), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_648), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_648), .B(n_644), .C(n_640), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_652), .B(n_80), .C(n_81), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_654), .Y(n_657) );
INVx3_ASAP7_75t_L g658 ( .A(n_653), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_655), .A2(n_651), .B1(n_649), .B2(n_650), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_657), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_658), .Y(n_661) );
AOI222xp33_ASAP7_75t_SL g662 ( .A1(n_661), .A2(n_659), .B1(n_646), .B2(n_656), .C1(n_651), .C2(n_88), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_661), .B1(n_660), .B2(n_213), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_167), .B(n_83), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_82), .B1(n_84), .B2(n_87), .C1(n_221), .C2(n_223), .Y(n_665) );
endmodule