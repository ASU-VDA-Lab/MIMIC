module fake_jpeg_21688_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_51),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_31),
.B1(n_36),
.B2(n_17),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_41),
.B1(n_49),
.B2(n_42),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_18),
.B1(n_19),
.B2(n_34),
.Y(n_80)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_79),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_41),
.B1(n_23),
.B2(n_33),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_35),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_80),
.A2(n_93),
.B1(n_27),
.B2(n_32),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_103),
.Y(n_130)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_84),
.Y(n_131)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_86),
.B(n_107),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_49),
.B1(n_50),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_102),
.B1(n_32),
.B2(n_27),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_41),
.B1(n_44),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_42),
.B1(n_44),
.B2(n_19),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_106),
.Y(n_132)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_37),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_21),
.Y(n_121)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_18),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_115),
.A2(n_118),
.B1(n_127),
.B2(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_116),
.B(n_16),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_125),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_36),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_101),
.B1(n_111),
.B2(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_47),
.B1(n_45),
.B2(n_30),
.Y(n_135)
);

NOR2x1p5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_47),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_149),
.B(n_113),
.C(n_92),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_83),
.B1(n_84),
.B2(n_94),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_25),
.A3(n_24),
.B1(n_16),
.B2(n_95),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_151),
.A2(n_179),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_83),
.B1(n_90),
.B2(n_108),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_154),
.B1(n_142),
.B2(n_28),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_136),
.B1(n_120),
.B2(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_159),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_85),
.B1(n_88),
.B2(n_109),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_168),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_21),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_81),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_81),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_176),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_140),
.B1(n_105),
.B2(n_131),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_170),
.A2(n_172),
.B1(n_167),
.B2(n_131),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_117),
.A2(n_124),
.B(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_183),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_76),
.B1(n_88),
.B2(n_109),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_76),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_180),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_16),
.B1(n_28),
.B2(n_26),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_126),
.B(n_16),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_126),
.B(n_125),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_135),
.B1(n_146),
.B2(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_189),
.B1(n_198),
.B2(n_202),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_162),
.A2(n_146),
.B1(n_137),
.B2(n_119),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_137),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_119),
.C(n_133),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_205),
.C(n_207),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_142),
.B1(n_28),
.B2(n_26),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_21),
.B(n_26),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_212),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_181),
.C(n_168),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_17),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_17),
.C(n_8),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_214),
.B1(n_9),
.B2(n_15),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_211),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_8),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_158),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_163),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_224),
.B(n_231),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_151),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_165),
.C(n_156),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_242),
.C(n_207),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_169),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_175),
.B(n_154),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_154),
.B(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_238),
.B1(n_212),
.B2(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_190),
.B(n_9),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_241),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_160),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_10),
.C(n_14),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_262),
.B1(n_228),
.B2(n_227),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_189),
.B1(n_187),
.B2(n_211),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_251),
.B1(n_261),
.B2(n_236),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_203),
.B(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_258),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_202),
.B1(n_203),
.B2(n_194),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_237),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_222),
.Y(n_258)
);

OAI22x1_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_193),
.B1(n_215),
.B2(n_199),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_216),
.A2(n_191),
.B1(n_210),
.B2(n_197),
.Y(n_262)
);

XOR2x1_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_225),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_274),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_276),
.B1(n_278),
.B2(n_280),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_244),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_225),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_220),
.C(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_228),
.B1(n_220),
.B2(n_248),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_241),
.C(n_226),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_277),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_244),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_245),
.A2(n_227),
.B1(n_235),
.B2(n_238),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_235),
.B1(n_210),
.B2(n_185),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_242),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_239),
.C(n_10),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_260),
.B1(n_255),
.B2(n_249),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_292),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_256),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_274),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_259),
.B1(n_247),
.B2(n_256),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_247),
.B1(n_257),
.B2(n_250),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_293),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_264),
.A2(n_257),
.B1(n_263),
.B2(n_6),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_282),
.B1(n_280),
.B2(n_273),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_305),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_303),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_286),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.C(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_306),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_285),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_267),
.B(n_286),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_13),
.B(n_15),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_287),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_277),
.B1(n_12),
.B2(n_8),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_318),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_296),
.B1(n_271),
.B2(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_4),
.C(n_5),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_307),
.B(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_320),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_322),
.B(n_319),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_325),
.C(n_315),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_318),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_15),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_7),
.C(n_4),
.Y(n_331)
);


endmodule