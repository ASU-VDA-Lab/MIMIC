module real_aes_3122_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_666;
wire n_320;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_904;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_996;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_363;
wire n_449;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_997;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_968;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
HB1xp67_ASAP7_75t_L g278 ( .A(n_0), .Y(n_278) );
AND2x4_ASAP7_75t_L g747 ( .A(n_0), .B(n_748), .Y(n_747) );
AND2x4_ASAP7_75t_L g753 ( .A(n_0), .B(n_265), .Y(n_753) );
AO22x1_ASAP7_75t_L g751 ( .A1(n_1), .A2(n_3), .B1(n_752), .B2(n_754), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_2), .A2(n_103), .B1(n_412), .B2(n_413), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_4), .A2(n_175), .B1(n_397), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_5), .A2(n_201), .B1(n_744), .B2(n_759), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_6), .A2(n_141), .B1(n_363), .B2(n_433), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_7), .A2(n_168), .B1(n_409), .B2(n_410), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_8), .A2(n_56), .B1(n_433), .B2(n_434), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_9), .B(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_10), .A2(n_90), .B1(n_327), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_11), .A2(n_111), .B1(n_982), .B2(n_983), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_12), .A2(n_208), .B1(n_375), .B2(n_378), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_13), .A2(n_252), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_14), .A2(n_220), .B1(n_439), .B2(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_15), .A2(n_615), .B(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_16), .A2(n_236), .B1(n_397), .B2(n_398), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_17), .A2(n_28), .B1(n_361), .B2(n_434), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_18), .A2(n_125), .B1(n_761), .B2(n_762), .Y(n_760) );
AO22x1_ASAP7_75t_L g417 ( .A1(n_19), .A2(n_151), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_20), .A2(n_52), .B1(n_447), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_21), .A2(n_160), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_22), .A2(n_240), .B1(n_381), .B2(n_383), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_23), .A2(n_195), .B1(n_363), .B2(n_482), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_24), .A2(n_211), .B1(n_349), .B2(n_566), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_25), .A2(n_153), .B1(n_489), .B2(n_603), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_26), .A2(n_245), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g313 ( .A(n_27), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_29), .A2(n_101), .B1(n_395), .B2(n_403), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_30), .A2(n_107), .B1(n_682), .B2(n_986), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_31), .A2(n_127), .B1(n_525), .B2(n_688), .Y(n_993) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_32), .A2(n_403), .B(n_404), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_33), .B(n_210), .Y(n_276) );
INVx1_ASAP7_75t_L g309 ( .A(n_33), .Y(n_309) );
INVxp67_ASAP7_75t_L g324 ( .A(n_33), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_34), .A2(n_123), .B1(n_361), .B2(n_363), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_35), .A2(n_216), .B1(n_315), .B2(n_442), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_36), .A2(n_70), .B1(n_354), .B2(n_525), .Y(n_524) );
AOI21xp33_ASAP7_75t_SL g589 ( .A1(n_37), .A2(n_537), .B(n_590), .Y(n_589) );
AO22x1_ASAP7_75t_L g411 ( .A1(n_38), .A2(n_143), .B1(n_412), .B2(n_413), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_39), .A2(n_69), .B1(n_395), .B2(n_403), .C(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_40), .A2(n_87), .B1(n_660), .B2(n_662), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_41), .B(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_42), .A2(n_110), .B1(n_409), .B2(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_43), .B(n_294), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_44), .A2(n_164), .B1(n_680), .B2(n_682), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_45), .A2(n_264), .B1(n_596), .B2(n_597), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_46), .A2(n_225), .B1(n_401), .B2(n_451), .Y(n_638) );
INVx1_ASAP7_75t_SL g543 ( .A(n_47), .Y(n_543) );
OAI21x1_ASAP7_75t_L g455 ( .A1(n_48), .A2(n_456), .B(n_473), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g473 ( .A(n_48), .B(n_457), .C(n_462), .D(n_469), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_49), .A2(n_75), .B1(n_288), .B2(n_375), .C(n_720), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_50), .A2(n_184), .B1(n_437), .B2(n_439), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_51), .A2(n_190), .B1(n_439), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_53), .A2(n_88), .B1(n_400), .B2(n_401), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_54), .A2(n_248), .B1(n_381), .B2(n_725), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_55), .A2(n_174), .B1(n_754), .B2(n_770), .Y(n_785) );
INVx1_ASAP7_75t_L g547 ( .A(n_57), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_58), .A2(n_163), .B1(n_368), .B2(n_371), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_59), .A2(n_112), .B1(n_381), .B2(n_383), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_60), .A2(n_241), .B1(n_418), .B2(n_419), .Y(n_650) );
INVx2_ASAP7_75t_L g273 ( .A(n_61), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_62), .B(n_395), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_63), .A2(n_451), .B(n_452), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_64), .A2(n_218), .B1(n_596), .B2(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g746 ( .A(n_65), .Y(n_746) );
AND2x4_ASAP7_75t_L g750 ( .A(n_65), .B(n_273), .Y(n_750) );
INVx1_ASAP7_75t_SL g758 ( .A(n_65), .Y(n_758) );
INVx1_ASAP7_75t_L g969 ( .A(n_66), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_67), .A2(n_203), .B1(n_410), .B2(n_416), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_68), .A2(n_215), .B1(n_418), .B2(n_419), .Y(n_708) );
XNOR2x1_ASAP7_75t_L g611 ( .A(n_71), .B(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_71), .A2(n_193), .B1(n_752), .B2(n_771), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_72), .A2(n_74), .B1(n_346), .B2(n_489), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_73), .A2(n_286), .B(n_312), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_76), .A2(n_156), .B1(n_433), .B2(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_77), .Y(n_294) );
XOR2x2_ASAP7_75t_L g509 ( .A(n_78), .B(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_79), .A2(n_154), .B1(n_397), .B2(n_398), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_80), .A2(n_191), .B1(n_400), .B2(n_401), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_81), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_82), .A2(n_185), .B1(n_397), .B2(n_398), .Y(n_467) );
INVx1_ASAP7_75t_L g540 ( .A(n_83), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_84), .A2(n_256), .B1(n_409), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_85), .A2(n_227), .B1(n_471), .B2(n_482), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_86), .A2(n_239), .B1(n_430), .B2(n_487), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_89), .A2(n_162), .B1(n_744), .B2(n_749), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_91), .A2(n_99), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_92), .A2(n_200), .B1(n_754), .B2(n_770), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_93), .A2(n_180), .B1(n_752), .B2(n_754), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_94), .A2(n_178), .B1(n_413), .B2(n_415), .Y(n_649) );
INVx1_ASAP7_75t_L g295 ( .A(n_95), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_95), .B(n_209), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_96), .A2(n_166), .B1(n_562), .B2(n_609), .Y(n_624) );
INVx1_ASAP7_75t_L g465 ( .A(n_97), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_98), .A2(n_104), .B1(n_349), .B2(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g453 ( .A(n_100), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_102), .A2(n_122), .B1(n_664), .B2(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_105), .A2(n_171), .B1(n_744), .B2(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g974 ( .A(n_106), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_108), .A2(n_116), .B1(n_744), .B2(n_759), .Y(n_780) );
INVx1_ASAP7_75t_L g405 ( .A(n_109), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_113), .A2(n_187), .B1(n_346), .B2(n_489), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_114), .A2(n_261), .B1(n_409), .B2(n_412), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_115), .A2(n_144), .B1(n_553), .B2(n_669), .C(n_671), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_115), .A2(n_144), .B1(n_553), .B2(n_669), .C(n_671), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_117), .A2(n_181), .B1(n_409), .B2(n_412), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_118), .A2(n_217), .B1(n_445), .B2(n_447), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_119), .A2(n_213), .B1(n_767), .B2(n_847), .Y(n_846) );
OA21x2_ASAP7_75t_L g635 ( .A1(n_120), .A2(n_636), .B(n_651), .Y(n_635) );
INVx1_ASAP7_75t_L g654 ( .A(n_120), .Y(n_654) );
INVx1_ASAP7_75t_L g499 ( .A(n_121), .Y(n_499) );
XNOR2x1_ASAP7_75t_L g478 ( .A(n_124), .B(n_479), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_126), .A2(n_255), .B1(n_744), .B2(n_759), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_128), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_129), .A2(n_263), .B1(n_349), .B2(n_354), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_130), .A2(n_189), .B1(n_340), .B2(n_346), .Y(n_339) );
AO22x1_ASAP7_75t_L g414 ( .A1(n_131), .A2(n_260), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_132), .A2(n_139), .B1(n_340), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_133), .A2(n_197), .B1(n_437), .B2(n_989), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_134), .A2(n_219), .B1(n_410), .B2(n_416), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_135), .A2(n_237), .B1(n_413), .B2(n_415), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_136), .A2(n_229), .B1(n_363), .B2(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g519 ( .A(n_137), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_138), .A2(n_233), .B1(n_730), .B2(n_731), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_140), .A2(n_238), .B1(n_349), .B2(n_354), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_142), .A2(n_188), .B1(n_687), .B2(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g515 ( .A(n_145), .Y(n_515) );
INVx1_ASAP7_75t_L g574 ( .A(n_146), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_147), .A2(n_221), .B1(n_412), .B2(n_413), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_148), .A2(n_152), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI21xp33_ASAP7_75t_SL g536 ( .A1(n_149), .A2(n_537), .B(n_539), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_150), .A2(n_161), .B1(n_561), .B2(n_562), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_155), .A2(n_253), .B1(n_757), .B2(n_759), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_157), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g643 ( .A(n_158), .Y(n_643) );
CKINVDCx14_ASAP7_75t_R g696 ( .A(n_159), .Y(n_696) );
INVx1_ASAP7_75t_L g979 ( .A(n_165), .Y(n_979) );
XNOR2x2_ASAP7_75t_L g391 ( .A(n_167), .B(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_169), .A2(n_224), .B1(n_762), .B2(n_770), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_170), .B(n_501), .Y(n_703) );
INVx1_ASAP7_75t_L g968 ( .A(n_172), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_173), .A2(n_965), .B1(n_998), .B2(n_999), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_173), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_176), .A2(n_243), .B1(n_349), .B2(n_484), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_177), .A2(n_222), .B1(n_494), .B2(n_496), .C(n_498), .Y(n_493) );
AO221x2_ASAP7_75t_L g743 ( .A1(n_179), .A2(n_231), .B1(n_744), .B2(n_749), .C(n_751), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_182), .B(n_327), .Y(n_619) );
OA22x2_ASAP7_75t_L g299 ( .A1(n_183), .A2(n_210), .B1(n_294), .B2(n_298), .Y(n_299) );
INVx1_ASAP7_75t_L g337 ( .A(n_183), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_186), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g528 ( .A(n_192), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_194), .A2(n_212), .B1(n_315), .B2(n_378), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_196), .A2(n_207), .B1(n_522), .B2(n_523), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_198), .A2(n_249), .B1(n_459), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_199), .A2(n_258), .B1(n_770), .B2(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g591 ( .A(n_202), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_204), .A2(n_232), .B1(n_371), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_205), .A2(n_251), .B1(n_378), .B2(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_206), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g311 ( .A(n_209), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_209), .B(n_334), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_210), .A2(n_228), .B(n_325), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_214), .Y(n_716) );
INVx1_ASAP7_75t_SL g550 ( .A(n_223), .Y(n_550) );
INVx1_ASAP7_75t_L g583 ( .A(n_224), .Y(n_583) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_226), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_228), .B(n_257), .Y(n_277) );
INVx1_ASAP7_75t_L g297 ( .A(n_228), .Y(n_297) );
CKINVDCx16_ASAP7_75t_R g617 ( .A(n_230), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_234), .A2(n_244), .B1(n_445), .B2(n_447), .Y(n_492) );
INVx1_ASAP7_75t_L g976 ( .A(n_235), .Y(n_976) );
INVx1_ASAP7_75t_SL g527 ( .A(n_242), .Y(n_527) );
INVx1_ASAP7_75t_L g426 ( .A(n_246), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_247), .A2(n_400), .B(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_250), .A2(n_259), .B1(n_349), .B2(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g672 ( .A(n_254), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_257), .B(n_304), .Y(n_303) );
AOI222xp33_ASAP7_75t_L g961 ( .A1(n_258), .A2(n_962), .B1(n_994), .B2(n_997), .C1(n_1000), .C2(n_1002), .Y(n_961) );
XNOR2x1_ASAP7_75t_L g964 ( .A(n_258), .B(n_965), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_262), .B(n_545), .Y(n_571) );
INVx1_ASAP7_75t_L g748 ( .A(n_265), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_266), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_279), .B(n_737), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx4_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .C(n_278), .Y(n_270) );
AND2x2_ASAP7_75t_L g994 ( .A(n_271), .B(n_995), .Y(n_994) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_271), .B(n_996), .Y(n_1001) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OA21x2_ASAP7_75t_L g1003 ( .A1(n_272), .A2(n_758), .B(n_1004), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g745 ( .A(n_273), .B(n_746), .Y(n_745) );
AND3x4_ASAP7_75t_L g757 ( .A(n_273), .B(n_747), .C(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_274), .B(n_996), .Y(n_995) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_275), .A2(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g996 ( .A(n_278), .Y(n_996) );
XNOR2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_577), .Y(n_279) );
XNOR2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_421), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_387), .B1(n_388), .B2(n_420), .Y(n_281) );
INVx2_ASAP7_75t_SL g420 ( .A(n_282), .Y(n_420) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
XNOR2x1_ASAP7_75t_L g283 ( .A(n_284), .B(n_386), .Y(n_283) );
NAND4xp75_ASAP7_75t_L g284 ( .A(n_285), .B(n_338), .C(n_359), .D(n_373), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g449 ( .A(n_289), .Y(n_449) );
INVx2_ASAP7_75t_L g645 ( .A(n_289), .Y(n_645) );
INVx2_ASAP7_75t_L g670 ( .A(n_289), .Y(n_670) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g535 ( .A(n_290), .Y(n_535) );
BUFx3_ASAP7_75t_L g573 ( .A(n_290), .Y(n_573) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_300), .Y(n_290) );
AND2x2_ASAP7_75t_L g350 ( .A(n_291), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g369 ( .A(n_291), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g379 ( .A(n_291), .B(n_345), .Y(n_379) );
AND2x2_ASAP7_75t_L g395 ( .A(n_291), .B(n_300), .Y(n_395) );
AND2x4_ASAP7_75t_L g397 ( .A(n_291), .B(n_345), .Y(n_397) );
AND2x4_ASAP7_75t_L g409 ( .A(n_291), .B(n_365), .Y(n_409) );
AND2x4_ASAP7_75t_L g412 ( .A(n_291), .B(n_351), .Y(n_412) );
AND2x2_ASAP7_75t_L g681 ( .A(n_291), .B(n_351), .Y(n_681) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_299), .Y(n_291) );
INVx1_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
NAND2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g298 ( .A(n_294), .Y(n_298) );
INVx3_ASAP7_75t_L g304 ( .A(n_294), .Y(n_304) );
NAND2xp33_ASAP7_75t_L g310 ( .A(n_294), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_294), .Y(n_320) );
INVx1_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_297), .A2(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g322 ( .A(n_299), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
AND2x2_ASAP7_75t_L g377 ( .A(n_299), .B(n_343), .Y(n_377) );
AND2x2_ASAP7_75t_L g347 ( .A(n_300), .B(n_342), .Y(n_347) );
AND2x4_ASAP7_75t_L g382 ( .A(n_300), .B(n_377), .Y(n_382) );
AND2x4_ASAP7_75t_L g385 ( .A(n_300), .B(n_357), .Y(n_385) );
AND2x4_ASAP7_75t_L g401 ( .A(n_300), .B(n_357), .Y(n_401) );
AND2x2_ASAP7_75t_L g403 ( .A(n_300), .B(n_377), .Y(n_403) );
AND2x4_ASAP7_75t_L g419 ( .A(n_300), .B(n_342), .Y(n_419) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_306), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g318 ( .A(n_302), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g345 ( .A(n_302), .B(n_306), .Y(n_345) );
AND2x4_ASAP7_75t_L g351 ( .A(n_302), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g366 ( .A(n_302), .B(n_353), .Y(n_366) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_304), .B(n_309), .Y(n_308) );
INVxp67_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_305), .B(n_333), .C(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g353 ( .A(n_307), .Y(n_353) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_326), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g553 ( .A(n_316), .Y(n_553) );
INVx2_ASAP7_75t_L g597 ( .A(n_316), .Y(n_597) );
INVx3_ASAP7_75t_L g982 ( .A(n_316), .Y(n_982) );
INVx5_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx4f_ASAP7_75t_L g443 ( .A(n_317), .Y(n_443) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
AND2x4_ASAP7_75t_L g398 ( .A(n_318), .B(n_322), .Y(n_398) );
AND2x2_ASAP7_75t_L g640 ( .A(n_318), .B(n_322), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
INVx2_ASAP7_75t_L g541 ( .A(n_327), .Y(n_541) );
INVx4_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_328), .B(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_328), .B(n_643), .Y(n_642) );
INVx4_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g454 ( .A(n_329), .Y(n_454) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_330), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_334), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g357 ( .A(n_335), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_348), .Y(n_338) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g438 ( .A(n_341), .Y(n_438) );
BUFx12f_ASAP7_75t_L g489 ( .A(n_341), .Y(n_489) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
AND2x4_ASAP7_75t_L g362 ( .A(n_342), .B(n_351), .Y(n_362) );
AND2x4_ASAP7_75t_L g364 ( .A(n_342), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g415 ( .A(n_342), .B(n_351), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_342), .B(n_370), .Y(n_416) );
AND2x4_ASAP7_75t_L g418 ( .A(n_342), .B(n_345), .Y(n_418) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x4_ASAP7_75t_L g376 ( .A(n_345), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g400 ( .A(n_345), .B(n_377), .Y(n_400) );
INVx1_ASAP7_75t_L g529 ( .A(n_346), .Y(n_529) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g439 ( .A(n_347), .Y(n_439) );
BUFx5_ASAP7_75t_L g603 ( .A(n_347), .Y(n_603) );
INVx1_ASAP7_75t_L g992 ( .A(n_347), .Y(n_992) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx8_ASAP7_75t_L g525 ( .A(n_350), .Y(n_525) );
AND2x4_ASAP7_75t_L g356 ( .A(n_351), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g413 ( .A(n_351), .B(n_357), .Y(n_413) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx4_ASAP7_75t_L g484 ( .A(n_355), .Y(n_484) );
INVx4_ASAP7_75t_L g566 ( .A(n_355), .Y(n_566) );
INVx2_ASAP7_75t_L g605 ( .A(n_355), .Y(n_605) );
INVx8_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g372 ( .A(n_357), .B(n_365), .Y(n_372) );
AND2x4_ASAP7_75t_L g410 ( .A(n_357), .B(n_365), .Y(n_410) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_367), .Y(n_359) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx12f_ASAP7_75t_L g433 ( .A(n_362), .Y(n_433) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_362), .Y(n_482) );
BUFx3_ASAP7_75t_L g677 ( .A(n_363), .Y(n_677) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_364), .Y(n_434) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_364), .Y(n_471) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g370 ( .A(n_366), .Y(n_370) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_369), .Y(n_487) );
BUFx12f_ASAP7_75t_L g561 ( .A(n_369), .Y(n_561) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_369), .Y(n_609) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_369), .Y(n_730) );
BUFx3_ASAP7_75t_L g678 ( .A(n_371), .Y(n_678) );
BUFx12f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx6_ASAP7_75t_L g431 ( .A(n_372), .Y(n_431) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_380), .Y(n_373) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g442 ( .A(n_376), .Y(n_442) );
INVx1_ASAP7_75t_L g538 ( .A(n_376), .Y(n_538) );
BUFx3_ASAP7_75t_L g570 ( .A(n_376), .Y(n_570) );
INVx3_ASAP7_75t_L g551 ( .A(n_378), .Y(n_551) );
BUFx3_ASAP7_75t_L g662 ( .A(n_378), .Y(n_662) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g446 ( .A(n_379), .Y(n_446) );
BUFx3_ASAP7_75t_L g596 ( .A(n_379), .Y(n_596) );
BUFx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_382), .Y(n_451) );
INVx2_ASAP7_75t_L g495 ( .A(n_382), .Y(n_495) );
INVx2_ASAP7_75t_L g546 ( .A(n_382), .Y(n_546) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_382), .Y(n_665) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g725 ( .A(n_384), .Y(n_725) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_385), .Y(n_447) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_385), .Y(n_600) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_406), .Y(n_392) );
AND4x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .C(n_399), .D(n_402), .Y(n_393) );
INVx2_ASAP7_75t_L g497 ( .A(n_395), .Y(n_497) );
INVx4_ASAP7_75t_L g618 ( .A(n_398), .Y(n_618) );
NOR4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .C(n_414), .D(n_417), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
XOR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_506), .Y(n_421) );
AO22x2_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_475), .B1(n_503), .B2(n_505), .Y(n_422) );
INVx1_ASAP7_75t_L g505 ( .A(n_423), .Y(n_505) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_455), .B2(n_474), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
XNOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_440), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_429), .B(n_432), .C(n_435), .D(n_436), .Y(n_428) );
INVx1_ASAP7_75t_L g518 ( .A(n_430), .Y(n_518) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g461 ( .A(n_431), .Y(n_461) );
INVx5_ASAP7_75t_L g562 ( .A(n_431), .Y(n_562) );
INVx2_ASAP7_75t_L g731 ( .A(n_431), .Y(n_731) );
BUFx12f_ASAP7_75t_L g522 ( .A(n_433), .Y(n_522) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_433), .Y(n_687) );
BUFx3_ASAP7_75t_L g523 ( .A(n_434), .Y(n_523) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g459 ( .A(n_438), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_438), .A2(n_527), .B1(n_528), .B2(n_529), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .C(n_448), .D(n_450), .Y(n_440) );
INVx2_ASAP7_75t_L g661 ( .A(n_442), .Y(n_661) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g972 ( .A(n_446), .Y(n_972) );
INVx3_ASAP7_75t_L g548 ( .A(n_447), .Y(n_548) );
BUFx3_ASAP7_75t_L g666 ( .A(n_447), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_454), .B(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g983 ( .A(n_454), .Y(n_983) );
INVx2_ASAP7_75t_L g474 ( .A(n_455), .Y(n_474) );
AND3x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_462), .C(n_469), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g504 ( .A(n_477), .Y(n_504) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND4xp75_ASAP7_75t_L g479 ( .A(n_480), .B(n_485), .C(n_490), .D(n_493), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
BUFx3_ASAP7_75t_L g514 ( .A(n_487), .Y(n_514) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g599 ( .A(n_495), .Y(n_599) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
NOR2xp33_ASAP7_75t_R g671 ( .A(n_500), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g593 ( .A(n_502), .Y(n_593) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_502), .Y(n_722) );
INVxp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_554), .B2(n_575), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_530), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .C(n_526), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_515), .B1(n_516), .B2(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g986 ( .A(n_518), .Y(n_986) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_521), .B(n_524), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .C(n_549), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_536), .Y(n_531) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_535), .Y(n_588) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g622 ( .A(n_538), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_547), .B2(n_548), .Y(n_542) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g576 ( .A(n_555), .Y(n_576) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
XOR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_574), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_559), .B(n_567), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .C(n_564), .D(n_565), .Y(n_559) );
BUFx3_ASAP7_75t_L g682 ( .A(n_561), .Y(n_682) );
BUFx2_ASAP7_75t_L g688 ( .A(n_566), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .C(n_571), .D(n_572), .Y(n_567) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
XNOR2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_631), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_610), .B1(n_628), .B2(n_630), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g629 ( .A(n_582), .Y(n_629) );
XNOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NOR4xp75_ASAP7_75t_L g584 ( .A(n_585), .B(n_594), .C(n_601), .D(n_606), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g980 ( .A(n_587), .Y(n_980) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g615 ( .A(n_588), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
INVx2_ASAP7_75t_L g975 ( .A(n_599), .Y(n_975) );
INVx4_ASAP7_75t_L g977 ( .A(n_600), .Y(n_977) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
BUFx3_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g630 ( .A(n_610), .Y(n_630) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_623), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_620), .C(n_621), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_619), .Y(n_616) );
NAND4xp25_ASAP7_75t_SL g623 ( .A(n_624), .B(n_625), .C(n_626), .D(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_693), .B2(n_736), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_655), .B1(n_691), .B2(n_692), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g691 ( .A(n_635), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_646), .Y(n_636) );
INVxp67_ASAP7_75t_L g652 ( .A(n_637), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .C(n_641), .D(n_644), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_646), .B(n_654), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .C(n_649), .D(n_650), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_SL g692 ( .A(n_655), .Y(n_692) );
AO22x2_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_673), .B1(n_674), .B2(n_689), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_667), .C(n_673), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND4xp75_ASAP7_75t_SL g689 ( .A(n_658), .B(n_675), .C(n_683), .D(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_663), .Y(n_658) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_661), .A2(n_968), .B1(n_969), .B2(n_970), .Y(n_967) );
BUFx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_683), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVx2_ASAP7_75t_SL g736 ( .A(n_693), .Y(n_736) );
AO22x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_712), .B1(n_733), .B2(n_735), .Y(n_693) );
INVx2_ASAP7_75t_L g735 ( .A(n_694), .Y(n_735) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI21x1_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_709), .Y(n_695) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_696), .B(n_710), .C(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_704), .Y(n_698) );
INVx1_ASAP7_75t_L g711 ( .A(n_699), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .C(n_702), .D(n_703), .Y(n_699) );
INVxp67_ASAP7_75t_L g710 ( .A(n_704), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .C(n_707), .D(n_708), .Y(n_704) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_715), .Y(n_734) );
XNOR2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
OR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_726), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .C(n_724), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NAND4xp25_ASAP7_75t_SL g726 ( .A(n_727), .B(n_728), .C(n_729), .D(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_959), .B(n_961), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_886), .C(n_924), .Y(n_738) );
OAI221xp5_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_844), .B1(n_845), .B2(n_850), .C(n_870), .Y(n_739) );
NOR4xp25_ASAP7_75t_L g740 ( .A(n_741), .B(n_815), .C(n_829), .D(n_837), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_763), .B(n_781), .C(n_808), .Y(n_741) );
INVx1_ASAP7_75t_L g813 ( .A(n_742), .Y(n_813) );
NOR2x1_ASAP7_75t_L g912 ( .A(n_742), .B(n_818), .Y(n_912) );
OR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_755), .Y(n_742) );
INVx1_ASAP7_75t_L g799 ( .A(n_743), .Y(n_799) );
AND2x2_ASAP7_75t_L g828 ( .A(n_743), .B(n_792), .Y(n_828) );
AND2x2_ASAP7_75t_L g834 ( .A(n_743), .B(n_755), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_743), .B(n_789), .Y(n_922) );
OAI321xp33_ASAP7_75t_L g943 ( .A1(n_743), .A2(n_826), .A3(n_918), .B1(n_944), .B2(n_945), .C(n_947), .Y(n_943) );
AND2x2_ASAP7_75t_L g957 ( .A(n_743), .B(n_788), .Y(n_957) );
INVx3_ASAP7_75t_L g848 ( .A(n_744), .Y(n_848) );
AND2x4_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
AND2x4_ASAP7_75t_L g752 ( .A(n_745), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g761 ( .A(n_745), .B(n_753), .Y(n_761) );
AND2x2_ASAP7_75t_L g770 ( .A(n_745), .B(n_753), .Y(n_770) );
AND2x4_ASAP7_75t_L g749 ( .A(n_747), .B(n_750), .Y(n_749) );
AND2x4_ASAP7_75t_L g759 ( .A(n_747), .B(n_750), .Y(n_759) );
AND2x2_ASAP7_75t_L g754 ( .A(n_750), .B(n_753), .Y(n_754) );
AND2x2_ASAP7_75t_L g762 ( .A(n_750), .B(n_753), .Y(n_762) );
AND2x4_ASAP7_75t_L g771 ( .A(n_750), .B(n_753), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_753), .Y(n_1004) );
INVx1_ASAP7_75t_L g792 ( .A(n_755), .Y(n_792) );
AND2x2_ASAP7_75t_L g804 ( .A(n_755), .B(n_789), .Y(n_804) );
AND2x2_ASAP7_75t_L g823 ( .A(n_755), .B(n_799), .Y(n_823) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .Y(n_755) );
INVx2_ASAP7_75t_SL g768 ( .A(n_759), .Y(n_768) );
INVx1_ASAP7_75t_L g940 ( .A(n_763), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_772), .Y(n_763) );
AND2x2_ASAP7_75t_L g800 ( .A(n_764), .B(n_777), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_764), .B(n_802), .Y(n_824) );
AND2x2_ASAP7_75t_L g836 ( .A(n_764), .B(n_826), .Y(n_836) );
OR2x2_ASAP7_75t_L g862 ( .A(n_764), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_764), .B(n_784), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_764), .B(n_844), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_764), .B(n_843), .Y(n_954) );
INVx4_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g853 ( .A(n_765), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g859 ( .A(n_765), .B(n_778), .Y(n_859) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_765), .B(n_823), .C(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g876 ( .A(n_765), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_765), .B(n_845), .Y(n_898) );
AND2x2_ASAP7_75t_L g901 ( .A(n_765), .B(n_826), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_765), .B(n_855), .Y(n_946) );
NOR3xp33_ASAP7_75t_SL g948 ( .A(n_765), .B(n_879), .C(n_915), .Y(n_948) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx2_ASAP7_75t_L g960 ( .A(n_771), .Y(n_960) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI332xp33_ASAP7_75t_L g913 ( .A1(n_773), .A2(n_858), .A3(n_914), .B1(n_917), .B2(n_918), .B3(n_919), .C1(n_920), .C2(n_923), .Y(n_913) );
OAI222xp33_ASAP7_75t_SL g930 ( .A1(n_773), .A2(n_788), .B1(n_843), .B2(n_931), .C1(n_935), .C2(n_936), .Y(n_930) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .Y(n_773) );
INVx4_ASAP7_75t_L g797 ( .A(n_774), .Y(n_797) );
OR2x2_ASAP7_75t_L g843 ( .A(n_774), .B(n_778), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_774), .B(n_807), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_774), .B(n_784), .Y(n_865) );
AND2x2_ASAP7_75t_L g868 ( .A(n_774), .B(n_777), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_774), .B(n_807), .Y(n_879) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g802 ( .A(n_777), .Y(n_802) );
OR2x2_ASAP7_75t_L g855 ( .A(n_777), .B(n_797), .Y(n_855) );
INVxp67_ASAP7_75t_L g863 ( .A(n_777), .Y(n_863) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_793), .B(n_800), .C(n_801), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
AND2x2_ASAP7_75t_L g831 ( .A(n_783), .B(n_827), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_783), .B(n_892), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_783), .B(n_822), .Y(n_905) );
AND2x2_ASAP7_75t_L g958 ( .A(n_783), .B(n_854), .Y(n_958) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g807 ( .A(n_784), .Y(n_807) );
AND2x2_ASAP7_75t_L g814 ( .A(n_784), .B(n_788), .Y(n_814) );
INVx3_ASAP7_75t_L g819 ( .A(n_784), .Y(n_819) );
AOI211xp5_ASAP7_75t_L g850 ( .A1(n_784), .A2(n_851), .B(n_856), .C(n_866), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_784), .B(n_922), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_784), .B(n_868), .Y(n_935) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g892 ( .A(n_787), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_792), .Y(n_787) );
AND2x2_ASAP7_75t_L g821 ( .A(n_788), .B(n_813), .Y(n_821) );
AND2x2_ASAP7_75t_L g833 ( .A(n_788), .B(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_788), .B(n_823), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_788), .B(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g880 ( .A(n_788), .B(n_828), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_788), .B(n_912), .Y(n_911) );
CKINVDCx6p67_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_789), .B(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g822 ( .A(n_789), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g827 ( .A(n_789), .B(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_L g842 ( .A(n_789), .B(n_813), .Y(n_842) );
AND2x2_ASAP7_75t_L g884 ( .A(n_789), .B(n_818), .Y(n_884) );
AND2x2_ASAP7_75t_L g928 ( .A(n_789), .B(n_874), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_789), .B(n_792), .Y(n_934) );
AND2x2_ASAP7_75t_L g941 ( .A(n_789), .B(n_792), .Y(n_941) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_792), .B(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_798), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_794), .B(n_883), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_794), .A2(n_926), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_925) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_795), .Y(n_929) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g806 ( .A(n_796), .Y(n_806) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g826 ( .A(n_797), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_799), .A2(n_817), .B1(n_888), .B2(n_890), .C(n_893), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_800), .A2(n_907), .B1(n_908), .B2(n_910), .C(n_913), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_800), .B(n_904), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx3_ASAP7_75t_SL g817 ( .A(n_802), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_802), .B(n_844), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_802), .B(n_845), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g919 ( .A(n_804), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g811 ( .A(n_806), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_807), .B(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_809), .B(n_911), .Y(n_910) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g904 ( .A(n_811), .Y(n_904) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x2_ASAP7_75t_L g883 ( .A(n_813), .B(n_884), .Y(n_883) );
INVxp67_ASAP7_75t_L g917 ( .A(n_814), .Y(n_917) );
OAI22xp33_ASAP7_75t_SL g815 ( .A1(n_816), .A2(n_820), .B1(n_824), .B2(n_825), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_817), .A2(n_940), .B1(n_941), .B2(n_942), .C(n_943), .Y(n_939) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_818), .B(n_840), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_818), .B(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g907 ( .A(n_818), .B(n_869), .Y(n_907) );
INVx3_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g874 ( .A(n_819), .B(n_834), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g955 ( .A(n_821), .Y(n_955) );
INVx1_ASAP7_75t_L g857 ( .A(n_822), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g956 ( .A1(n_822), .A2(n_957), .B(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g915 ( .A(n_823), .Y(n_915) );
INVx1_ASAP7_75t_L g871 ( .A(n_824), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
O2A1O1Ixp33_ASAP7_75t_L g881 ( .A1(n_826), .A2(n_832), .B(n_882), .C(n_885), .Y(n_881) );
INVx1_ASAP7_75t_L g936 ( .A(n_827), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_828), .B(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_828), .B(n_884), .Y(n_896) );
INVx1_ASAP7_75t_L g916 ( .A(n_828), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_832), .B(n_835), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_834), .B(n_884), .Y(n_927) );
INVx1_ASAP7_75t_L g944 ( .A(n_834), .Y(n_944) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
AOI21xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_841), .B(n_843), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g869 ( .A(n_840), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_841), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
OAI221xp5_ASAP7_75t_SL g886 ( .A1(n_845), .A2(n_887), .B1(n_897), .B2(n_899), .C(n_906), .Y(n_886) );
OAI221xp5_ASAP7_75t_SL g924 ( .A1(n_845), .A2(n_925), .B1(n_937), .B2(n_939), .C(n_949), .Y(n_924) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_853), .A2(n_890), .B1(n_950), .B2(n_951), .C(n_952), .Y(n_949) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_860), .B2(n_862), .C(n_864), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g889 ( .A(n_868), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_868), .B(n_895), .Y(n_894) );
AOI211xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B(n_875), .C(n_881), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_872), .A2(n_900), .B(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_885), .Y(n_951) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g950 ( .A(n_905), .Y(n_950) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g942 ( .A(n_911), .Y(n_942) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVxp67_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVxp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
OAI21xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .B(n_956), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_965), .Y(n_999) );
AND2x4_ASAP7_75t_L g965 ( .A(n_966), .B(n_984), .Y(n_965) );
NOR3xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_973), .C(n_978), .Y(n_966) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_974), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_973) );
OAI21xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_980), .B(n_981), .Y(n_978) );
AND4x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_987), .C(n_988), .D(n_993), .Y(n_984) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
endmodule