module fake_jpeg_13020_n_48 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_48);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_17),
.C(n_21),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.C(n_22),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_23),
.B1(n_5),
.B2(n_6),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_31),
.B(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.C(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_41),
.B1(n_7),
.B2(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_42),
.B1(n_36),
.B2(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.B(n_40),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_43),
.C(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_7),
.Y(n_48)
);


endmodule