module real_aes_9272_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_13;
wire n_41;
wire n_56;
wire n_34;
wire n_55;
wire n_12;
wire n_62;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_59;
wire n_53;
wire n_25;
wire n_47;
wire n_58;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_51;
wire n_54;
wire n_35;
wire n_42;
wire n_39;
wire n_60;
wire n_15;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_61;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_57;
wire n_44;
wire n_64;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_63;
wire n_33;
wire n_36;
INVx2_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
INVx1_ASAP7_75t_L g33 ( .A(n_0), .Y(n_33) );
INVx1_ASAP7_75t_L g39 ( .A(n_1), .Y(n_39) );
NAND2xp5_ASAP7_75t_L g41 ( .A(n_2), .B(n_42), .Y(n_41) );
HB1xp67_ASAP7_75t_L g58 ( .A(n_2), .Y(n_58) );
BUFx2_ASAP7_75t_L g54 ( .A(n_3), .Y(n_54) );
INVx1_ASAP7_75t_L g42 ( .A(n_4), .Y(n_42) );
INVx2_ASAP7_75t_L g26 ( .A(n_5), .Y(n_26) );
INVx1_ASAP7_75t_L g49 ( .A(n_6), .Y(n_49) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
INVx2_ASAP7_75t_L g23 ( .A(n_8), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_9), .B(n_38), .Y(n_37) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_11), .A2(n_34), .B1(n_43), .B2(n_60), .C(n_61), .Y(n_10) );
OAI21xp33_ASAP7_75t_L g11 ( .A1(n_12), .A2(n_24), .B(n_27), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_13), .B(n_17), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_13), .B(n_29), .Y(n_28) );
INVxp67_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_18), .B(n_21), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_23), .B(n_26), .Y(n_31) );
INVx2_ASAP7_75t_L g60 ( .A(n_24), .Y(n_60) );
INVx1_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
INVx1_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
OR2x6_ASAP7_75t_L g29 ( .A(n_30), .B(n_32), .Y(n_29) );
BUFx6f_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVx2_ASAP7_75t_SL g32 ( .A(n_33), .Y(n_32) );
BUFx2_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
AND2x4_ASAP7_75t_L g35 ( .A(n_36), .B(n_40), .Y(n_35) );
HB1xp67_ASAP7_75t_L g59 ( .A(n_36), .Y(n_59) );
INVx1_ASAP7_75t_L g36 ( .A(n_37), .Y(n_36) );
INVx1_ASAP7_75t_L g38 ( .A(n_39), .Y(n_38) );
INVx1_ASAP7_75t_L g40 ( .A(n_41), .Y(n_40) );
HB1xp67_ASAP7_75t_L g46 ( .A(n_42), .Y(n_46) );
INVx1_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
NOR2xp33_ASAP7_75t_L g44 ( .A(n_45), .B(n_47), .Y(n_44) );
INVx1_ASAP7_75t_SL g45 ( .A(n_46), .Y(n_45) );
NAND2xp5_ASAP7_75t_L g64 ( .A(n_46), .B(n_57), .Y(n_64) );
OAI22xp33_ASAP7_75t_SL g47 ( .A1(n_48), .A2(n_55), .B1(n_56), .B2(n_59), .Y(n_47) );
NAND2xp5_ASAP7_75t_L g62 ( .A(n_48), .B(n_63), .Y(n_62) );
NOR2xp33_ASAP7_75t_L g48 ( .A(n_49), .B(n_50), .Y(n_48) );
INVx5_ASAP7_75t_L g50 ( .A(n_51), .Y(n_50) );
BUFx8_ASAP7_75t_SL g51 ( .A(n_52), .Y(n_51) );
INVx2_ASAP7_75t_L g52 ( .A(n_53), .Y(n_52) );
BUFx2_ASAP7_75t_L g53 ( .A(n_54), .Y(n_53) );
CKINVDCx20_ASAP7_75t_R g55 ( .A(n_56), .Y(n_55) );
HB1xp67_ASAP7_75t_L g56 ( .A(n_57), .Y(n_56) );
INVx1_ASAP7_75t_L g57 ( .A(n_58), .Y(n_57) );
CKINVDCx16_ASAP7_75t_R g61 ( .A(n_62), .Y(n_61) );
INVx1_ASAP7_75t_L g63 ( .A(n_64), .Y(n_63) );
endmodule