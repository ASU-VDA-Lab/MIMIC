module fake_netlist_1_1065_n_653 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_653);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_653;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_10), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_64), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_56), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_51), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_46), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_37), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_10), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_54), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_43), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_27), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_30), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_2), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_25), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_34), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_59), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_31), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_22), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_66), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_44), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_73), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_71), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_28), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_75), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_45), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_53), .Y(n_102) );
NOR2xp67_ASAP7_75t_L g103 ( .A(n_1), .B(n_14), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_55), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_1), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_48), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_24), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_42), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_58), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_26), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_13), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_20), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_8), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_50), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_86), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_79), .B(n_0), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_79), .B(n_0), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_121), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_93), .B(n_3), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_119), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_78), .Y(n_140) );
BUFx3_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_77), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_78), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
BUFx8_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_113), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_81), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_111), .B(n_3), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_112), .B(n_4), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_112), .B(n_4), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_120), .B(n_5), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_101), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
OAI21x1_ASAP7_75t_L g160 ( .A1(n_104), .A2(n_38), .B(n_69), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_105), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_108), .B(n_5), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_76), .B(n_6), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_124), .A2(n_109), .B1(n_110), .B2(n_83), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_124), .B(n_115), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_150), .B(n_82), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_125), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_152), .A2(n_116), .B(n_114), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_134), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_135), .B(n_106), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_135), .B(n_85), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_135), .B(n_103), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_135), .B(n_122), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_125), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_125), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_137), .B(n_87), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_125), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_146), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_163), .B(n_97), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_126), .B(n_117), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_163), .B(n_123), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_163), .B(n_84), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_126), .B(n_102), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_141), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_125), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_133), .Y(n_205) );
AND2x6_ASAP7_75t_L g206 ( .A(n_157), .B(n_80), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_130), .B(n_123), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_144), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_161), .B(n_96), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_142), .B(n_98), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
INVx6_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_133), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_163), .B(n_99), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_133), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_137), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_161), .B(n_96), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_133), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_142), .B(n_92), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_133), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_220), .B(n_137), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_198), .A2(n_157), .B1(n_131), .B2(n_132), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_207), .B(n_130), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_210), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_165), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_165), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_220), .A2(n_128), .B1(n_157), .B2(n_152), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_169), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_210), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_171), .A2(n_128), .B1(n_118), .B2(n_106), .Y(n_236) );
BUFx4f_ASAP7_75t_SL g237 ( .A(n_179), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_179), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_167), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_207), .B(n_131), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
AND2x6_ASAP7_75t_L g243 ( .A(n_218), .B(n_154), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_171), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_221), .B(n_149), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_221), .B(n_132), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_213), .B(n_136), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_197), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_225), .B(n_136), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_182), .B(n_146), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_182), .B(n_146), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_185), .B(n_149), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_215), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_199), .B(n_146), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_199), .B(n_158), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_197), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_185), .A2(n_89), .B1(n_107), .B2(n_118), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_206), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_184), .B(n_155), .Y(n_262) );
AND3x2_ASAP7_75t_SL g263 ( .A(n_198), .B(n_87), .C(n_160), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_185), .B(n_158), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_206), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_167), .Y(n_266) );
OR2x6_ASAP7_75t_L g267 ( .A(n_185), .B(n_164), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_166), .B(n_164), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_202), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_218), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_172), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_198), .A2(n_156), .B1(n_153), .B2(n_161), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_204), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_223), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_208), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_215), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_184), .B(n_162), .Y(n_280) );
BUFx4f_ASAP7_75t_L g281 ( .A(n_206), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_218), .B(n_162), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_208), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_218), .B(n_155), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_206), .A2(n_148), .B1(n_139), .B2(n_156), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_184), .B(n_138), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_173), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_238), .B(n_169), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_231), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_270), .A2(n_206), .B1(n_183), .B2(n_166), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_237), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_267), .A2(n_206), .B1(n_223), .B2(n_209), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_231), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_281), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_256), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_244), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_245), .B(n_206), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_232), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_244), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_245), .B(n_184), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_230), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_235), .B(n_223), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_267), .A2(n_194), .B1(n_196), .B2(n_209), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_242), .Y(n_305) );
OAI21xp33_ASAP7_75t_L g306 ( .A1(n_228), .A2(n_170), .B(n_195), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_254), .Y(n_307) );
BUFx10_ASAP7_75t_L g308 ( .A(n_245), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_232), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_239), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_254), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_254), .Y(n_312) );
AND2x4_ASAP7_75t_SL g313 ( .A(n_267), .B(n_169), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_234), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_228), .A2(n_209), .B1(n_212), .B2(n_215), .Y(n_315) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_243), .B(n_191), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_267), .A2(n_209), .B1(n_178), .B2(n_169), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_256), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_243), .Y(n_319) );
AO32x2_ASAP7_75t_L g320 ( .A1(n_263), .A2(n_178), .A3(n_160), .B1(n_148), .B2(n_154), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_252), .B(n_212), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_259), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_252), .B(n_212), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_252), .B(n_212), .Y(n_324) );
BUFx2_ASAP7_75t_SL g325 ( .A(n_243), .Y(n_325) );
BUFx12f_ASAP7_75t_L g326 ( .A(n_227), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_239), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_255), .A2(n_191), .B(n_251), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_227), .B(n_178), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_246), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_268), .B(n_100), .C(n_90), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_281), .B(n_191), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_247), .B(n_178), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_330), .B(n_264), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_290), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_290), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_319), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_313), .A2(n_272), .B1(n_285), .B2(n_264), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_294), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_322), .A2(n_281), .B1(n_279), .B2(n_243), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_326), .A2(n_243), .B1(n_279), .B2(n_265), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_326), .A2(n_243), .B1(n_261), .B2(n_264), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_319), .B(n_234), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_300), .A2(n_285), .B1(n_280), .B2(n_262), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_SL g347 ( .A1(n_328), .A2(n_250), .B(n_229), .C(n_241), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_305), .B(n_257), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_313), .A2(n_233), .B1(n_282), .B2(n_284), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_302), .A2(n_280), .B1(n_262), .B2(n_236), .C(n_249), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_319), .A2(n_286), .B1(n_287), .B2(n_266), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_297), .A2(n_276), .B1(n_274), .B2(n_283), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_331), .A2(n_276), .B1(n_260), .B2(n_277), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_301), .B(n_276), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_292), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_288), .B1(n_258), .B2(n_275), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_297), .A2(n_263), .B1(n_85), .B2(n_92), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_308), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_298), .A2(n_248), .B1(n_269), .B2(n_273), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_211), .B1(n_217), .B2(n_222), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_323), .A2(n_287), .B1(n_266), .B2(n_273), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_339), .A2(n_329), .B1(n_291), .B2(n_325), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_348), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_338), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_357), .A2(n_329), .B1(n_308), .B2(n_333), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_356), .A2(n_308), .B1(n_333), .B2(n_303), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_309), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_345), .A2(n_293), .B1(n_304), .B2(n_317), .C(n_321), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_321), .B1(n_315), .B2(n_324), .C(n_316), .Y(n_371) );
CKINVDCx6p67_ASAP7_75t_R g372 ( .A(n_348), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_321), .B1(n_324), .B2(n_316), .C(n_139), .Y(n_373) );
INVx11_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_340), .B(n_309), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_347), .B(n_311), .C(n_312), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_310), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_349), .A2(n_303), .B1(n_321), .B2(n_323), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_346), .B(n_310), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_160), .B(n_332), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_335), .A2(n_327), .B1(n_314), .B2(n_332), .Y(n_382) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_355), .A2(n_303), .B1(n_289), .B2(n_323), .C1(n_217), .C2(n_222), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_336), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_363), .A2(n_327), .B1(n_289), .B2(n_334), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_360), .A2(n_148), .B1(n_138), .B2(n_154), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_352), .A2(n_295), .B1(n_334), .B2(n_318), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_354), .A2(n_192), .B1(n_193), .B2(n_173), .C(n_175), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_359), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_365), .B(n_343), .Y(n_391) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_366), .B(n_338), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_366), .A2(n_338), .B1(n_358), .B2(n_337), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_379), .A2(n_341), .B1(n_361), .B2(n_358), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_384), .Y(n_395) );
OAI31xp33_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_342), .A3(n_344), .B(n_337), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_365), .B(n_154), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_372), .Y(n_399) );
XNOR2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_6), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_377), .A2(n_362), .B(n_147), .Y(n_401) );
AOI33xp33_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_147), .A3(n_159), .B1(n_151), .B2(n_145), .B3(n_140), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_368), .A2(n_364), .B1(n_370), .B2(n_382), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
OAI22xp5_ASAP7_75t_SL g405 ( .A1(n_366), .A2(n_97), .B1(n_90), .B2(n_344), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_386), .Y(n_407) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_375), .Y(n_408) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_377), .A2(n_362), .B(n_151), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_373), .B(n_296), .Y(n_410) );
NOR2xp33_ASAP7_75t_R g411 ( .A(n_369), .B(n_344), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_383), .A2(n_334), .B1(n_318), .B2(n_296), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_369), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_384), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_383), .A2(n_318), .B1(n_296), .B2(n_295), .Y(n_415) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_387), .B(n_138), .C(n_141), .D(n_147), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_385), .A2(n_312), .B1(n_311), .B2(n_307), .Y(n_417) );
NAND4xp25_ASAP7_75t_SL g418 ( .A(n_374), .B(n_7), .C(n_9), .D(n_11), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_376), .B(n_138), .Y(n_419) );
OAI33xp33_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_145), .A3(n_140), .B1(n_147), .B2(n_151), .B3(n_159), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_376), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_378), .B(n_9), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_380), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_403), .A2(n_388), .B1(n_384), .B2(n_389), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_414), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_418), .A2(n_381), .B1(n_312), .B2(n_311), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_408), .A2(n_141), .B1(n_312), .B2(n_311), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_417), .A2(n_381), .B(n_145), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_414), .Y(n_431) );
NAND4xp75_ASAP7_75t_L g432 ( .A(n_392), .B(n_320), .C(n_145), .D(n_151), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_307), .B1(n_271), .B2(n_320), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_398), .B(n_127), .Y(n_434) );
OAI31xp33_ASAP7_75t_SL g435 ( .A1(n_394), .A2(n_320), .A3(n_14), .B(n_15), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_423), .B(n_12), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_402), .B(n_159), .C(n_140), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_391), .A2(n_159), .B1(n_127), .B2(n_140), .C(n_177), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_406), .B(n_320), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_411), .A2(n_127), .B(n_143), .Y(n_444) );
OAI33xp33_ASAP7_75t_L g445 ( .A1(n_407), .A2(n_127), .A3(n_16), .B1(n_17), .B2(n_18), .B3(n_19), .Y(n_445) );
OAI31xp33_ASAP7_75t_L g446 ( .A1(n_405), .A2(n_271), .A3(n_201), .B(n_200), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_307), .B1(n_143), .B2(n_133), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_15), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_413), .B(n_16), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_424), .B(n_17), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_421), .B(n_18), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_411), .A2(n_307), .B1(n_133), .B2(n_143), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_422), .B(n_399), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_19), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_390), .B(n_410), .C(n_397), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_401), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_398), .B(n_143), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_392), .B(n_143), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_401), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_419), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_416), .A2(n_176), .A3(n_226), .B1(n_224), .B2(n_219), .B3(n_216), .Y(n_461) );
OAI31xp33_ASAP7_75t_L g462 ( .A1(n_396), .A2(n_200), .A3(n_201), .B(n_177), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_409), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_409), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_409), .B(n_143), .Y(n_465) );
AO31x2_ASAP7_75t_L g466 ( .A1(n_420), .A2(n_402), .A3(n_180), .B(n_181), .Y(n_466) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_412), .A2(n_174), .B(n_226), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_393), .Y(n_469) );
OAI33xp33_ASAP7_75t_L g470 ( .A1(n_404), .A2(n_168), .A3(n_226), .B1(n_224), .B2(n_219), .B3(n_216), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_414), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_414), .Y(n_472) );
OAI221xp5_ASAP7_75t_SL g473 ( .A1(n_400), .A2(n_181), .B1(n_192), .B2(n_193), .C(n_219), .Y(n_473) );
OAI21x1_ASAP7_75t_L g474 ( .A1(n_417), .A2(n_188), .B(n_168), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_423), .B(n_143), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_442), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_436), .B(n_29), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_443), .B(n_471), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_453), .B(n_460), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_448), .B(n_32), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_443), .B(n_33), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_454), .B(n_35), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_426), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_448), .B(n_36), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_455), .B(n_168), .C(n_174), .D(n_176), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_471), .B(n_39), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_445), .B(n_174), .C(n_176), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_437), .Y(n_489) );
NOR2xp67_ASAP7_75t_SL g490 ( .A(n_458), .B(n_254), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_473), .B(n_214), .C(n_188), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_427), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_449), .B(n_40), .Y(n_493) );
INVx5_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_471), .B(n_41), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_444), .B(n_278), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_469), .B(n_47), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_444), .A2(n_240), .B(n_253), .C(n_57), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
OR2x6_ASAP7_75t_L g500 ( .A(n_472), .B(n_278), .Y(n_500) );
AOI31xp33_ASAP7_75t_L g501 ( .A1(n_452), .A2(n_49), .A3(n_52), .B(n_60), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_468), .A2(n_190), .B1(n_186), .B2(n_203), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_472), .B(n_61), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_427), .B(n_63), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_438), .B(n_188), .C(n_214), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_426), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_431), .B(n_65), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_431), .B(n_67), .Y(n_508) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_433), .B(n_68), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_449), .B(n_70), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_426), .B(n_186), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_437), .B(n_214), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_451), .B(n_216), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_475), .B(n_205), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_451), .B(n_205), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_463), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_468), .B(n_205), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_468), .B(n_224), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_435), .A2(n_187), .B1(n_186), .B2(n_190), .C(n_203), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_456), .B(n_187), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_435), .B(n_187), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_456), .B(n_186), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_463), .B(n_186), .Y(n_527) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_465), .A2(n_186), .B(n_190), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_428), .B(n_190), .C(n_203), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_429), .B(n_190), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_459), .B(n_441), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g532 ( .A(n_462), .B(n_240), .C(n_253), .D(n_190), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_441), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_501), .A2(n_505), .B(n_523), .C(n_497), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_489), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_519), .B(n_425), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_511), .B(n_425), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_497), .B(n_461), .C(n_470), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_479), .B(n_434), .Y(n_540) );
NAND2xp33_ASAP7_75t_SL g541 ( .A(n_483), .B(n_433), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_486), .B(n_432), .Y(n_542) );
AOI211xp5_ASAP7_75t_L g543 ( .A1(n_485), .A2(n_446), .B(n_462), .C(n_429), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_515), .B(n_459), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_506), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_514), .B(n_434), .Y(n_546) );
OAI22xp5_ASAP7_75t_SL g547 ( .A1(n_494), .A2(n_447), .B1(n_463), .B2(n_457), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_478), .B(n_499), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_478), .B(n_467), .Y(n_550) );
OAI21xp33_ASAP7_75t_L g551 ( .A1(n_525), .A2(n_434), .B(n_439), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_531), .B(n_467), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_494), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_494), .B(n_467), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_494), .B(n_446), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_483), .B(n_441), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_494), .B(n_464), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_481), .B(n_434), .Y(n_561) );
NAND2xp33_ASAP7_75t_L g562 ( .A(n_498), .B(n_432), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_533), .B(n_464), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_507), .B(n_464), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_477), .B(n_439), .C(n_440), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_508), .B(n_466), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_518), .B(n_466), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_503), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_482), .B(n_430), .Y(n_569) );
OR2x6_ASAP7_75t_L g570 ( .A(n_509), .B(n_465), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_503), .B(n_466), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_477), .B(n_457), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_487), .B(n_457), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_528), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_548), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_549), .B(n_552), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_554), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_537), .B(n_484), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_534), .Y(n_580) );
NAND2xp33_ASAP7_75t_SL g581 ( .A(n_547), .B(n_490), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_544), .B(n_520), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_537), .B(n_520), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_557), .A2(n_498), .B1(n_496), .B2(n_529), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_574), .Y(n_585) );
OAI22x1_ASAP7_75t_L g586 ( .A1(n_545), .A2(n_496), .B1(n_480), .B2(n_495), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_540), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_540), .B(n_527), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_559), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_563), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_553), .B(n_526), .Y(n_591) );
OAI22xp33_ASAP7_75t_SL g592 ( .A1(n_570), .A2(n_510), .B1(n_493), .B2(n_500), .Y(n_592) );
OAI32xp33_ASAP7_75t_L g593 ( .A1(n_541), .A2(n_532), .A3(n_530), .B1(n_516), .B2(n_502), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_538), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_567), .B(n_524), .Y(n_595) );
NAND3xp33_ASAP7_75t_SL g596 ( .A(n_535), .B(n_502), .C(n_488), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_561), .B(n_517), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_535), .B(n_527), .Y(n_599) );
INVx4_ASAP7_75t_L g600 ( .A(n_570), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_542), .B(n_512), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_572), .A2(n_457), .B(n_522), .Y(n_602) );
NAND4xp75_ASAP7_75t_L g603 ( .A(n_569), .B(n_517), .C(n_521), .D(n_430), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_562), .A2(n_512), .B(n_474), .C(n_491), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_539), .A2(n_500), .B1(n_512), .B2(n_430), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_570), .A2(n_500), .B1(n_474), .B2(n_513), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_556), .Y(n_608) );
XNOR2xp5_ASAP7_75t_L g609 ( .A(n_543), .B(n_500), .Y(n_609) );
INVx3_ASAP7_75t_SL g610 ( .A(n_573), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_558), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_560), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_551), .B(n_566), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_568), .B(n_564), .Y(n_614) );
AOI22x1_ASAP7_75t_L g615 ( .A1(n_555), .A2(n_539), .B1(n_565), .B2(n_571), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_565), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_557), .A2(n_494), .B1(n_554), .B2(n_535), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_537), .B(n_519), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_557), .A2(n_494), .B1(n_554), .B2(n_535), .Y(n_620) );
XOR2xp5_ASAP7_75t_L g621 ( .A(n_609), .B(n_597), .Y(n_621) );
NAND3xp33_ASAP7_75t_SL g622 ( .A(n_604), .B(n_599), .C(n_617), .Y(n_622) );
NOR4xp25_ASAP7_75t_L g623 ( .A(n_616), .B(n_596), .C(n_599), .D(n_620), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_576), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_579), .A2(n_613), .B1(n_594), .B2(n_583), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_592), .A2(n_593), .B(n_581), .C(n_584), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_581), .A2(n_600), .B(n_607), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_576), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_615), .A2(n_606), .B(n_585), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_600), .A2(n_587), .B1(n_606), .B2(n_619), .C1(n_601), .C2(n_589), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_600), .A2(n_586), .B(n_601), .Y(n_631) );
XNOR2xp5_ASAP7_75t_L g632 ( .A(n_598), .B(n_588), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_579), .A2(n_585), .B(n_610), .C(n_602), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_622), .A2(n_595), .B1(n_605), .B2(n_612), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_626), .A2(n_614), .B1(n_603), .B2(n_589), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_624), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_623), .A2(n_578), .B1(n_611), .B2(n_608), .C(n_618), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_633), .B(n_590), .Y(n_638) );
AO22x2_ASAP7_75t_L g639 ( .A1(n_627), .A2(n_578), .B1(n_575), .B2(n_580), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_631), .A2(n_577), .B1(n_582), .B2(n_591), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_636), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_635), .A2(n_623), .B1(n_625), .B2(n_629), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_639), .A2(n_621), .B1(n_632), .B2(n_628), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_640), .B(n_630), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_642), .B(n_637), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_641), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_643), .B(n_634), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_646), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_647), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_648), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_650), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_649), .B(n_645), .C(n_644), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_639), .B(n_638), .Y(n_653) );
endmodule