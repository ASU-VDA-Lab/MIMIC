module fake_jpeg_11344_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_54),
.Y(n_148)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_63),
.B(n_85),
.Y(n_112)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_106),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_10),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_103),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_48),
.Y(n_101)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_105),
.Y(n_130)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_72),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_51),
.B1(n_47),
.B2(n_48),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_122),
.A2(n_135),
.B1(n_141),
.B2(n_147),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_42),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_60),
.A2(n_47),
.B1(n_51),
.B2(n_50),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_54),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_136),
.B(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_43),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_142),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_62),
.A2(n_51),
.B1(n_47),
.B2(n_30),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_43),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_62),
.A2(n_84),
.B1(n_50),
.B2(n_96),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_75),
.A2(n_50),
.B1(n_49),
.B2(n_21),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_151),
.A2(n_155),
.B1(n_35),
.B2(n_31),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_72),
.A2(n_50),
.B1(n_49),
.B2(n_21),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_64),
.B(n_22),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_169),
.B(n_172),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_65),
.B(n_104),
.C(n_103),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_69),
.B(n_22),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_112),
.A2(n_21),
.B1(n_49),
.B2(n_34),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_175),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_20),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_178),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_45),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_182),
.Y(n_237)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_102),
.B1(n_98),
.B2(n_86),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_181),
.A2(n_191),
.B1(n_233),
.B2(n_162),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_134),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_44),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_189),
.A2(n_196),
.B(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_77),
.B1(n_82),
.B2(n_76),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_44),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_20),
.Y(n_197)
);

INVx5_ASAP7_75t_SL g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_198),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_147),
.A2(n_66),
.B1(n_61),
.B2(n_34),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_214),
.B1(n_216),
.B2(n_227),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_134),
.A2(n_34),
.B1(n_45),
.B2(n_41),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_202),
.B(n_206),
.Y(n_265)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_111),
.B(n_31),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_135),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_210),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_113),
.B(n_46),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_224),
.Y(n_258)
);

AO22x2_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_151),
.A2(n_45),
.B1(n_41),
.B2(n_44),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_218),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_141),
.A2(n_46),
.B1(n_37),
.B2(n_36),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_232),
.B1(n_120),
.B2(n_164),
.Y(n_261)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_220),
.B(n_222),
.Y(n_280)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_127),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_223),
.A2(n_0),
.B(n_1),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_114),
.B(n_46),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_234),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_117),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_127),
.A2(n_41),
.B1(n_35),
.B2(n_33),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_119),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_108),
.A2(n_37),
.B1(n_36),
.B2(n_20),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_120),
.B1(n_119),
.B2(n_131),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_37),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_231),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_159),
.B(n_36),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_143),
.A2(n_33),
.B1(n_10),
.B2(n_11),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_143),
.A2(n_10),
.B1(n_17),
.B2(n_16),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_137),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_0),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_152),
.B1(n_150),
.B2(n_153),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_239),
.A2(n_228),
.B1(n_203),
.B2(n_193),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_139),
.C(n_160),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_246),
.B(n_254),
.C(n_257),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_260),
.B1(n_264),
.B2(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_167),
.C(n_108),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_189),
.A2(n_204),
.B1(n_196),
.B2(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_256),
.A2(n_261),
.B1(n_273),
.B2(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_167),
.C(n_159),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_197),
.A2(n_162),
.B1(n_150),
.B2(n_131),
.Y(n_260)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

AO21x2_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_3),
.B(n_4),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_176),
.B(n_2),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_281),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_189),
.B1(n_196),
.B2(n_204),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_173),
.A2(n_229),
.B1(n_212),
.B2(n_179),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_277),
.A2(n_284),
.B1(n_287),
.B2(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_3),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_213),
.A2(n_220),
.B1(n_225),
.B2(n_226),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_177),
.B(n_11),
.C(n_16),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_185),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_213),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_213),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_293),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_213),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_300),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_198),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_298),
.B(n_306),
.Y(n_377)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

OA21x2_ASAP7_75t_R g300 ( 
.A1(n_258),
.A2(n_232),
.B(n_187),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_301),
.B(n_340),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_238),
.A2(n_209),
.B1(n_210),
.B2(n_223),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_333),
.B1(n_335),
.B2(n_295),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_241),
.A2(n_221),
.B(n_208),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_303),
.A2(n_339),
.B(n_311),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_190),
.C(n_194),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_276),
.C(n_288),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_305),
.A2(n_307),
.B1(n_312),
.B2(n_318),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_240),
.B(n_235),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_260),
.A2(n_234),
.B1(n_180),
.B2(n_217),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_251),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_313),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_314),
.B(n_320),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_240),
.B(n_192),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_326),
.Y(n_366)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_317),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_184),
.B1(n_183),
.B2(n_207),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_238),
.A2(n_195),
.B1(n_7),
.B2(n_8),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_319),
.A2(n_330),
.B1(n_255),
.B2(n_270),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_8),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_265),
.Y(n_323)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_6),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_334),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_237),
.B(n_12),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_262),
.B(n_12),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_329),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_287),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_332),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_275),
.A2(n_6),
.B1(n_13),
.B2(n_14),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_6),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_261),
.A2(n_6),
.B1(n_18),
.B2(n_242),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_336),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_254),
.B(n_18),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_338),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_271),
.B(n_18),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_241),
.A2(n_242),
.B(n_246),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_248),
.B(n_285),
.CI(n_273),
.CON(n_340),
.SN(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_341),
.A2(n_342),
.B1(n_259),
.B2(n_247),
.Y(n_373)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_343),
.A2(n_325),
.B1(n_310),
.B2(n_321),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_315),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_345),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_297),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

OA22x2_ASAP7_75t_L g347 ( 
.A1(n_300),
.A2(n_269),
.B1(n_289),
.B2(n_264),
.Y(n_347)
);

AOI22x1_ASAP7_75t_L g423 ( 
.A1(n_347),
.A2(n_381),
.B1(n_361),
.B2(n_355),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_348),
.A2(n_374),
.B1(n_387),
.B2(n_341),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_339),
.A2(n_243),
.B(n_269),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_353),
.A2(n_356),
.B(n_365),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_312),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_371),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_303),
.A2(n_269),
.B(n_283),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_302),
.A2(n_283),
.B1(n_250),
.B2(n_266),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_359),
.A2(n_360),
.B1(n_367),
.B2(n_307),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_335),
.A2(n_250),
.B1(n_266),
.B2(n_279),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_316),
.A2(n_236),
.B(n_290),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_276),
.B1(n_249),
.B2(n_279),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_249),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_376),
.C(n_381),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_318),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_336),
.A2(n_247),
.B1(n_259),
.B2(n_290),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_301),
.B(n_288),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_304),
.B(n_244),
.C(n_337),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_368),
.C(n_365),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_292),
.A2(n_244),
.B1(n_319),
.B2(n_333),
.Y(n_387)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_388),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_370),
.B(n_327),
.Y(n_389)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_345),
.A2(n_308),
.B1(n_292),
.B2(n_305),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_390),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_426)
);

NAND3xp33_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_294),
.C(n_296),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_391),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g392 ( 
.A(n_351),
.B(n_309),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_398),
.B(n_355),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_344),
.A2(n_305),
.B1(n_294),
.B2(n_330),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_348),
.A2(n_305),
.B1(n_296),
.B2(n_299),
.Y(n_396)
);

A2O1A1O1Ixp25_ASAP7_75t_L g398 ( 
.A1(n_351),
.A2(n_340),
.B(n_326),
.C(n_334),
.D(n_338),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_378),
.A2(n_305),
.B(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_388),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_353),
.A2(n_322),
.B(n_331),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_401),
.A2(n_349),
.B(n_362),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_357),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_406),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_356),
.A2(n_367),
.B1(n_375),
.B2(n_347),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_404),
.A2(n_409),
.B1(n_419),
.B2(n_379),
.Y(n_434)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_377),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_410),
.B1(n_420),
.B2(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_375),
.A2(n_340),
.B1(n_317),
.B2(n_342),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_343),
.A2(n_293),
.B1(n_324),
.B2(n_244),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_411),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_346),
.A2(n_244),
.B(n_384),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_416),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_380),
.C(n_363),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_349),
.Y(n_416)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_357),
.B(n_366),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_347),
.A2(n_354),
.B1(n_371),
.B2(n_360),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_364),
.A2(n_347),
.B1(n_376),
.B2(n_366),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_424),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_359),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_358),
.A2(n_379),
.B1(n_363),
.B2(n_372),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_425),
.A2(n_386),
.B1(n_369),
.B2(n_382),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_427),
.B(n_446),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_383),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_428),
.B(n_430),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_383),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_434),
.A2(n_392),
.B1(n_405),
.B2(n_408),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_435),
.B(n_439),
.C(n_443),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_423),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_448),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_380),
.C(n_372),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_400),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_362),
.C(n_385),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_369),
.B1(n_382),
.B2(n_385),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_447),
.B1(n_453),
.B2(n_458),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_425),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_421),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_412),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_455),
.C(n_456),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_402),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_422),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_420),
.A2(n_418),
.B1(n_407),
.B2(n_424),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_404),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_399),
.B(n_401),
.C(n_419),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_410),
.A2(n_390),
.B1(n_396),
.B2(n_403),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_459),
.Y(n_460)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_437),
.B(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_463),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_458),
.A2(n_393),
.B1(n_403),
.B2(n_400),
.Y(n_465)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_467),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_451),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_472),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_475),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_426),
.A2(n_392),
.B1(n_411),
.B2(n_414),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_476),
.Y(n_511)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_481),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_453),
.A2(n_398),
.B1(n_416),
.B2(n_449),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_426),
.A2(n_434),
.B1(n_441),
.B2(n_457),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_455),
.Y(n_492)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_430),
.C(n_428),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_436),
.C(n_448),
.Y(n_493)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g496 ( 
.A1(n_483),
.A2(n_485),
.B(n_486),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_450),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_484),
.B(n_487),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g485 ( 
.A(n_429),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_431),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_431),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_447),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_459),
.Y(n_509)
);

XNOR2x1_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_494),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_498),
.C(n_505),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_443),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_439),
.C(n_432),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_471),
.B(n_456),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_504),
.B(n_466),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_427),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_432),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_508),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_440),
.C(n_441),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_507),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_479),
.C(n_470),
.Y(n_508)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_479),
.B(n_445),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_469),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_503),
.A2(n_464),
.B1(n_478),
.B2(n_465),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_513),
.A2(n_525),
.B1(n_510),
.B2(n_511),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g541 ( 
.A(n_515),
.B(n_505),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_520),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_502),
.A2(n_480),
.B1(n_475),
.B2(n_460),
.Y(n_518)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_487),
.Y(n_519)
);

CKINVDCx14_ASAP7_75t_R g539 ( 
.A(n_519),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_502),
.A2(n_460),
.B1(n_488),
.B2(n_467),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_489),
.A2(n_472),
.B(n_464),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_523),
.A2(n_531),
.B(n_519),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_500),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_503),
.A2(n_483),
.B1(n_476),
.B2(n_474),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_491),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_526),
.B(n_527),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_489),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_530),
.Y(n_547)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_486),
.B(n_462),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_498),
.C(n_512),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_533),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_490),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_515),
.B(n_492),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_535),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_516),
.B(n_493),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_528),
.A2(n_500),
.B(n_501),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_537),
.A2(n_546),
.B(n_523),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_530),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_541),
.B(n_542),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_531),
.B(n_514),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_543),
.A2(n_544),
.B1(n_522),
.B2(n_525),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_513),
.A2(n_496),
.B1(n_506),
.B2(n_463),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_518),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_551),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_549),
.A2(n_550),
.B(n_540),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_546),
.A2(n_520),
.B(n_517),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_545),
.B(n_517),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_555),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_522),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_536),
.A2(n_504),
.B1(n_509),
.B2(n_529),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_557),
.B(n_558),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_529),
.C(n_494),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_537),
.Y(n_562)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_560),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_562),
.A2(n_549),
.B(n_547),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_552),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_SL g567 ( 
.A1(n_563),
.A2(n_539),
.B(n_547),
.C(n_554),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_550),
.B(n_544),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_566),
.B(n_538),
.C(n_540),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_567),
.B(n_570),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_569),
.A2(n_561),
.B(n_564),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_SL g572 ( 
.A1(n_568),
.A2(n_560),
.B(n_556),
.C(n_562),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_573),
.C(n_566),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_575),
.B(n_557),
.Y(n_576)
);

MAJx2_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_565),
.C(n_558),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_553),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_543),
.C(n_477),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_481),
.Y(n_579)
);


endmodule