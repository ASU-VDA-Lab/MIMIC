module fake_jpeg_8407_n_65 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_34),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_3),
.B(n_5),
.Y(n_38)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_9),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_7),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.C(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_55),
.B(n_49),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_48),
.B(n_53),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_46),
.B1(n_47),
.B2(n_43),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_51),
.C(n_52),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_45),
.Y(n_65)
);


endmodule