module fake_jpeg_19292_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_38),
.B1(n_24),
.B2(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_30),
.Y(n_94)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_84),
.B1(n_30),
.B2(n_24),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_34),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_22),
.B(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_83),
.Y(n_109)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_74),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_23),
.B1(n_21),
.B2(n_31),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_22),
.B1(n_28),
.B2(n_16),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_37),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_40),
.B1(n_35),
.B2(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_111),
.B1(n_24),
.B2(n_18),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_27),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_101),
.B(n_103),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_80),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_27),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_20),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_18),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_28),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_29),
.C(n_20),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_29),
.C(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_115),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_138),
.C(n_139),
.Y(n_150)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_82),
.B1(n_57),
.B2(n_72),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_124),
.B1(n_136),
.B2(n_77),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_129),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_132),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_70),
.B1(n_59),
.B2(n_23),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_131),
.Y(n_153)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_61),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_15),
.B1(n_21),
.B2(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_70),
.B1(n_59),
.B2(n_23),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_91),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_61),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_73),
.B(n_1),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_117),
.B(n_118),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_141),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_152),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_103),
.A3(n_101),
.B1(n_91),
.B2(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_147),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_0),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_101),
.C(n_86),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_155),
.C(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_87),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_96),
.C(n_88),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_162),
.B(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_163),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_96),
.C(n_92),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_95),
.B(n_15),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_172),
.B(n_144),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_111),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_90),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_90),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_117),
.A2(n_98),
.B1(n_110),
.B2(n_89),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_170),
.B1(n_140),
.B2(n_29),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_77),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_58),
.B1(n_15),
.B2(n_28),
.Y(n_169)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_95),
.B1(n_29),
.B2(n_20),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_73),
.B(n_1),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_161),
.B(n_143),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_194),
.B(n_157),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_204),
.B1(n_205),
.B2(n_166),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_190),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_25),
.B1(n_20),
.B2(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_0),
.Y(n_227)
);

XOR2x2_ASAP7_75t_SL g189 ( 
.A(n_146),
.B(n_25),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_167),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_154),
.A2(n_26),
.B1(n_17),
.B2(n_2),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_26),
.B1(n_17),
.B2(n_2),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_17),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_196),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_0),
.B(n_1),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_8),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_170),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_149),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_202),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_164),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_160),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_159),
.C(n_150),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_219),
.C(n_226),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_182),
.B(n_188),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_148),
.C(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_212),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_151),
.C(n_162),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_193),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_183),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_173),
.C(n_7),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_9),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_243),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_182),
.B1(n_198),
.B2(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_188),
.C(n_185),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_240),
.C(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_184),
.C(n_196),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_184),
.C(n_205),
.Y(n_241)
);

BUFx6f_ASAP7_75t_SL g242 ( 
.A(n_208),
.Y(n_242)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_221),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_217),
.B(n_208),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_256),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_228),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_212),
.C(n_215),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_258),
.C(n_244),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_213),
.C(n_211),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_176),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_231),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_229),
.A2(n_194),
.B(n_227),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_227),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_267),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_239),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_239),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_270),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_241),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_273),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_207),
.C(n_244),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_260),
.B1(n_255),
.B2(n_263),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_189),
.CI(n_181),
.CON(n_276),
.SN(n_276)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_278),
.B1(n_277),
.B2(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_181),
.C(n_195),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_186),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_204),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_252),
.B1(n_259),
.B2(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_284),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_2),
.C(n_3),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_255),
.B1(n_261),
.B2(n_276),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_286),
.B(n_289),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_260),
.B(n_190),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_191),
.B(n_10),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_6),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_10),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_13),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_14),
.C(n_3),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_14),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_297),
.B(n_14),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_283),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_302),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_289),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_291),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_307),
.B(n_300),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_298),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_306),
.C(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_293),
.B(n_301),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_285),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_4),
.Y(n_313)
);


endmodule