module fake_aes_1306_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_7), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_11), .B(n_8), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g17 ( .A(n_9), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_0), .B(n_1), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
NAND3xp33_ASAP7_75t_SL g20 ( .A(n_18), .B(n_16), .C(n_14), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_20), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B(n_17), .Y(n_22) );
OAI21xp5_ASAP7_75t_SL g23 ( .A1(n_22), .A2(n_3), .B(n_4), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_5), .B1(n_10), .B2(n_12), .Y(n_26) );
endmodule