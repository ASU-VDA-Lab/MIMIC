module fake_aes_10469_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_11), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
INVxp67_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g19 ( .A(n_15), .B(n_0), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_1), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_22), .Y(n_23) );
NOR3xp33_ASAP7_75t_SL g24 ( .A(n_23), .B(n_19), .C(n_16), .Y(n_24) );
OAI222xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_13), .B1(n_17), .B2(n_1), .C1(n_2), .C2(n_21), .Y(n_25) );
BUFx6f_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI221xp5_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_2), .B1(n_14), .B2(n_5), .C(n_6), .Y(n_27) );
OAI222xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_26), .B1(n_7), .B2(n_9), .C1(n_3), .C2(n_14), .Y(n_28) );
INVxp67_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
endmodule