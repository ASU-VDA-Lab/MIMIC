module fake_jpeg_3051_n_388 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_49),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_8),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_56),
.Y(n_111)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_18),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_51),
.Y(n_124)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_54),
.B(n_62),
.Y(n_94)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_9),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_14),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_73),
.Y(n_126)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_75),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_81),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_7),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_84),
.B1(n_86),
.B2(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_10),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_46),
.B(n_10),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_10),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_13),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_50),
.B1(n_91),
.B2(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_37),
.B1(n_24),
.B2(n_23),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_119),
.B1(n_128),
.B2(n_75),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_122),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_21),
.B1(n_19),
.B2(n_27),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_118),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_21),
.B1(n_19),
.B2(n_27),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_45),
.B1(n_28),
.B2(n_37),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_52),
.A2(n_19),
.B1(n_27),
.B2(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_20),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_22),
.B1(n_45),
.B2(n_20),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_73),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_97),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_64),
.B1(n_89),
.B2(n_84),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_137),
.B1(n_136),
.B2(n_106),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_51),
.A2(n_41),
.B(n_39),
.C(n_35),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_76),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_86),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_51),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_139),
.B(n_140),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_150),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_82),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_76),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_146),
.A2(n_165),
.B1(n_174),
.B2(n_175),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_94),
.B(n_14),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_103),
.B(n_41),
.CI(n_63),
.CON(n_151),
.SN(n_151)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_157),
.Y(n_203)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

OR2x4_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_67),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_155),
.A2(n_156),
.B1(n_178),
.B2(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_13),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_99),
.A2(n_57),
.A3(n_53),
.B1(n_41),
.B2(n_63),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_11),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_11),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_168),
.Y(n_208)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_11),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_102),
.B1(n_131),
.B2(n_123),
.Y(n_205)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_1),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_177),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_132),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_105),
.A2(n_41),
.B1(n_25),
.B2(n_18),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_95),
.B1(n_100),
.B2(n_129),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_191),
.B1(n_193),
.B2(n_202),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_93),
.B1(n_110),
.B2(n_104),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_115),
.B1(n_105),
.B2(n_126),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_117),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_151),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_171),
.B1(n_146),
.B2(n_164),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_153),
.B(n_145),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_143),
.A2(n_155),
.B(n_151),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_161),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_215),
.B(n_217),
.Y(n_252)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_138),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_233),
.B1(n_205),
.B2(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_228),
.Y(n_250)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_227),
.Y(n_237)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_167),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_234),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_126),
.B1(n_116),
.B2(n_98),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_203),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_206),
.B(n_201),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_232),
.B(n_196),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_181),
.B1(n_186),
.B2(n_183),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_242),
.B1(n_222),
.B2(n_219),
.Y(n_266)
);

OAI22x1_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_201),
.B1(n_209),
.B2(n_183),
.Y(n_241)
);

AOI22x1_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_226),
.B1(n_233),
.B2(n_228),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_193),
.B1(n_203),
.B2(n_185),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_256),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_253),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_234),
.A2(n_209),
.B1(n_201),
.B2(n_185),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_252),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_258),
.B(n_260),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_261),
.B(n_249),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_213),
.C(n_192),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_272),
.C(n_277),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_204),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

AOI22x1_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_222),
.B1(n_211),
.B2(n_214),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_268),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_255),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_222),
.B1(n_220),
.B2(n_224),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_204),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_273),
.C(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_222),
.B1(n_184),
.B2(n_229),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_249),
.B1(n_237),
.B2(n_225),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_180),
.C(n_198),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_184),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_208),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_195),
.Y(n_292)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_276),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_180),
.C(n_198),
.Y(n_277)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_253),
.B(n_246),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g309 ( 
.A(n_279),
.B(n_194),
.C(n_131),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_187),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_255),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_259),
.B(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_231),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_289),
.C(n_294),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_257),
.A2(n_237),
.B1(n_256),
.B2(n_236),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_290),
.B1(n_268),
.B2(n_271),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_237),
.C(n_195),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_257),
.A2(n_236),
.B1(n_251),
.B2(n_218),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_275),
.C(n_266),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_257),
.B1(n_259),
.B2(n_265),
.Y(n_298)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_315),
.B(n_290),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_294),
.B1(n_292),
.B2(n_289),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_174),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_251),
.B1(n_227),
.B2(n_190),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_303),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_148),
.B1(n_116),
.B2(n_188),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_282),
.A2(n_194),
.B1(n_114),
.B2(n_178),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_114),
.B1(n_152),
.B2(n_170),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_175),
.B(n_176),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_291),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_327),
.Y(n_336)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_313),
.A3(n_299),
.B1(n_304),
.B2(n_308),
.C1(n_300),
.C2(n_298),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_321),
.A2(n_331),
.B(n_127),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_301),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_329),
.Y(n_339)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_281),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_283),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_134),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_280),
.C(n_286),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_332),
.Y(n_341)
);

AOI321xp33_ASAP7_75t_L g331 ( 
.A1(n_305),
.A2(n_280),
.A3(n_134),
.B1(n_177),
.B2(n_123),
.C(n_169),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_158),
.C(n_141),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_315),
.C(n_307),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_335),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_316),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_310),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_338),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_306),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_13),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_323),
.B(n_12),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_343),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_324),
.B(n_319),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_344),
.A2(n_331),
.B(n_324),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_317),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_339),
.A2(n_333),
.B1(n_318),
.B2(n_320),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_357),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_358),
.C(n_25),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_354),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_334),
.A2(n_325),
.B1(n_333),
.B2(n_320),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_355),
.B(n_336),
.Y(n_360)
);

FAx1_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_319),
.CI(n_332),
.CON(n_354),
.SN(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_345),
.A2(n_134),
.B(n_177),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_12),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_120),
.C(n_132),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_349),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_363),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_367),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_338),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_362),
.A2(n_365),
.B(n_366),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_356),
.B(n_346),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_120),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_132),
.B(n_25),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_354),
.A2(n_18),
.B(n_3),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_SL g369 ( 
.A(n_368),
.B(n_354),
.C(n_358),
.Y(n_369)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_351),
.C(n_4),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_372),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_364),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_1),
.B(n_4),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_374),
.A2(n_6),
.B(n_371),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_375),
.A2(n_1),
.B(n_4),
.Y(n_377)
);

AOI21xp33_ASAP7_75t_L g382 ( 
.A1(n_377),
.A2(n_379),
.B(n_376),
.Y(n_382)
);

OAI21x1_ASAP7_75t_SL g378 ( 
.A1(n_375),
.A2(n_4),
.B(n_5),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_380),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_373),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_6),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_381),
.C(n_6),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_385),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_387),
.Y(n_388)
);


endmodule