module real_jpeg_546_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_0),
.B(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_1),
.B(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

AO21x2_ASAP7_75t_L g9 ( 
.A1(n_3),
.A2(n_10),
.B(n_11),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_20),
.Y(n_19)
);

NAND2x1_ASAP7_75t_SL g21 ( 
.A(n_4),
.B(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_12),
.B(n_22),
.C(n_32),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_9),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_16),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_17),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_16),
.A2(n_17),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_21),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_35),
.B(n_36),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);


endmodule