module real_jpeg_16338_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_382),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_0),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_2),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_2),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_2),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_2),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_2),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_2),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

NAND2x1_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_74),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_3),
.B(n_79),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_3),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_3),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_4),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_5),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_5),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_5),
.B(n_113),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_9),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_9),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_9),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_9),
.B(n_181),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_9),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_9),
.B(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_12),
.Y(n_383)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_163),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_162),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_19),
.B(n_139),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_90),
.C(n_117),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_20),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.C(n_84),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_21),
.B(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.C(n_45),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_22),
.B(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_23),
.A2(n_33),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.Y(n_23)
);

NAND2x1p5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_24),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_102),
.C(n_105),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_24),
.A2(n_86),
.B1(n_102),
.B2(n_103),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_24),
.A2(n_86),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_27),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_37),
.B(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_31),
.C(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_28),
.A2(n_230),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_28),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_28),
.A2(n_37),
.B1(n_236),
.B2(n_242),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_30),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_30),
.B(n_31),
.C(n_200),
.Y(n_283)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_31),
.A2(n_34),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_31),
.A2(n_34),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_33),
.A2(n_173),
.B(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_34),
.B(n_70),
.C(n_94),
.Y(n_93)
);

XOR2x1_ASAP7_75t_L g344 ( 
.A(n_35),
.B(n_45),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_36),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_37),
.A2(n_174),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_37),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_37),
.A2(n_66),
.B1(n_242),
.B2(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_37),
.B(n_66),
.C(n_213),
.Y(n_310)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_41),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_41),
.B(n_330),
.Y(n_329)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_58),
.Y(n_45)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_47),
.A2(n_48),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_47),
.A2(n_48),
.B1(n_102),
.B2(n_103),
.Y(n_208)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_48),
.B(n_53),
.C(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_48),
.B(n_88),
.C(n_122),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_48),
.A2(n_103),
.B(n_185),
.C(n_244),
.Y(n_268)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_57),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_58),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_58),
.B(n_156),
.C(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_58),
.A2(n_73),
.B1(n_134),
.B2(n_156),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_58),
.A2(n_134),
.B1(n_200),
.B2(n_203),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_106),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_59),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_63),
.B(n_84),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_77),
.C(n_80),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_64),
.A2(n_65),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.C(n_73),
.Y(n_65)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_66),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_66),
.A2(n_73),
.B1(n_156),
.B2(n_272),
.Y(n_333)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_70),
.A2(n_94),
.B1(n_95),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_70),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_70),
.A2(n_138),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_70),
.B(n_81),
.C(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_73),
.A2(n_110),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_73),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_73),
.B(n_116),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_73),
.A2(n_158),
.B(n_159),
.Y(n_331)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_77),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_77),
.B(n_81),
.Y(n_324)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_78),
.B(n_216),
.C(n_305),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_80),
.A2(n_81),
.B1(n_319),
.B2(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_85),
.C(n_88),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_81),
.B(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_81),
.B(n_319),
.C(n_321),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_86),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_89),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_88),
.A2(n_89),
.B1(n_109),
.B2(n_115),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_88),
.B(n_103),
.C(n_110),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_90),
.B(n_117),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_108),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_100),
.B2(n_101),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_101),
.C(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_102),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_102),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_102),
.B(n_251),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_104),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_130),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_105),
.A2(n_278),
.B(n_282),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_105),
.B(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_112),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_R g240 ( 
.A1(n_110),
.A2(n_180),
.B(n_241),
.C(n_244),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_110),
.B(n_180),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_110),
.A2(n_155),
.B1(n_180),
.B2(n_182),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_110),
.A2(n_155),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_155),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_128),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_127),
.C(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.C(n_135),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_129),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_133),
.B(n_135),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_134),
.B(n_203),
.C(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_138),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_161),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_151),
.B1(n_152),
.B2(n_160),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_376),
.B(n_380),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI321xp33_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_313),
.A3(n_364),
.B1(n_369),
.B2(n_370),
.C(n_375),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_285),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_261),
.B(n_284),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_220),
.B(n_260),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_195),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_195),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_183),
.C(n_188),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_183),
.A2(n_188),
.B1(n_189),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_185),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_185),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_192),
.A2(n_213),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_204),
.B2(n_205),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_198),
.B(n_204),
.C(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_211),
.C(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_216),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_216),
.A2(n_219),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_229),
.B(n_230),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_238),
.B(n_259),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_225),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.C(n_234),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_248),
.B(n_258),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_245),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_255),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_254),
.B(n_257),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.B(n_253),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_274),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.C(n_274),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_270),
.C(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_283),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_277),
.C(n_283),
.Y(n_312)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_282),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_286),
.B(n_287),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_288),
.B(n_301),
.C(n_312),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_298),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_294),
.C(n_298),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_310),
.C(n_311),
.Y(n_336)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_352),
.Y(n_313)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_345),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_315),
.B(n_345),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_334),
.C(n_342),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_343),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_327),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_322),
.B1(n_325),
.B2(n_326),
.Y(n_317)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_326),
.C(n_327),
.Y(n_346)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.C(n_332),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

XOR2x2_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.C(n_338),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_348),
.C(n_350),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

AOI31xp67_ASAP7_75t_L g370 ( 
.A1(n_352),
.A2(n_365),
.A3(n_371),
.B(n_374),
.Y(n_370)
);

NAND2x1p5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

NOR2x1_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_355),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.C(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_361),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_368),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

AND2x4_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_378),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);


endmodule