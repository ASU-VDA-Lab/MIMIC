module fake_jpeg_15535_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_8),
.B(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_52),
.Y(n_90)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_49),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_3),
.C(n_4),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_5),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_6),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_7),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_35),
.B1(n_36),
.B2(n_28),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_74),
.B1(n_87),
.B2(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_35),
.B1(n_36),
.B2(n_28),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_20),
.B(n_29),
.C(n_22),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_34),
.B1(n_29),
.B2(n_22),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_79),
.B1(n_83),
.B2(n_88),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_17),
.B1(n_34),
.B2(n_16),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_42),
.A2(n_21),
.B1(n_33),
.B2(n_30),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_43),
.A2(n_21),
.B1(n_30),
.B2(n_11),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_21),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_10),
.B(n_11),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_80),
.B(n_81),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_44),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_50),
.B1(n_71),
.B2(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_117),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_13),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_124),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_54),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_123),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_45),
.CON(n_113),
.SN(n_113)
);

NOR4xp25_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_131),
.C(n_123),
.D(n_118),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_48),
.B(n_50),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_127),
.C(n_130),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_48),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_103),
.B1(n_78),
.B2(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_101),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_66),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_72),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_73),
.B(n_94),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_66),
.A2(n_78),
.B(n_67),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_135),
.A2(n_95),
.B1(n_130),
.B2(n_134),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_140),
.B1(n_146),
.B2(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_95),
.B1(n_103),
.B2(n_112),
.Y(n_140)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_108),
.CI(n_106),
.CON(n_174),
.SN(n_174)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_122),
.B1(n_115),
.B2(n_110),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_128),
.B1(n_132),
.B2(n_106),
.Y(n_170)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_158),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_108),
.Y(n_172)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_110),
.C(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_114),
.C(n_126),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_169),
.B1(n_181),
.B2(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_114),
.B1(n_105),
.B2(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_127),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_174),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_105),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_179),
.C(n_180),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_117),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_177),
.B(n_182),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_143),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_129),
.C(n_135),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_135),
.B1(n_104),
.B2(n_129),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_156),
.B(n_139),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_194),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_192),
.Y(n_206)
);

AOI211xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_139),
.B(n_149),
.C(n_140),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_144),
.A3(n_174),
.B1(n_148),
.B2(n_154),
.C1(n_181),
.C2(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_159),
.B(n_161),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_137),
.B1(n_150),
.B2(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_197),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_144),
.B1(n_136),
.B2(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_169),
.Y(n_203)
);

AO221x1_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_178),
.B1(n_168),
.B2(n_142),
.C(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_173),
.C(n_179),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_202),
.C(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_172),
.C(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_185),
.B1(n_199),
.B2(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_187),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_208),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_144),
.A3(n_104),
.B1(n_168),
.B2(n_142),
.C1(n_135),
.C2(n_153),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_153),
.B(n_157),
.C(n_198),
.D(n_193),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_194),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_218),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_210),
.C(n_203),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_198),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_219),
.C(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_222),
.C(n_225),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_211),
.C(n_207),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_209),
.B(n_211),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_204),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_227),
.B(n_228),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_210),
.B(n_215),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_184),
.A3(n_191),
.B1(n_214),
.B2(n_185),
.C1(n_195),
.C2(n_219),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_233),
.B(n_212),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_184),
.B(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_188),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_235),
.B1(n_189),
.B2(n_229),
.C(n_217),
.Y(n_236)
);


endmodule