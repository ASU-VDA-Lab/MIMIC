module real_jpeg_6534_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_1),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_63),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_1),
.A2(n_63),
.B1(n_109),
.B2(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_3),
.A2(n_136),
.B1(n_265),
.B2(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_3),
.A2(n_69),
.B1(n_136),
.B2(n_286),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_3),
.A2(n_136),
.B1(n_227),
.B2(n_363),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_4),
.A2(n_54),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_4),
.A2(n_54),
.B1(n_212),
.B2(n_287),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_182),
.B1(n_183),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_6),
.Y(n_100)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_7),
.Y(n_219)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_7),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_8),
.A2(n_72),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_9),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_10),
.Y(n_103)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_11),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_122),
.B1(n_163),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_12),
.A2(n_122),
.B1(n_174),
.B2(n_271),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_12),
.A2(n_69),
.B1(n_122),
.B2(n_212),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_13),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_13),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_13),
.A2(n_162),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_13),
.A2(n_162),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_13),
.A2(n_162),
.B1(n_265),
.B2(n_334),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_14),
.A2(n_86),
.B1(n_237),
.B2(n_241),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_16),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_16),
.A2(n_203),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_16),
.B(n_277),
.C(n_280),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_16),
.B(n_111),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_16),
.B(n_180),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_16),
.B(n_56),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_16),
.B(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_255),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_254),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_231),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_21),
.B(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.C(n_187),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_22),
.A2(n_23),
.B1(n_166),
.B2(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_91),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_24),
.B(n_92),
.C(n_165),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_67),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_25),
.B(n_67),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_52),
.B1(n_55),
.B2(n_57),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_26),
.A2(n_264),
.B(n_269),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_26),
.A2(n_55),
.B1(n_297),
.B2(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_26),
.A2(n_269),
.B(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_27),
.A2(n_56),
.B1(n_58),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_27),
.A2(n_56),
.B1(n_168),
.B2(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_27),
.B(n_270),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_42),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_31),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_31),
.Y(n_265)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_31),
.Y(n_273)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_40),
.Y(n_242)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_42),
.A2(n_297),
.B(n_299),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_47),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_50),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_52),
.A2(n_55),
.B(n_299),
.Y(n_392)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_56),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_75),
.B1(n_81),
.B2(n_89),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_68),
.Y(n_220)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_71),
.Y(n_185)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_75),
.B(n_293),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_75),
.A2(n_218),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_75),
.A2(n_210),
.B1(n_347),
.B2(n_370),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_77),
.Y(n_244)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_82),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_176)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_85),
.Y(n_213)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_85),
.Y(n_290)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_131),
.B1(n_164),
.B2(n_165),
.Y(n_91)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

AOI22x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_111),
.B1(n_117),
.B2(n_126),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_93),
.A2(n_222),
.B(n_229),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_93),
.A2(n_229),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_93),
.B(n_117),
.Y(n_366)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_94),
.A2(n_127),
.B1(n_230),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_94),
.A2(n_223),
.B1(n_230),
.B2(n_362),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_111),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_101),
.B1(n_104),
.B2(n_108),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_103),
.Y(n_343)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_109),
.A2(n_203),
.B(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_110),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_111),
.Y(n_230)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g348 ( 
.A1(n_115),
.A2(n_265),
.A3(n_339),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_116),
.Y(n_351)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_118),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_125),
.Y(n_251)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_140),
.B1(n_151),
.B2(n_159),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_132),
.A2(n_190),
.B(n_192),
.Y(n_189)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_140),
.A2(n_159),
.B(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_141),
.A2(n_387),
.B(n_389),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_151),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_198),
.A3(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_197)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_151),
.B(n_203),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_157),
.Y(n_151)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g349 ( 
.A(n_156),
.Y(n_349)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_166),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_176),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_167),
.B(n_176),
.Y(n_247)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_172),
.Y(n_298)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_209),
.B1(n_217),
.B2(n_220),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_177),
.A2(n_181),
.B(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_177),
.A2(n_285),
.B(n_291),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_177),
.A2(n_203),
.B(n_291),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_180),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_187),
.B(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.C(n_221),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_188),
.A2(n_189),
.B1(n_221),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_191),
.B(n_193),
.Y(n_253)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_196),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_207),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_197),
.A2(n_207),
.B1(n_208),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_197),
.Y(n_380)
);

OAI21xp33_ASAP7_75t_SL g387 ( 
.A1(n_202),
.A2(n_203),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_217),
.A2(n_316),
.B(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_221),
.Y(n_402)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_230),
.A2(n_362),
.B(n_366),
.Y(n_361)
);

BUFx24_ASAP7_75t_SL g417 ( 
.A(n_231),
.Y(n_417)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.CI(n_246),
.CON(n_231),
.SN(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_243),
.B2(n_245),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_253),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_395),
.B(n_414),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_375),
.B(n_394),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_353),
.B(n_374),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_327),
.B(n_352),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_302),
.B(n_326),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_283),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_262),
.B(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_274),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_263),
.A2(n_274),
.B1(n_275),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_294),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_295),
.C(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_300),
.B2(n_301),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp33_ASAP7_75t_SL g350 ( 
.A(n_298),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_319),
.B(n_325),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_312),
.B(n_318),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_317),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_329),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_344),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_335),
.B2(n_336),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_335),
.C(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_348),
.Y(n_359)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_354),
.B(n_355),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_360),
.B2(n_373),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_359),
.C(n_373),
.Y(n_376)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_367),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_368),
.C(n_369),
.Y(n_381)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_376),
.B(n_377),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_384),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_378)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_382),
.C(n_384),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_390),
.B2(n_393),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_391),
.C(n_392),
.Y(n_405)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_390),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_409),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_415),
.B(n_416),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_406),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_406),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.C(n_405),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_403),
.A2(n_404),
.B1(n_405),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_405),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_411),
.Y(n_415)
);


endmodule