module fake_jpeg_14095_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx4f_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx24_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_1),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_20),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_13),
.A3(n_10),
.B1(n_8),
.B2(n_7),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_13),
.B1(n_10),
.B2(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_32),
.B1(n_24),
.B2(n_30),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_18),
.B1(n_16),
.B2(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_37),
.B(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_23),
.C(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_42),
.C(n_43),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_24),
.C(n_21),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_30),
.C(n_25),
.Y(n_43)
);

BUFx24_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_37),
.C(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_18),
.B1(n_34),
.B2(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_6),
.B1(n_2),
.B2(n_4),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_1),
.B1(n_5),
.B2(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_5),
.C(n_51),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_49),
.B(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);


endmodule