module fake_jpeg_15255_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_44),
.Y(n_52)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_1),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_31),
.B1(n_26),
.B2(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_21),
.B1(n_26),
.B2(n_29),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_61),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_21),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_39),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_33),
.B1(n_25),
.B2(n_27),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_19),
.B1(n_30),
.B2(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_44),
.B1(n_39),
.B2(n_36),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_68),
.B1(n_79),
.B2(n_2),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_85),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_43),
.B1(n_37),
.B2(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_76),
.Y(n_99)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_81),
.B1(n_32),
.B2(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_88),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_27),
.B1(n_19),
.B2(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_60),
.B1(n_18),
.B2(n_53),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_16),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_2),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_73),
.B1(n_71),
.B2(n_70),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_77),
.C(n_89),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_34),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_110),
.C(n_34),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_3),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_16),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_32),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_111),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_83),
.C(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_72),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_82),
.B(n_76),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_98),
.B1(n_90),
.B2(n_96),
.C(n_95),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_103),
.B1(n_93),
.B2(n_6),
.Y(n_143)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_128),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_109),
.B1(n_107),
.B2(n_94),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_124),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_133),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_34),
.B(n_41),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_53),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_126),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_135),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_143),
.B(n_118),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_93),
.C(n_94),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_113),
.Y(n_152)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_127),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_120),
.B1(n_116),
.B2(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_151),
.C(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_158),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_115),
.B1(n_116),
.B2(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_162),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_115),
.B1(n_130),
.B2(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_165),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_147),
.B(n_137),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_124),
.B1(n_121),
.B2(n_128),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_151),
.C(n_137),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_32),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_171),
.C(n_80),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_143),
.C(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_153),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_135),
.B(n_144),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_163),
.B1(n_158),
.B2(n_80),
.Y(n_180)
);

AOI321xp33_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_146),
.A3(n_14),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_162),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_179),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_180),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_184),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_7),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_167),
.B(n_172),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_189),
.B(n_190),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_167),
.B1(n_172),
.B2(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_4),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_53),
.C(n_8),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_194),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_195),
.B(n_15),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_12),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_15),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_196),
.B(n_5),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule