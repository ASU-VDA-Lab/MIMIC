module fake_jpeg_22237_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_49),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_20),
.C(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_34),
.B1(n_37),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_73),
.B1(n_23),
.B2(n_20),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_34),
.B1(n_37),
.B2(n_22),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_36),
.B1(n_23),
.B2(n_20),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_69),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_34),
.B1(n_24),
.B2(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_37),
.B1(n_22),
.B2(n_23),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_35),
.B1(n_25),
.B2(n_29),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_84),
.A2(n_111),
.B1(n_55),
.B2(n_8),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_26),
.B1(n_24),
.B2(n_32),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_91),
.B1(n_108),
.B2(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_92),
.B1(n_61),
.B2(n_51),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_36),
.B1(n_31),
.B2(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_97),
.Y(n_150)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_35),
.B1(n_25),
.B2(n_29),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_117),
.B1(n_71),
.B2(n_27),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_103),
.Y(n_148)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_105),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_63),
.B(n_57),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_61),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_26),
.B1(n_24),
.B2(n_32),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_31),
.B1(n_18),
.B2(n_19),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_83),
.B1(n_82),
.B2(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_38),
.B1(n_17),
.B2(n_29),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_35),
.B1(n_25),
.B2(n_27),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_38),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_0),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_27),
.B1(n_38),
.B2(n_9),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_127),
.B1(n_142),
.B2(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_69),
.C(n_65),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_124),
.B(n_129),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_75),
.B1(n_53),
.B2(n_54),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_38),
.B1(n_55),
.B2(n_51),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_86),
.B1(n_94),
.B2(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_133),
.B(n_141),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_61),
.C(n_64),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_149),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_61),
.A3(n_59),
.B1(n_55),
.B2(n_51),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_136),
.B(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_59),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_96),
.B1(n_97),
.B2(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_86),
.A2(n_94),
.B1(n_114),
.B2(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_164),
.Y(n_202)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_152),
.B1(n_120),
.B2(n_138),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_165),
.B1(n_171),
.B2(n_177),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_119),
.B1(n_115),
.B2(n_105),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_113),
.B1(n_98),
.B2(n_2),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_180),
.B1(n_151),
.B2(n_128),
.Y(n_215)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_173),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_182),
.B(n_150),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_175),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_147),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_179),
.B1(n_187),
.B2(n_131),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_5),
.B1(n_16),
.B2(n_7),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_137),
.B(n_6),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_10),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_7),
.B(n_9),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_136),
.B1(n_120),
.B2(n_126),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_129),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_192),
.B(n_206),
.Y(n_243)
);

CKINVDCx6p67_ASAP7_75t_R g189 ( 
.A(n_175),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_149),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_127),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_140),
.Y(n_207)
);

OAI31xp33_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_168),
.A3(n_164),
.B(n_158),
.Y(n_221)
);

INVx6_ASAP7_75t_SL g208 ( 
.A(n_175),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_15),
.B(n_11),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_145),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_218),
.C(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_183),
.B1(n_171),
.B2(n_178),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_153),
.B(n_123),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_160),
.A2(n_140),
.B(n_11),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_225),
.B(n_231),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_163),
.B1(n_166),
.B2(n_183),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_233),
.B1(n_234),
.B2(n_238),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_170),
.B(n_157),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_195),
.B1(n_216),
.B2(n_210),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_163),
.B1(n_180),
.B2(n_157),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_177),
.B1(n_181),
.B2(n_168),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_189),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_177),
.B(n_174),
.C(n_176),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_201),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_177),
.B1(n_172),
.B2(n_182),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_239),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_195),
.B1(n_199),
.B2(n_204),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_14),
.C(n_15),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_213),
.C(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_252),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_243),
.B(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_240),
.B1(n_230),
.B2(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_212),
.C(n_194),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_249),
.C(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_200),
.C(n_205),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_206),
.C(n_196),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_232),
.B(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_189),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_236),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_208),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_197),
.C(n_241),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_238),
.C(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_234),
.B1(n_235),
.B2(n_220),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_266),
.A2(n_248),
.B1(n_220),
.B2(n_226),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_221),
.CI(n_234),
.CON(n_270),
.SN(n_270)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_246),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_224),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_276),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_279),
.C(n_244),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_264),
.B(n_274),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_222),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_263),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_258),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_291),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_262),
.B1(n_260),
.B2(n_248),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_228),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_279),
.C(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_295),
.C(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_302),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_272),
.C(n_269),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_285),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_227),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_219),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_219),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_302),
.C(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_319),
.C(n_297),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_296),
.B(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_272),
.A3(n_288),
.B1(n_283),
.B2(n_282),
.C1(n_287),
.C2(n_271),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_317),
.C(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_316),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.C(n_321),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_255),
.C(n_281),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_270),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_270),
.Y(n_328)
);


endmodule