module fake_jpeg_12553_n_365 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_365);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_365;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g149 ( 
.A(n_56),
.Y(n_149)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_19),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_83),
.Y(n_116)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_71),
.B(n_78),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_10),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_38),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_81),
.B(n_88),
.Y(n_167)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_87),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_27),
.B(n_2),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_93),
.Y(n_118)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_98),
.B(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_100),
.Y(n_143)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_49),
.B(n_37),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_28),
.B(n_3),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_108),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_32),
.B(n_4),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_107),
.B(n_60),
.Y(n_163)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_34),
.B(n_41),
.C(n_40),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_37),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_126),
.B(n_134),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_54),
.B1(n_41),
.B2(n_40),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_142),
.B1(n_134),
.B2(n_136),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_76),
.B1(n_35),
.B2(n_86),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_157),
.B1(n_138),
.B2(n_125),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_61),
.A2(n_54),
.B1(n_29),
.B2(n_23),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_136),
.B1(n_142),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_29),
.B1(n_39),
.B2(n_23),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_39),
.B1(n_21),
.B2(n_45),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_78),
.A2(n_107),
.B1(n_103),
.B2(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_159),
.B1(n_169),
.B2(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_52),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_158),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_94),
.A2(n_52),
.B1(n_49),
.B2(n_45),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_35),
.B1(n_0),
.B2(n_13),
.Y(n_151)
);

NOR2x1_ASAP7_75t_R g154 ( 
.A(n_81),
.B(n_4),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_154),
.B(n_160),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_87),
.A2(n_0),
.B1(n_13),
.B2(n_14),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_79),
.B(n_15),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_64),
.A2(n_84),
.B1(n_104),
.B2(n_56),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_168),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_102),
.A2(n_81),
.B(n_17),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_71),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_162),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_58),
.B(n_89),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_78),
.A2(n_107),
.B1(n_103),
.B2(n_98),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_174),
.B(n_189),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_175),
.B(n_182),
.Y(n_246)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_137),
.B1(n_113),
.B2(n_112),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_179),
.A2(n_184),
.B1(n_216),
.B2(n_188),
.Y(n_250)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_118),
.B(n_111),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_154),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_188),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_109),
.B1(n_153),
.B2(n_164),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_185),
.A2(n_187),
.B1(n_201),
.B2(n_204),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_151),
.B1(n_131),
.B2(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_124),
.B(n_123),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_197),
.Y(n_222)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_117),
.B(n_115),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_138),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_196),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_115),
.B(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_206),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_140),
.B1(n_153),
.B2(n_121),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_202),
.B(n_205),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_160),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_109),
.A2(n_121),
.B1(n_157),
.B2(n_145),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_140),
.A2(n_161),
.B1(n_135),
.B2(n_120),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_135),
.A2(n_132),
.B1(n_152),
.B2(n_156),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_145),
.A2(n_127),
.B1(n_152),
.B2(n_130),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_216),
.B1(n_202),
.B2(n_191),
.Y(n_244)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_130),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_211),
.Y(n_227)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_147),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_127),
.B(n_166),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_215),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g213 ( 
.A(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_139),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_174),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_163),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_129),
.A2(n_113),
.B1(n_137),
.B2(n_119),
.Y(n_216)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_135),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_149),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_220),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_201),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_173),
.B(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_200),
.C(n_199),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_172),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_233),
.B(n_240),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_179),
.B1(n_187),
.B2(n_177),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_244),
.B1(n_250),
.B2(n_209),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_170),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_200),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_196),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_196),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_250),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_272),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_219),
.B(n_205),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_267),
.B(n_248),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_171),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_204),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_265),
.C(n_275),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_199),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_195),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_199),
.B(n_206),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_221),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_239),
.B(n_218),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_239),
.B(n_192),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_274),
.A2(n_281),
.B1(n_282),
.B2(n_280),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_224),
.B(n_176),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_222),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_248),
.Y(n_291)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_221),
.B(n_210),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_217),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_237),
.A2(n_208),
.B1(n_190),
.B2(n_183),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_183),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_264),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_225),
.A2(n_183),
.B1(n_252),
.B2(n_235),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_248),
.B1(n_252),
.B2(n_236),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_267),
.B(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.Y(n_303)
);

AO22x1_ASAP7_75t_L g292 ( 
.A1(n_259),
.A2(n_236),
.B1(n_241),
.B2(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_294),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_238),
.B1(n_231),
.B2(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_297),
.Y(n_318)
);

AO22x1_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_227),
.B1(n_242),
.B2(n_253),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_258),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_256),
.B1(n_268),
.B2(n_276),
.C(n_260),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_302),
.B(n_289),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_277),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_306),
.C(n_308),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_275),
.C(n_269),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_275),
.C(n_257),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_312),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_313),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_275),
.C(n_265),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_287),
.B1(n_288),
.B2(n_294),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_256),
.A3(n_262),
.B1(n_272),
.B2(n_279),
.C1(n_281),
.C2(n_226),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_284),
.B1(n_290),
.B2(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_261),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_290),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_318),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_320),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_285),
.B(n_292),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_327),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_331),
.B1(n_307),
.B2(n_304),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_301),
.B1(n_288),
.B2(n_287),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_323),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_317),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_318),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_330),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_308),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_335),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_306),
.C(n_313),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_337),
.C(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_334),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_305),
.C(n_303),
.Y(n_337)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_338),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_346),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_333),
.C(n_336),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_329),
.B1(n_319),
.B2(n_331),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_335),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_347),
.B(n_324),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_350),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_345),
.A2(n_340),
.B(n_327),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_353),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_345),
.A2(n_324),
.B(n_320),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_SL g355 ( 
.A1(n_352),
.A2(n_321),
.B(n_343),
.C(n_320),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_322),
.Y(n_358)
);

AOI31xp67_ASAP7_75t_SL g356 ( 
.A1(n_352),
.A2(n_328),
.A3(n_329),
.B(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_356),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_359),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_354),
.C(n_344),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_362),
.A2(n_348),
.B(n_343),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_363),
.B(n_347),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_361),
.Y(n_365)
);


endmodule