module fake_ibex_946_n_3714 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_3714);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_3714;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_3456;
wire n_2687;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3211;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2924;
wire n_2456;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_3544;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_3558;
wire n_2751;
wire n_2785;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1395;
wire n_998;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3401;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_1400;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_3557;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_3398;
wire n_2376;
wire n_2476;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_3314;
wire n_961;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_991;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3269;
wire n_3029;
wire n_3609;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1348;
wire n_1289;
wire n_838;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_3216;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_3066;
wire n_2714;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2653;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3343;
wire n_3163;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_3225;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_3067;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2148;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_3056;
wire n_2453;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_3406;
wire n_2678;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_318),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_387),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_576),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_526),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_432),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_738),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_76),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_309),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_343),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_182),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_76),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_488),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_623),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_774),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_799),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_747),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_776),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_497),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_410),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_575),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_548),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_789),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_569),
.Y(n_825)
);

BUFx10_ASAP7_75t_L g826 ( 
.A(n_371),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_670),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_670),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_504),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_788),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_382),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_54),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_488),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_480),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_60),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_411),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_239),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_685),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_326),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_351),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_447),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_147),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_630),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_175),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_39),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_668),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_131),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_4),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_357),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_134),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_482),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_231),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_11),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_777),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_224),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_640),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_400),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_590),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_531),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_299),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_786),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_254),
.Y(n_862)
);

BUFx10_ASAP7_75t_L g863 ( 
.A(n_630),
.Y(n_863)
);

BUFx5_ASAP7_75t_L g864 ( 
.A(n_775),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_32),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_83),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_123),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_13),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_299),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_496),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_96),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_500),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_58),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_542),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_108),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_288),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_715),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_170),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_679),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_599),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_699),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_271),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_495),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_280),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_795),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_395),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_497),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_350),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_350),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_770),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_28),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_335),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_446),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_673),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_714),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_513),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_586),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_66),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_508),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_772),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_9),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_690),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_196),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_678),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_270),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_52),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_617),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_351),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_131),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_796),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_482),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_608),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_475),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_618),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_53),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_15),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_55),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_758),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_170),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_771),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_201),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_573),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_493),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_441),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_757),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_748),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_538),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_176),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_537),
.Y(n_929)
);

INVxp33_ASAP7_75t_L g930 ( 
.A(n_370),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_452),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_696),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_296),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_615),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_198),
.Y(n_935)
);

BUFx10_ASAP7_75t_L g936 ( 
.A(n_391),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_390),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_384),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_329),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_548),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_261),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_686),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_778),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_481),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_631),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_27),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_103),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_579),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_164),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_456),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_377),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_21),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_72),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_560),
.Y(n_954)
);

BUFx8_ASAP7_75t_SL g955 ( 
.A(n_769),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_199),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_133),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_515),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_85),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_2),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_125),
.Y(n_961)
);

INVxp33_ASAP7_75t_R g962 ( 
.A(n_614),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_363),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_3),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_366),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_67),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_133),
.Y(n_967)
);

BUFx8_ASAP7_75t_SL g968 ( 
.A(n_429),
.Y(n_968)
);

BUFx5_ASAP7_75t_L g969 ( 
.A(n_75),
.Y(n_969)
);

BUFx5_ASAP7_75t_L g970 ( 
.A(n_232),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_426),
.Y(n_971)
);

BUFx8_ASAP7_75t_SL g972 ( 
.A(n_1),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_317),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_669),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_419),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_231),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_430),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_101),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_457),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_587),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_320),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_204),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_292),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_84),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_694),
.Y(n_985)
);

CKINVDCx14_ASAP7_75t_R g986 ( 
.A(n_741),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_434),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_355),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_71),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_536),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_582),
.Y(n_991)
);

INVx4_ASAP7_75t_R g992 ( 
.A(n_584),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_179),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_111),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_55),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_787),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_561),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_645),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_174),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_235),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_271),
.Y(n_1001)
);

BUFx2_ASAP7_75t_SL g1002 ( 
.A(n_654),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_594),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_780),
.Y(n_1004)
);

CKINVDCx14_ASAP7_75t_R g1005 ( 
.A(n_742),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_469),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_665),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_584),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_664),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_210),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_650),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_592),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_81),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_545),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_5),
.Y(n_1015)
);

CKINVDCx16_ASAP7_75t_R g1016 ( 
.A(n_704),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_297),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_703),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_3),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_187),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_552),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_334),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_293),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_752),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_115),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_688),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_622),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_298),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_139),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_131),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_540),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_61),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_227),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_61),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_595),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_554),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_674),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_226),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_689),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_336),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_642),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_546),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_633),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_57),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_570),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_729),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_49),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_184),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_161),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_787),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_356),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_349),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_296),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_786),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_619),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_402),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_286),
.Y(n_1057)
);

BUFx10_ASAP7_75t_L g1058 ( 
.A(n_43),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_287),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_335),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_419),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_649),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_653),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_732),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_124),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_228),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_719),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_717),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_767),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_185),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_795),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_234),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_465),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_525),
.Y(n_1074)
);

BUFx5_ASAP7_75t_L g1075 ( 
.A(n_406),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_93),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_367),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_439),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_281),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_699),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_610),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_583),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_627),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_40),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_572),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_29),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_147),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_417),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_658),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_605),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_189),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_779),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_572),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_451),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_798),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_774),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_379),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_775),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_782),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_613),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_267),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_691),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_164),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_546),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_328),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_325),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_15),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_401),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_480),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_513),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_364),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_396),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_104),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_263),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_362),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_118),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_695),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_124),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_388),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_327),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_462),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_81),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_387),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_440),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_161),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_579),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_265),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_473),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_535),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_7),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_18),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_6),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_425),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_617),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_405),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_783),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_773),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_279),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_376),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_319),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_562),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_523),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_255),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_353),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_646),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_790),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_354),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_273),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_222),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_557),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_715),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_324),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_452),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_498),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_217),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_631),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_38),
.Y(n_1157)
);

BUFx8_ASAP7_75t_SL g1158 ( 
.A(n_691),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_641),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_429),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_367),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_680),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_322),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_742),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_186),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_644),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_788),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_286),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_674),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_784),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_29),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_494),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_230),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_545),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_694),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_781),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_37),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_197),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_486),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_408),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_785),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_171),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_81),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_544),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_708),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_647),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_739),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_972),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_972),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_935),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_915),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_986),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_949),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_986),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1005),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1005),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_955),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1084),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_853),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_812),
.B(n_0),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1183),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_907),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_955),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_851),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_842),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_853),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_866),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_867),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_968),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_875),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_969),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1039),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_898),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_875),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_903),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_968),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_966),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1158),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_930),
.B(n_0),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_848),
.Y(n_1220)
);

INVxp33_ASAP7_75t_SL g1221 ( 
.A(n_1155),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_813),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_832),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_969),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_835),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_966),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_917),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_844),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_919),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_845),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_847),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1025),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_993),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_858),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_873),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_865),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_850),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1025),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1020),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1118),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_868),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1030),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_930),
.B(n_1),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1032),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_871),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_850),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_878),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_850),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1070),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1107),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_891),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_809),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1003),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_969),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_959),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1113),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_901),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1021),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_909),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1118),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_947),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_820),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1126),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_947),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_916),
.Y(n_1265)
);

CKINVDCx16_ASAP7_75t_R g1266 ( 
.A(n_947),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_921),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_951),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_928),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1016),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_959),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1191),
.B(n_1198),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1237),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1220),
.Y(n_1274)
);

INVx5_ASAP7_75t_L g1275 ( 
.A(n_1246),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1222),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1252),
.Y(n_1277)
);

AND2x6_ASAP7_75t_L g1278 ( 
.A(n_1264),
.B(n_978),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1235),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1201),
.B(n_1136),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1248),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1190),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1202),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1255),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1271),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1224),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1205),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1224),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1254),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1261),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1223),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1207),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1208),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1213),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1215),
.B(n_969),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1253),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1266),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1219),
.A2(n_1182),
.B1(n_952),
.B2(n_953),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1204),
.B(n_1139),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1227),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1234),
.B(n_958),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1229),
.A2(n_961),
.B(n_960),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1225),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1263),
.B(n_1212),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1233),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_SL g1306 ( 
.A(n_1192),
.B(n_946),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1239),
.B(n_1242),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1244),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1252),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1249),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1188),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1250),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1228),
.B(n_956),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1230),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1256),
.A2(n_961),
.B(n_960),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1258),
.B(n_1117),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1231),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1252),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1226),
.A2(n_822),
.B1(n_823),
.B2(n_816),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1243),
.B(n_978),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1243),
.B(n_1165),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1221),
.B(n_1165),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1236),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1200),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1200),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1241),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1245),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1247),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1251),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1257),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1259),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1265),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1267),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1269),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1194),
.B(n_1195),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1196),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1193),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1197),
.A2(n_994),
.B(n_967),
.Y(n_1338)
);

INVx5_ASAP7_75t_L g1339 ( 
.A(n_1203),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1209),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1193),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1216),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1218),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1262),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1268),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1270),
.B(n_956),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1189),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1199),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1206),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1210),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1214),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1217),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1232),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1260),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1226),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1238),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1238),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1240),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1240),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1220),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1246),
.B(n_957),
.Y(n_1361)
);

CKINVDCx16_ASAP7_75t_R g1362 ( 
.A(n_1246),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1252),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1220),
.B(n_864),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1220),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1191),
.B(n_1149),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1220),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1220),
.B(n_864),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1220),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1220),
.B(n_864),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1220),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1220),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1220),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1220),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1264),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1220),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1246),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1211),
.A2(n_994),
.B(n_967),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1246),
.B(n_957),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1220),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1222),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1246),
.B(n_957),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1222),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1191),
.B(n_1161),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1220),
.B(n_864),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1246),
.B(n_1058),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1252),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1220),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1201),
.A2(n_816),
.B1(n_823),
.B2(n_822),
.Y(n_1389)
);

CKINVDCx6p67_ASAP7_75t_R g1390 ( 
.A(n_1246),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1237),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1264),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1237),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1220),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1220),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1211),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1252),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1220),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1246),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1220),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1246),
.B(n_1058),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1220),
.B(n_864),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1237),
.B(n_933),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1211),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1220),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1246),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1252),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_L g1408 ( 
.A(n_1278),
.B(n_1375),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1275),
.Y(n_1409)
);

NAND2x1_ASAP7_75t_L g1410 ( 
.A(n_1302),
.B(n_992),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_SL g1411 ( 
.A(n_1375),
.B(n_1028),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1305),
.B(n_1048),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1305),
.B(n_1177),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1296),
.Y(n_1414)
);

AND2x2_ASAP7_75t_SL g1415 ( 
.A(n_1362),
.B(n_1077),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1312),
.B(n_1178),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1275),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1278),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1390),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1392),
.B(n_1049),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1302),
.Y(n_1421)
);

AND2x6_ASAP7_75t_L g1422 ( 
.A(n_1361),
.B(n_1382),
.Y(n_1422)
);

INVx4_ASAP7_75t_SL g1423 ( 
.A(n_1278),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1392),
.Y(n_1424)
);

INVx8_ASAP7_75t_L g1425 ( 
.A(n_1401),
.Y(n_1425)
);

INVx4_ASAP7_75t_L g1426 ( 
.A(n_1290),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1304),
.B(n_826),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1315),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1315),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1324),
.B(n_1325),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1391),
.B(n_944),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1378),
.Y(n_1432)
);

AND2x6_ASAP7_75t_L g1433 ( 
.A(n_1334),
.B(n_1103),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1282),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1327),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1327),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1307),
.Y(n_1437)
);

INVx8_ASAP7_75t_L g1438 ( 
.A(n_1278),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1283),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1307),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1297),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1273),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1399),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1327),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1299),
.B(n_856),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1377),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1281),
.B(n_1029),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1285),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1339),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1281),
.B(n_1276),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1299),
.B(n_856),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1393),
.B(n_980),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1328),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1280),
.B(n_1291),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1393),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1322),
.B(n_964),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1406),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1272),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1334),
.B(n_1041),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1362),
.B(n_1122),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_SL g1461 ( 
.A(n_1314),
.B(n_843),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1381),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1274),
.A2(n_1131),
.B1(n_1125),
.B2(n_809),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1383),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1330),
.Y(n_1465)
);

AND2x6_ASAP7_75t_L g1466 ( 
.A(n_1330),
.B(n_1131),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1279),
.B(n_984),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1330),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1303),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1317),
.B(n_863),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1337),
.B(n_1002),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1272),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1284),
.B(n_989),
.Y(n_1473)
);

BUFx24_ASAP7_75t_SL g1474 ( 
.A(n_1298),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1339),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1360),
.B(n_995),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1339),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1389),
.B(n_1171),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1298),
.B(n_863),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1365),
.B(n_999),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1338),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1343),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1338),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1343),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1367),
.B(n_1013),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_R g1486 ( 
.A(n_1311),
.B(n_1179),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1369),
.B(n_1015),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1295),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1323),
.B(n_1019),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1371),
.B(n_1034),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1372),
.B(n_1044),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1389),
.B(n_1047),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1326),
.B(n_805),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1295),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1373),
.B(n_1065),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1346),
.B(n_1076),
.Y(n_1496)
);

CKINVDCx8_ASAP7_75t_R g1497 ( 
.A(n_1341),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1319),
.A2(n_852),
.B1(n_855),
.B2(n_843),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1374),
.B(n_1086),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1364),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1316),
.B(n_1376),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1364),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1380),
.B(n_1087),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1368),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1348),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1368),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1329),
.B(n_805),
.Y(n_1507)
);

CKINVDCx16_ASAP7_75t_R g1508 ( 
.A(n_1319),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1352),
.B(n_1116),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1370),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1388),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1316),
.B(n_863),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1354),
.B(n_1132),
.Y(n_1513)
);

AND2x2_ASAP7_75t_SL g1514 ( 
.A(n_1345),
.B(n_962),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1331),
.B(n_905),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1350),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1343),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1350),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1394),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1395),
.B(n_1157),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1287),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1366),
.Y(n_1522)
);

CKINVDCx6p67_ASAP7_75t_R g1523 ( 
.A(n_1351),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1398),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1400),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1332),
.B(n_905),
.Y(n_1526)
);

AND2x2_ASAP7_75t_SL g1527 ( 
.A(n_1344),
.B(n_846),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1405),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1370),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1301),
.B(n_874),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1292),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1384),
.B(n_803),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1301),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1293),
.Y(n_1534)
);

BUFx4f_ASAP7_75t_L g1535 ( 
.A(n_1351),
.Y(n_1535)
);

AND2x6_ASAP7_75t_L g1536 ( 
.A(n_1333),
.B(n_906),
.Y(n_1536)
);

AND2x6_ASAP7_75t_L g1537 ( 
.A(n_1320),
.B(n_906),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1336),
.B(n_806),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1340),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1294),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1313),
.B(n_1027),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1306),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1300),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1379),
.B(n_874),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1335),
.B(n_807),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1335),
.B(n_808),
.Y(n_1546)
);

BUFx8_ASAP7_75t_SL g1547 ( 
.A(n_1356),
.Y(n_1547)
);

CKINVDCx16_ASAP7_75t_R g1548 ( 
.A(n_1347),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1321),
.B(n_1308),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1386),
.B(n_1027),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1356),
.Y(n_1551)
);

AND2x4_ASAP7_75t_SL g1552 ( 
.A(n_1342),
.B(n_874),
.Y(n_1552)
);

BUFx10_ASAP7_75t_L g1553 ( 
.A(n_1403),
.Y(n_1553)
);

BUFx10_ASAP7_75t_L g1554 ( 
.A(n_1310),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1385),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1385),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1402),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1286),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1321),
.A2(n_1130),
.B1(n_1091),
.B2(n_1082),
.Y(n_1559)
);

INVx5_ASAP7_75t_L g1560 ( 
.A(n_1288),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1359),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1277),
.Y(n_1563)
);

AND2x6_ASAP7_75t_L g1564 ( 
.A(n_1289),
.B(n_1091),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_1349),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1277),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1353),
.Y(n_1567)
);

INVxp33_ASAP7_75t_L g1568 ( 
.A(n_1355),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1277),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1309),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1396),
.Y(n_1571)
);

AND2x6_ASAP7_75t_L g1572 ( 
.A(n_1404),
.B(n_1130),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1309),
.B(n_810),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1309),
.B(n_852),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1318),
.B(n_1056),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1363),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1363),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1363),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1407),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1387),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1387),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1387),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1397),
.Y(n_1583)
);

INVx5_ASAP7_75t_L g1584 ( 
.A(n_1397),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1305),
.B(n_970),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1302),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1305),
.B(n_1075),
.Y(n_1587)
);

INVx5_ASAP7_75t_L g1588 ( 
.A(n_1278),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1375),
.B(n_1153),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1375),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1375),
.B(n_849),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1305),
.B(n_1075),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1302),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1302),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1375),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1437),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1440),
.B(n_814),
.Y(n_1597)
);

NAND2x1p5_ASAP7_75t_L g1598 ( 
.A(n_1424),
.B(n_815),
.Y(n_1598)
);

AO22x2_ASAP7_75t_L g1599 ( 
.A1(n_1590),
.A2(n_1492),
.B1(n_1478),
.B2(n_1595),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1554),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1554),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1414),
.B(n_879),
.Y(n_1602)
);

BUFx8_ASAP7_75t_L g1603 ( 
.A(n_1446),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1462),
.B(n_923),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1605)
);

OAI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1474),
.A2(n_1411),
.B1(n_1496),
.B2(n_1458),
.C(n_1456),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1446),
.Y(n_1607)
);

AO22x1_ASAP7_75t_L g1608 ( 
.A1(n_1464),
.A2(n_881),
.B1(n_888),
.B2(n_879),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1450),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1540),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1479),
.A2(n_821),
.B1(n_824),
.B2(n_819),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1409),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1511),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1447),
.A2(n_1160),
.B1(n_1119),
.B2(n_829),
.C(n_830),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1508),
.A2(n_888),
.B1(n_892),
.B2(n_881),
.Y(n_1615)
);

AO22x2_ASAP7_75t_L g1616 ( 
.A1(n_1429),
.A2(n_897),
.B1(n_938),
.B2(n_892),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1519),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1524),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1454),
.B(n_1469),
.Y(n_1619)
);

NAND2x1p5_ASAP7_75t_L g1620 ( 
.A(n_1419),
.B(n_1174),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1525),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1504),
.B(n_1506),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1427),
.A2(n_833),
.B1(n_834),
.B2(n_828),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1528),
.Y(n_1624)
);

AO22x2_ASAP7_75t_L g1625 ( 
.A1(n_1429),
.A2(n_1460),
.B1(n_1498),
.B2(n_1589),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1545),
.B(n_839),
.C(n_837),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1457),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1488),
.Y(n_1628)
);

AO22x2_ASAP7_75t_L g1629 ( 
.A1(n_1589),
.A2(n_938),
.B1(n_940),
.B2(n_897),
.Y(n_1629)
);

NAND2x1p5_ASAP7_75t_L g1630 ( 
.A(n_1426),
.B(n_804),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1575),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1441),
.B(n_940),
.Y(n_1632)
);

AO22x2_ASAP7_75t_L g1633 ( 
.A1(n_1461),
.A2(n_985),
.B1(n_991),
.B2(n_983),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1488),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1443),
.B(n_983),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1574),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1494),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1448),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1481),
.A2(n_991),
.B1(n_996),
.B2(n_985),
.Y(n_1639)
);

BUFx8_ASAP7_75t_L g1640 ( 
.A(n_1567),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1521),
.Y(n_1641)
);

AO22x2_ASAP7_75t_L g1642 ( 
.A1(n_1586),
.A2(n_1594),
.B1(n_1593),
.B2(n_1423),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1531),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1472),
.B(n_1007),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1556),
.B(n_857),
.Y(n_1645)
);

AO22x2_ASAP7_75t_L g1646 ( 
.A1(n_1423),
.A2(n_1011),
.B1(n_1017),
.B2(n_1007),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1534),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1486),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1510),
.B(n_859),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1543),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1516),
.B(n_1011),
.Y(n_1651)
);

AO22x2_ASAP7_75t_L g1652 ( 
.A1(n_1574),
.A2(n_1038),
.B1(n_1054),
.B2(n_1033),
.Y(n_1652)
);

BUFx8_ASAP7_75t_L g1653 ( 
.A(n_1567),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1549),
.A2(n_817),
.B(n_818),
.C(n_811),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1457),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1575),
.Y(n_1656)
);

AO22x2_ASAP7_75t_L g1657 ( 
.A1(n_1410),
.A2(n_1067),
.B1(n_1093),
.B2(n_1054),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1509),
.A2(n_877),
.B1(n_883),
.B2(n_872),
.C(n_861),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1513),
.A2(n_887),
.B1(n_889),
.B2(n_886),
.C(n_885),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1445),
.B(n_1067),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1439),
.B(n_825),
.Y(n_1661)
);

AO22x2_ASAP7_75t_L g1662 ( 
.A1(n_1410),
.A2(n_1101),
.B1(n_1112),
.B2(n_1093),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1555),
.Y(n_1663)
);

AO22x2_ASAP7_75t_L g1664 ( 
.A1(n_1550),
.A2(n_1112),
.B1(n_1124),
.B2(n_1101),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1421),
.Y(n_1665)
);

AO22x2_ASAP7_75t_L g1666 ( 
.A1(n_1550),
.A2(n_1147),
.B1(n_1156),
.B2(n_1124),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1425),
.Y(n_1667)
);

AO22x2_ASAP7_75t_L g1668 ( 
.A1(n_1562),
.A2(n_1156),
.B1(n_1179),
.B2(n_1147),
.Y(n_1668)
);

AO22x2_ASAP7_75t_L g1669 ( 
.A1(n_1459),
.A2(n_831),
.B1(n_836),
.B2(n_827),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1522),
.Y(n_1670)
);

CKINVDCx14_ASAP7_75t_R g1671 ( 
.A(n_1518),
.Y(n_1671)
);

AO22x2_ASAP7_75t_L g1672 ( 
.A1(n_1459),
.A2(n_840),
.B1(n_841),
.B2(n_838),
.Y(n_1672)
);

CKINVDCx11_ASAP7_75t_R g1673 ( 
.A(n_1497),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1425),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1501),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1451),
.B(n_936),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1434),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1476),
.A2(n_925),
.B1(n_927),
.B2(n_920),
.C(n_913),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_1523),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1493),
.Y(n_1680)
);

AO22x2_ASAP7_75t_L g1681 ( 
.A1(n_1420),
.A2(n_854),
.B1(n_869),
.B2(n_860),
.Y(n_1681)
);

AO22x2_ASAP7_75t_L g1682 ( 
.A1(n_1432),
.A2(n_876),
.B1(n_880),
.B2(n_870),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1493),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1529),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1557),
.Y(n_1685)
);

AO22x2_ASAP7_75t_L g1686 ( 
.A1(n_1432),
.A2(n_890),
.B1(n_893),
.B2(n_884),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1412),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1471),
.B(n_894),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1435),
.Y(n_1689)
);

AO22x2_ASAP7_75t_L g1690 ( 
.A1(n_1507),
.A2(n_896),
.B1(n_899),
.B2(n_895),
.Y(n_1690)
);

OR2x6_ASAP7_75t_L g1691 ( 
.A(n_1471),
.B(n_846),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1585),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1415),
.B(n_982),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1587),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1592),
.Y(n_1695)
);

NAND2x1_ASAP7_75t_L g1696 ( 
.A(n_1466),
.B(n_849),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1455),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1413),
.B(n_931),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1490),
.A2(n_942),
.B1(n_943),
.B2(n_941),
.C(n_934),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1416),
.B(n_945),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1433),
.Y(n_1701)
);

NAND2x1p5_ASAP7_75t_L g1702 ( 
.A(n_1417),
.B(n_900),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1535),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1442),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1422),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1470),
.B(n_982),
.Y(n_1706)
);

AO22x2_ASAP7_75t_L g1707 ( 
.A1(n_1507),
.A2(n_904),
.B1(n_908),
.B2(n_902),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1467),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1473),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1560),
.B(n_950),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1512),
.B(n_982),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1421),
.Y(n_1712)
);

AO22x2_ASAP7_75t_L g1713 ( 
.A1(n_1515),
.A2(n_911),
.B1(n_914),
.B2(n_910),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1480),
.Y(n_1714)
);

AO22x2_ASAP7_75t_L g1715 ( 
.A1(n_1515),
.A2(n_1526),
.B1(n_1483),
.B2(n_1541),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1527),
.B(n_1129),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1485),
.Y(n_1717)
);

AO22x2_ASAP7_75t_L g1718 ( 
.A1(n_1526),
.A2(n_922),
.B1(n_924),
.B2(n_918),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1435),
.B(n_926),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1487),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1530),
.B(n_1129),
.Y(n_1721)
);

AO22x2_ASAP7_75t_L g1722 ( 
.A1(n_1541),
.A2(n_932),
.B1(n_937),
.B2(n_929),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1503),
.B(n_1129),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1533),
.B(n_948),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1491),
.Y(n_1725)
);

AND2x6_ASAP7_75t_L g1726 ( 
.A(n_1436),
.B(n_862),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1495),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1499),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1552),
.B(n_954),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1436),
.B(n_963),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1520),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1565),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1546),
.A2(n_1009),
.B1(n_1012),
.B2(n_1008),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1505),
.Y(n_1734)
);

AO22x2_ASAP7_75t_L g1735 ( 
.A1(n_1468),
.A2(n_971),
.B1(n_974),
.B2(n_965),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1547),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1553),
.B(n_1544),
.Y(n_1737)
);

AO22x2_ASAP7_75t_L g1738 ( 
.A1(n_1430),
.A2(n_976),
.B1(n_977),
.B2(n_975),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1532),
.A2(n_1022),
.B1(n_1023),
.B2(n_1018),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1539),
.B(n_979),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1538),
.A2(n_1042),
.B1(n_1045),
.B2(n_1040),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1489),
.B(n_981),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1452),
.A2(n_1052),
.B1(n_1055),
.B2(n_1050),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1542),
.A2(n_1060),
.B1(n_1061),
.B2(n_1057),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1548),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1568),
.A2(n_1068),
.B1(n_1069),
.B2(n_1064),
.C(n_1062),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_SL g1747 ( 
.A(n_1514),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1431),
.A2(n_1074),
.B1(n_1079),
.B2(n_1073),
.C(n_1071),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1428),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1551),
.B(n_987),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1571),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1542),
.B(n_1561),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1558),
.B(n_1083),
.Y(n_1753)
);

NAND2x1p5_ASAP7_75t_L g1754 ( 
.A(n_1444),
.B(n_990),
.Y(n_1754)
);

AO22x2_ASAP7_75t_L g1755 ( 
.A1(n_1517),
.A2(n_998),
.B1(n_1000),
.B2(n_997),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1466),
.Y(n_1756)
);

AO22x2_ASAP7_75t_L g1757 ( 
.A1(n_1482),
.A2(n_1004),
.B1(n_1006),
.B2(n_1001),
.Y(n_1757)
);

AO22x2_ASAP7_75t_L g1758 ( 
.A1(n_1591),
.A2(n_1014),
.B1(n_1024),
.B2(n_1010),
.Y(n_1758)
);

AO22x2_ASAP7_75t_L g1759 ( 
.A1(n_1408),
.A2(n_1035),
.B1(n_1043),
.B2(n_1026),
.Y(n_1759)
);

NAND2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1453),
.B(n_1046),
.Y(n_1760)
);

AO22x2_ASAP7_75t_L g1761 ( 
.A1(n_1438),
.A2(n_1059),
.B1(n_1063),
.B2(n_1051),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1465),
.B(n_1088),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1475),
.B(n_1089),
.Y(n_1763)
);

AO22x2_ASAP7_75t_L g1764 ( 
.A1(n_1438),
.A2(n_1072),
.B1(n_1078),
.B2(n_1066),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1463),
.A2(n_1094),
.B1(n_1096),
.B2(n_1090),
.Y(n_1765)
);

OAI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1559),
.A2(n_1099),
.B1(n_1102),
.B2(n_1098),
.C(n_1097),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1484),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1477),
.B(n_1080),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1573),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1418),
.B(n_1588),
.Y(n_1770)
);

AO22x2_ASAP7_75t_L g1771 ( 
.A1(n_1418),
.A2(n_1085),
.B1(n_1092),
.B2(n_1081),
.Y(n_1771)
);

AO22x2_ASAP7_75t_L g1772 ( 
.A1(n_1418),
.A2(n_1100),
.B1(n_1104),
.B2(n_1095),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1588),
.B(n_1105),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1537),
.A2(n_1111),
.B1(n_1115),
.B2(n_1109),
.Y(n_1774)
);

BUFx8_ASAP7_75t_L g1775 ( 
.A(n_1536),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1537),
.B(n_1120),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1588),
.B(n_1106),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1449),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1578),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1536),
.B(n_1108),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_SL g1781 ( 
.A(n_1564),
.Y(n_1781)
);

AO22x2_ASAP7_75t_L g1782 ( 
.A1(n_1582),
.A2(n_1114),
.B1(n_1121),
.B2(n_1110),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1572),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1576),
.B(n_1123),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1584),
.B(n_1128),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1572),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1572),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1584),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1584),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1563),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1580),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1580),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1581),
.A2(n_1138),
.B1(n_1141),
.B2(n_1137),
.C(n_1133),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1577),
.B(n_1142),
.Y(n_1794)
);

NAND2x1_ASAP7_75t_L g1795 ( 
.A(n_1583),
.B(n_849),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1579),
.A2(n_1145),
.B1(n_1146),
.B2(n_1144),
.C(n_1143),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1566),
.B(n_862),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1607),
.B(n_1186),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1600),
.B(n_1187),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1601),
.B(n_1148),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1605),
.B(n_1151),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1596),
.B(n_1622),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1598),
.B(n_1152),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1732),
.B(n_1154),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1684),
.B(n_1685),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1640),
.B(n_1169),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1653),
.B(n_1170),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1609),
.B(n_1172),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1603),
.B(n_1173),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1604),
.B(n_1630),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1627),
.B(n_1159),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1663),
.B(n_1162),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1767),
.B(n_1164),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1774),
.B(n_1184),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1628),
.B(n_1166),
.Y(n_1815)
);

NAND2xp33_ASAP7_75t_SL g1816 ( 
.A(n_1634),
.B(n_849),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1637),
.B(n_1180),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1687),
.B(n_1127),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1661),
.B(n_1566),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1708),
.B(n_1134),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1790),
.B(n_1569),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1632),
.B(n_1570),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1635),
.B(n_1570),
.Y(n_1823)
);

NAND2xp33_ASAP7_75t_SL g1824 ( 
.A(n_1756),
.B(n_912),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1709),
.B(n_1140),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1655),
.B(n_912),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1714),
.B(n_1150),
.Y(n_1827)
);

XNOR2xp5_ASAP7_75t_L g1828 ( 
.A(n_1633),
.B(n_4),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1717),
.B(n_1163),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1705),
.B(n_939),
.Y(n_1830)
);

NAND2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1638),
.B(n_939),
.Y(n_1831)
);

NAND2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1781),
.B(n_1641),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1779),
.B(n_1768),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1720),
.B(n_1168),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1702),
.B(n_1719),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1725),
.B(n_1175),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1727),
.B(n_1176),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1730),
.B(n_1754),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1760),
.B(n_1602),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1728),
.B(n_1181),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1734),
.B(n_939),
.Y(n_1841)
);

AND2x2_ASAP7_75t_SL g1842 ( 
.A(n_1636),
.B(n_988),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1679),
.B(n_1674),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1651),
.B(n_1036),
.Y(n_1844)
);

NAND2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1648),
.B(n_1036),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1731),
.B(n_1167),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1613),
.B(n_1185),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1675),
.B(n_882),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1737),
.B(n_973),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1608),
.B(n_1031),
.Y(n_1850)
);

NAND2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1786),
.B(n_1037),
.Y(n_1851)
);

NAND2xp33_ASAP7_75t_SL g1852 ( 
.A(n_1787),
.B(n_1053),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_SL g1853 ( 
.A(n_1787),
.B(n_1053),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1745),
.B(n_1135),
.Y(n_1854)
);

AND2x2_ASAP7_75t_SL g1855 ( 
.A(n_1639),
.B(n_4),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1617),
.B(n_5),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1762),
.B(n_7),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1763),
.B(n_1597),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1618),
.B(n_6),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1623),
.B(n_1752),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1716),
.B(n_8),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1644),
.B(n_9),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1785),
.B(n_9),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1706),
.B(n_10),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1744),
.B(n_10),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1740),
.B(n_10),
.Y(n_1866)
);

AND2x2_ASAP7_75t_SL g1867 ( 
.A(n_1782),
.B(n_8),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1711),
.B(n_11),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1621),
.B(n_8),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1729),
.B(n_12),
.Y(n_1870)
);

NAND2xp33_ASAP7_75t_SL g1871 ( 
.A(n_1703),
.B(n_11),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1606),
.B(n_12),
.Y(n_1872)
);

NAND2xp33_ASAP7_75t_SL g1873 ( 
.A(n_1667),
.B(n_12),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1676),
.B(n_16),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1784),
.B(n_16),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1721),
.B(n_16),
.Y(n_1876)
);

NAND2xp33_ASAP7_75t_SL g1877 ( 
.A(n_1610),
.B(n_14),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1765),
.B(n_18),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1688),
.B(n_19),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1733),
.B(n_19),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1753),
.B(n_19),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1669),
.B(n_17),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1750),
.B(n_21),
.Y(n_1883)
);

NAND2xp33_ASAP7_75t_SL g1884 ( 
.A(n_1747),
.B(n_20),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1624),
.B(n_20),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1620),
.B(n_23),
.Y(n_1886)
);

AND2x2_ASAP7_75t_SL g1887 ( 
.A(n_1782),
.B(n_22),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1701),
.B(n_1741),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1669),
.B(n_22),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1599),
.B(n_24),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1743),
.B(n_25),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1778),
.B(n_25),
.Y(n_1892)
);

NAND2xp33_ASAP7_75t_SL g1893 ( 
.A(n_1643),
.B(n_24),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1723),
.B(n_1612),
.Y(n_1894)
);

NAND2xp33_ASAP7_75t_SL g1895 ( 
.A(n_1647),
.B(n_24),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1611),
.B(n_27),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1599),
.B(n_26),
.Y(n_1897)
);

NAND2xp33_ASAP7_75t_SL g1898 ( 
.A(n_1650),
.B(n_26),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1739),
.B(n_30),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1654),
.B(n_29),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1776),
.B(n_32),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1660),
.B(n_33),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1775),
.B(n_33),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1680),
.B(n_31),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1665),
.B(n_31),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1689),
.B(n_35),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1626),
.B(n_1698),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1700),
.B(n_36),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1683),
.B(n_34),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1692),
.B(n_38),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1672),
.B(n_37),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_SL g1912 ( 
.A(n_1736),
.B(n_37),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1694),
.B(n_39),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1695),
.B(n_39),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1769),
.B(n_40),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1742),
.B(n_41),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1697),
.B(n_41),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1693),
.B(n_42),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1780),
.B(n_43),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1724),
.B(n_44),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1715),
.B(n_1722),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1722),
.B(n_41),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1658),
.B(n_45),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1682),
.B(n_45),
.Y(n_1924)
);

NAND2xp33_ASAP7_75t_SL g1925 ( 
.A(n_1712),
.B(n_46),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1773),
.B(n_47),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1777),
.B(n_47),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1751),
.B(n_47),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1682),
.B(n_46),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1686),
.B(n_48),
.Y(n_1930)
);

NAND2xp33_ASAP7_75t_SL g1931 ( 
.A(n_1615),
.B(n_48),
.Y(n_1931)
);

NAND2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1749),
.B(n_50),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1686),
.B(n_50),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1672),
.B(n_50),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1681),
.B(n_51),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1794),
.B(n_52),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1670),
.B(n_53),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1631),
.B(n_54),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1656),
.B(n_54),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1788),
.B(n_1645),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1681),
.B(n_56),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1649),
.B(n_57),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1677),
.B(n_56),
.Y(n_1943)
);

NAND2xp33_ASAP7_75t_SL g1944 ( 
.A(n_1789),
.B(n_59),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1704),
.B(n_59),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1710),
.B(n_62),
.Y(n_1946)
);

NAND2xp33_ASAP7_75t_SL g1947 ( 
.A(n_1696),
.B(n_59),
.Y(n_1947)
);

NAND2xp33_ASAP7_75t_SL g1948 ( 
.A(n_1791),
.B(n_63),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1792),
.B(n_64),
.Y(n_1949)
);

NAND2xp33_ASAP7_75t_SL g1950 ( 
.A(n_1642),
.B(n_63),
.Y(n_1950)
);

NAND2xp33_ASAP7_75t_SL g1951 ( 
.A(n_1642),
.B(n_65),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1770),
.B(n_67),
.Y(n_1952)
);

NAND2xp33_ASAP7_75t_SL g1953 ( 
.A(n_1783),
.B(n_65),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1757),
.B(n_69),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1797),
.B(n_69),
.Y(n_1955)
);

NAND2xp33_ASAP7_75t_SL g1956 ( 
.A(n_1625),
.B(n_1761),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1691),
.B(n_68),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1797),
.B(n_70),
.Y(n_1958)
);

NAND2xp33_ASAP7_75t_SL g1959 ( 
.A(n_1625),
.B(n_68),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1726),
.B(n_71),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_SL g1961 ( 
.A(n_1761),
.B(n_70),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1659),
.B(n_72),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1691),
.B(n_74),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1746),
.B(n_74),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1764),
.B(n_1771),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1690),
.B(n_73),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1764),
.B(n_74),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1690),
.B(n_73),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1707),
.B(n_73),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_SL g1970 ( 
.A(n_1772),
.B(n_75),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1707),
.B(n_77),
.Y(n_1971)
);

NAND2xp33_ASAP7_75t_SL g1972 ( 
.A(n_1652),
.B(n_76),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1713),
.B(n_79),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1718),
.B(n_79),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1718),
.B(n_79),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1738),
.B(n_78),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_SL g1977 ( 
.A(n_1652),
.B(n_78),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1795),
.B(n_78),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1657),
.B(n_82),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1657),
.B(n_82),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1616),
.B(n_1633),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1662),
.B(n_83),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1646),
.B(n_83),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1735),
.B(n_80),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1646),
.B(n_84),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_SL g1986 ( 
.A(n_1759),
.B(n_80),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1758),
.B(n_85),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1755),
.B(n_86),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_SL g1989 ( 
.A(n_1759),
.B(n_85),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1796),
.B(n_87),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1614),
.B(n_87),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1629),
.B(n_87),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1629),
.B(n_1793),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1616),
.B(n_86),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1664),
.B(n_88),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_SL g1996 ( 
.A(n_1664),
.B(n_86),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1666),
.B(n_89),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1666),
.B(n_89),
.Y(n_1998)
);

NAND2xp33_ASAP7_75t_SL g1999 ( 
.A(n_1668),
.B(n_88),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1748),
.B(n_90),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1673),
.B(n_90),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1668),
.B(n_90),
.Y(n_2002)
);

NAND2xp33_ASAP7_75t_SL g2003 ( 
.A(n_1678),
.B(n_1699),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1671),
.B(n_91),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1766),
.B(n_92),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1605),
.B(n_93),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1607),
.B(n_95),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1596),
.B(n_94),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1607),
.B(n_95),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1596),
.B(n_94),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_SL g2011 ( 
.A(n_1605),
.B(n_94),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1619),
.B(n_96),
.Y(n_2012)
);

NAND2xp33_ASAP7_75t_SL g2013 ( 
.A(n_1605),
.B(n_97),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1607),
.B(n_98),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1607),
.B(n_99),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1607),
.B(n_99),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1596),
.B(n_98),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1605),
.B(n_100),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1619),
.B(n_102),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1607),
.B(n_103),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1607),
.B(n_103),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1607),
.B(n_104),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1607),
.B(n_104),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1596),
.B(n_102),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1607),
.B(n_106),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1607),
.B(n_106),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1607),
.B(n_107),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1607),
.B(n_107),
.Y(n_2028)
);

NAND2xp33_ASAP7_75t_SL g2029 ( 
.A(n_1605),
.B(n_105),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1607),
.B(n_108),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_SL g2031 ( 
.A(n_1605),
.B(n_107),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1607),
.B(n_109),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1607),
.B(n_110),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1607),
.B(n_110),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1607),
.B(n_110),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1607),
.B(n_111),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1596),
.B(n_109),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1607),
.B(n_111),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1596),
.B(n_109),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1607),
.B(n_113),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1607),
.B(n_113),
.Y(n_2041)
);

NAND2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1605),
.B(n_112),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1607),
.B(n_115),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1600),
.B(n_114),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1607),
.B(n_115),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1607),
.B(n_116),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1607),
.B(n_117),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1607),
.B(n_119),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_SL g2049 ( 
.A(n_1605),
.B(n_118),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1607),
.B(n_118),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1607),
.B(n_120),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1600),
.B(n_119),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1607),
.B(n_120),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1607),
.B(n_120),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1607),
.B(n_122),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1596),
.B(n_121),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1607),
.B(n_123),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1619),
.B(n_122),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1607),
.B(n_125),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1607),
.B(n_126),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1607),
.B(n_126),
.Y(n_2061)
);

NAND2xp33_ASAP7_75t_SL g2062 ( 
.A(n_1605),
.B(n_126),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1607),
.B(n_128),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1607),
.B(n_128),
.Y(n_2064)
);

NAND2xp33_ASAP7_75t_SL g2065 ( 
.A(n_1605),
.B(n_127),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1619),
.B(n_127),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1607),
.B(n_129),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1596),
.B(n_128),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1607),
.B(n_130),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1619),
.B(n_132),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1607),
.B(n_135),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1607),
.B(n_135),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1607),
.B(n_135),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1607),
.B(n_137),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1607),
.B(n_137),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1607),
.B(n_138),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1607),
.B(n_138),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1607),
.B(n_138),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1619),
.B(n_136),
.Y(n_2079)
);

NAND2xp33_ASAP7_75t_SL g2080 ( 
.A(n_1605),
.B(n_136),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1619),
.B(n_140),
.Y(n_2081)
);

NAND2xp33_ASAP7_75t_SL g2082 ( 
.A(n_1605),
.B(n_140),
.Y(n_2082)
);

NAND2xp33_ASAP7_75t_SL g2083 ( 
.A(n_1605),
.B(n_141),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_SL g2084 ( 
.A(n_1605),
.B(n_141),
.Y(n_2084)
);

NAND2xp33_ASAP7_75t_SL g2085 ( 
.A(n_1605),
.B(n_142),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1607),
.B(n_143),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1607),
.B(n_143),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1607),
.B(n_143),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1607),
.B(n_144),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1607),
.B(n_144),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1607),
.B(n_145),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1607),
.B(n_146),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1619),
.B(n_145),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1607),
.B(n_148),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1600),
.B(n_147),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1607),
.B(n_149),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1607),
.B(n_149),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1607),
.B(n_149),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_1600),
.B(n_148),
.Y(n_2099)
);

NAND2xp33_ASAP7_75t_SL g2100 ( 
.A(n_1605),
.B(n_150),
.Y(n_2100)
);

NAND2xp33_ASAP7_75t_SL g2101 ( 
.A(n_1605),
.B(n_150),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1607),
.B(n_151),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1607),
.B(n_151),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1607),
.B(n_151),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1619),
.B(n_150),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1596),
.B(n_152),
.Y(n_2106)
);

NAND2xp33_ASAP7_75t_SL g2107 ( 
.A(n_1605),
.B(n_153),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1607),
.B(n_154),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1607),
.B(n_155),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1607),
.B(n_155),
.Y(n_2110)
);

NAND2xp33_ASAP7_75t_SL g2111 ( 
.A(n_1605),
.B(n_153),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1607),
.B(n_156),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1596),
.B(n_156),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1607),
.B(n_157),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1607),
.B(n_157),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1607),
.B(n_158),
.Y(n_2116)
);

AND2x2_ASAP7_75t_SL g2117 ( 
.A(n_1756),
.B(n_156),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1607),
.B(n_159),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1600),
.B(n_158),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1607),
.B(n_160),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1600),
.B(n_159),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1607),
.B(n_161),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1607),
.B(n_162),
.Y(n_2123)
);

NAND2xp33_ASAP7_75t_SL g2124 ( 
.A(n_1605),
.B(n_159),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1607),
.B(n_163),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1619),
.B(n_162),
.Y(n_2126)
);

NAND2xp33_ASAP7_75t_SL g2127 ( 
.A(n_1605),
.B(n_163),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1596),
.B(n_163),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1600),
.B(n_165),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1607),
.B(n_166),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1607),
.B(n_167),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1607),
.B(n_167),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1607),
.B(n_167),
.Y(n_2133)
);

NAND2xp33_ASAP7_75t_SL g2134 ( 
.A(n_1605),
.B(n_165),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1607),
.B(n_169),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1607),
.B(n_169),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1607),
.B(n_169),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_1860),
.B(n_168),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1945),
.Y(n_2139)
);

AOI21xp33_ASAP7_75t_L g2140 ( 
.A1(n_1872),
.A2(n_170),
.B(n_171),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1805),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1802),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1855),
.B(n_171),
.Y(n_2143)
);

INVx8_ASAP7_75t_L g2144 ( 
.A(n_1957),
.Y(n_2144)
);

OAI22x1_ASAP7_75t_L g2145 ( 
.A1(n_1828),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1882),
.B(n_1889),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2008),
.Y(n_2147)
);

AOI221xp5_ASAP7_75t_SL g2148 ( 
.A1(n_1965),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.C(n_178),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1816),
.A2(n_178),
.B(n_179),
.Y(n_2149)
);

AO21x2_ASAP7_75t_L g2150 ( 
.A1(n_1921),
.A2(n_1897),
.B(n_1890),
.Y(n_2150)
);

AOI21xp5_ASAP7_75t_L g2151 ( 
.A1(n_1816),
.A2(n_178),
.B(n_179),
.Y(n_2151)
);

AOI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_1831),
.A2(n_180),
.B(n_181),
.Y(n_2152)
);

AOI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_1831),
.A2(n_180),
.B(n_181),
.Y(n_2153)
);

CKINVDCx14_ASAP7_75t_R g2154 ( 
.A(n_1843),
.Y(n_2154)
);

OR2x6_ASAP7_75t_L g2155 ( 
.A(n_1957),
.B(n_182),
.Y(n_2155)
);

A2O1A1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_1956),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_1821),
.Y(n_2157)
);

NAND2x1p5_ASAP7_75t_L g2158 ( 
.A(n_1810),
.B(n_183),
.Y(n_2158)
);

AOI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_1907),
.A2(n_184),
.B(n_185),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_R g2160 ( 
.A(n_1832),
.B(n_185),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1855),
.B(n_186),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2012),
.B(n_186),
.Y(n_2162)
);

CKINVDCx11_ASAP7_75t_R g2163 ( 
.A(n_2001),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2019),
.B(n_187),
.Y(n_2164)
);

CKINVDCx11_ASAP7_75t_R g2165 ( 
.A(n_2001),
.Y(n_2165)
);

OA21x2_ASAP7_75t_L g2166 ( 
.A1(n_1987),
.A2(n_188),
.B(n_189),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2058),
.B(n_2066),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2003),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2168)
);

OAI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2010),
.A2(n_191),
.B(n_192),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1835),
.B(n_192),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_1957),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1869),
.Y(n_2172)
);

NAND2x1p5_ASAP7_75t_L g2173 ( 
.A(n_1842),
.B(n_193),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1858),
.A2(n_193),
.B(n_194),
.Y(n_2174)
);

NAND2x1p5_ASAP7_75t_L g2175 ( 
.A(n_1842),
.B(n_194),
.Y(n_2175)
);

INVx4_ASAP7_75t_L g2176 ( 
.A(n_1867),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1993),
.B(n_1981),
.Y(n_2177)
);

BUFx12f_ASAP7_75t_L g2178 ( 
.A(n_2001),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2070),
.B(n_195),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_1918),
.B(n_197),
.Y(n_2180)
);

BUFx10_ASAP7_75t_L g2181 ( 
.A(n_2004),
.Y(n_2181)
);

AO21x2_ASAP7_75t_L g2182 ( 
.A1(n_1954),
.A2(n_199),
.B(n_200),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1945),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2079),
.B(n_2081),
.Y(n_2184)
);

OAI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_1867),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2093),
.B(n_202),
.Y(n_2186)
);

BUFx4_ASAP7_75t_SL g2187 ( 
.A(n_1850),
.Y(n_2187)
);

OAI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_2017),
.A2(n_204),
.B(n_205),
.Y(n_2188)
);

NAND2x1p5_ASAP7_75t_L g2189 ( 
.A(n_1887),
.B(n_206),
.Y(n_2189)
);

BUFx5_ASAP7_75t_L g2190 ( 
.A(n_1945),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2105),
.B(n_206),
.Y(n_2191)
);

INVxp67_ASAP7_75t_SL g2192 ( 
.A(n_1869),
.Y(n_2192)
);

OAI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2024),
.A2(n_207),
.B(n_208),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2126),
.B(n_207),
.Y(n_2194)
);

NAND3xp33_ASAP7_75t_L g2195 ( 
.A(n_1959),
.B(n_208),
.C(n_209),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_2044),
.Y(n_2196)
);

INVx4_ASAP7_75t_L g2197 ( 
.A(n_1887),
.Y(n_2197)
);

OAI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_2037),
.A2(n_211),
.B(n_212),
.Y(n_2198)
);

INVx1_ASAP7_75t_SL g2199 ( 
.A(n_2044),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_L g2200 ( 
.A(n_1959),
.B(n_213),
.C(n_214),
.Y(n_2200)
);

NAND2xp33_ASAP7_75t_L g2201 ( 
.A(n_1830),
.B(n_793),
.Y(n_2201)
);

AO31x2_ASAP7_75t_L g2202 ( 
.A1(n_1976),
.A2(n_217),
.A3(n_215),
.B(n_216),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1885),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1885),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_2039),
.A2(n_218),
.B(n_219),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1820),
.B(n_219),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_SL g2207 ( 
.A(n_2117),
.B(n_1912),
.Y(n_2207)
);

BUFx5_ASAP7_75t_L g2208 ( 
.A(n_1885),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_SL g2209 ( 
.A(n_2117),
.B(n_220),
.Y(n_2209)
);

OAI22x1_ASAP7_75t_L g2210 ( 
.A1(n_1979),
.A2(n_222),
.B1(n_223),
.B2(n_221),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1820),
.B(n_224),
.Y(n_2211)
);

OAI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2056),
.A2(n_225),
.B(n_226),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1820),
.B(n_227),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1825),
.B(n_1827),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_2004),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2044),
.B(n_229),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_2004),
.Y(n_2217)
);

A2O1A1Ixp33_ASAP7_75t_L g2218 ( 
.A1(n_2006),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2068),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1825),
.B(n_233),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_2052),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1825),
.B(n_236),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2003),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_2223)
);

INVxp67_ASAP7_75t_L g2224 ( 
.A(n_2052),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1827),
.B(n_240),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1917),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1917),
.Y(n_2227)
);

NAND2x1p5_ASAP7_75t_L g2228 ( 
.A(n_1833),
.B(n_240),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1827),
.B(n_1847),
.Y(n_2229)
);

OA21x2_ASAP7_75t_L g2230 ( 
.A1(n_1935),
.A2(n_241),
.B(n_242),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1943),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1911),
.B(n_241),
.Y(n_2232)
);

OA22x2_ASAP7_75t_L g2233 ( 
.A1(n_1995),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_2233)
);

AOI221x1_ASAP7_75t_L g2234 ( 
.A1(n_1972),
.A2(n_1977),
.B1(n_1970),
.B2(n_1989),
.C(n_1986),
.Y(n_2234)
);

AND2x6_ASAP7_75t_L g2235 ( 
.A(n_1943),
.B(n_244),
.Y(n_2235)
);

NAND3xp33_ASAP7_75t_L g2236 ( 
.A(n_1972),
.B(n_245),
.C(n_246),
.Y(n_2236)
);

OAI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_2106),
.A2(n_245),
.B(n_246),
.Y(n_2237)
);

AOI21xp5_ASAP7_75t_SL g2238 ( 
.A1(n_2052),
.A2(n_247),
.B(n_248),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2113),
.Y(n_2239)
);

OA21x2_ASAP7_75t_L g2240 ( 
.A1(n_1941),
.A2(n_249),
.B(n_250),
.Y(n_2240)
);

NAND3x1_ASAP7_75t_L g2241 ( 
.A(n_1994),
.B(n_1934),
.C(n_1966),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2128),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1856),
.Y(n_2243)
);

A2O1A1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_2006),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2244)
);

AO32x2_ASAP7_75t_L g2245 ( 
.A1(n_1950),
.A2(n_1951),
.A3(n_1986),
.B1(n_1989),
.B2(n_1977),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1859),
.Y(n_2246)
);

NAND2x1p5_ASAP7_75t_L g2247 ( 
.A(n_2095),
.B(n_256),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2005),
.A2(n_257),
.B(n_258),
.Y(n_2248)
);

AO31x2_ASAP7_75t_L g2249 ( 
.A1(n_1924),
.A2(n_261),
.A3(n_259),
.B(n_260),
.Y(n_2249)
);

NOR4xp25_ASAP7_75t_L g2250 ( 
.A(n_1980),
.B(n_264),
.C(n_262),
.D(n_263),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1847),
.B(n_262),
.Y(n_2251)
);

INVx1_ASAP7_75t_SL g2252 ( 
.A(n_2095),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1902),
.B(n_264),
.Y(n_2253)
);

OAI22xp5_ASAP7_75t_L g2254 ( 
.A1(n_2095),
.A2(n_268),
.B1(n_265),
.B2(n_266),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1948),
.Y(n_2255)
);

AO31x2_ASAP7_75t_L g2256 ( 
.A1(n_1929),
.A2(n_269),
.A3(n_266),
.B(n_268),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1904),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1829),
.B(n_269),
.Y(n_2258)
);

INVx5_ASAP7_75t_L g2259 ( 
.A(n_2099),
.Y(n_2259)
);

INVx2_ASAP7_75t_SL g2260 ( 
.A(n_2099),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_1824),
.B(n_270),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1834),
.B(n_1836),
.Y(n_2262)
);

NAND2x1p5_ASAP7_75t_L g2263 ( 
.A(n_2099),
.B(n_272),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2119),
.B(n_272),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1837),
.B(n_273),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1840),
.B(n_274),
.Y(n_2266)
);

OAI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_1990),
.A2(n_274),
.B(n_275),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1846),
.B(n_275),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1923),
.B(n_276),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1978),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1978),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1962),
.B(n_277),
.Y(n_2272)
);

BUFx2_ASAP7_75t_L g2273 ( 
.A(n_2119),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2119),
.B(n_278),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1894),
.B(n_280),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1909),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1818),
.B(n_282),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1922),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2050),
.B(n_282),
.Y(n_2279)
);

BUFx2_ASAP7_75t_L g2280 ( 
.A(n_2121),
.Y(n_2280)
);

NOR4xp25_ASAP7_75t_L g2281 ( 
.A(n_1982),
.B(n_285),
.C(n_283),
.D(n_284),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1864),
.B(n_1862),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_1888),
.A2(n_283),
.B(n_284),
.Y(n_2283)
);

AND2x2_ASAP7_75t_SL g2284 ( 
.A(n_2121),
.B(n_2129),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1968),
.Y(n_2285)
);

CKINVDCx8_ASAP7_75t_R g2286 ( 
.A(n_2121),
.Y(n_2286)
);

OAI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_1908),
.A2(n_289),
.B(n_290),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1969),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2129),
.B(n_1997),
.Y(n_2289)
);

AO31x2_ASAP7_75t_L g2290 ( 
.A1(n_1930),
.A2(n_1933),
.A3(n_1900),
.B(n_1984),
.Y(n_2290)
);

AOI221x1_ASAP7_75t_L g2291 ( 
.A1(n_1970),
.A2(n_1961),
.B1(n_2002),
.B2(n_1999),
.C(n_1996),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1868),
.B(n_289),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2129),
.B(n_290),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1874),
.B(n_291),
.Y(n_2294)
);

AO32x2_ASAP7_75t_L g2295 ( 
.A1(n_1950),
.A2(n_294),
.A3(n_291),
.B1(n_292),
.B2(n_295),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_1876),
.B(n_297),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1978),
.Y(n_2297)
);

OAI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_1964),
.A2(n_300),
.B(n_301),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_1910),
.A2(n_1914),
.B(n_1913),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1896),
.B(n_302),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_1967),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_1861),
.Y(n_2302)
);

NOR4xp25_ASAP7_75t_L g2303 ( 
.A(n_1992),
.B(n_1998),
.C(n_1985),
.D(n_1983),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1949),
.Y(n_2304)
);

INVx3_ASAP7_75t_SL g2305 ( 
.A(n_1806),
.Y(n_2305)
);

A2O1A1Ixp33_ASAP7_75t_L g2306 ( 
.A1(n_2011),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1893),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1916),
.B(n_307),
.Y(n_2308)
);

BUFx3_ASAP7_75t_L g2309 ( 
.A(n_1848),
.Y(n_2309)
);

A2O1A1Ixp33_ASAP7_75t_L g2310 ( 
.A1(n_2011),
.A2(n_311),
.B(n_308),
.C(n_310),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_1971),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1893),
.Y(n_2312)
);

AO32x2_ASAP7_75t_L g2313 ( 
.A1(n_1951),
.A2(n_315),
.A3(n_313),
.B1(n_314),
.B2(n_316),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1839),
.B(n_318),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_1891),
.B(n_321),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_1940),
.A2(n_321),
.B(n_322),
.Y(n_2316)
);

NOR2xp67_ASAP7_75t_L g2317 ( 
.A(n_1803),
.B(n_323),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1895),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_1973),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2080),
.A2(n_331),
.B(n_332),
.Y(n_2320)
);

INVxp67_ASAP7_75t_L g2321 ( 
.A(n_1996),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1899),
.B(n_333),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_1819),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_1974),
.B(n_337),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1928),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_1878),
.A2(n_338),
.B(n_339),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_1975),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2327)
);

BUFx3_ASAP7_75t_L g2328 ( 
.A(n_1812),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1857),
.B(n_1875),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_L g2330 ( 
.A(n_2002),
.B(n_341),
.C(n_342),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1988),
.Y(n_2331)
);

BUFx5_ASAP7_75t_L g2332 ( 
.A(n_2080),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_1841),
.A2(n_344),
.B(n_345),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1938),
.Y(n_2334)
);

AOI221x1_ASAP7_75t_L g2335 ( 
.A1(n_1961),
.A2(n_347),
.B1(n_344),
.B2(n_346),
.C(n_348),
.Y(n_2335)
);

BUFx4f_ASAP7_75t_L g2336 ( 
.A(n_1832),
.Y(n_2336)
);

OAI21xp33_ASAP7_75t_L g2337 ( 
.A1(n_1991),
.A2(n_352),
.B(n_353),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_1838),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1880),
.B(n_355),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1865),
.B(n_358),
.Y(n_2340)
);

AO31x2_ASAP7_75t_L g2341 ( 
.A1(n_2082),
.A2(n_360),
.A3(n_358),
.B(n_359),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2083),
.A2(n_359),
.B(n_360),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1939),
.Y(n_2343)
);

AO32x2_ASAP7_75t_L g2344 ( 
.A1(n_1898),
.A2(n_363),
.A3(n_361),
.B1(n_362),
.B2(n_364),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_1854),
.B(n_365),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_1807),
.B(n_365),
.Y(n_2346)
);

A2O1A1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_2083),
.A2(n_369),
.B(n_366),
.C(n_368),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2084),
.A2(n_370),
.B(n_371),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_1798),
.B(n_1822),
.Y(n_2349)
);

A2O1A1Ixp33_ASAP7_75t_L g2350 ( 
.A1(n_2085),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2000),
.B(n_1863),
.Y(n_2351)
);

OAI22x1_ASAP7_75t_L g2352 ( 
.A1(n_1903),
.A2(n_378),
.B1(n_375),
.B2(n_376),
.Y(n_2352)
);

AO31x2_ASAP7_75t_L g2353 ( 
.A1(n_2100),
.A2(n_380),
.A3(n_378),
.B(n_379),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_1870),
.B(n_380),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_1955),
.Y(n_2355)
);

AO32x2_ASAP7_75t_L g2356 ( 
.A1(n_1898),
.A2(n_383),
.A3(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_2356)
);

NAND2x1p5_ASAP7_75t_L g2357 ( 
.A(n_1809),
.B(n_381),
.Y(n_2357)
);

OAI22x1_ASAP7_75t_L g2358 ( 
.A1(n_1963),
.A2(n_386),
.B1(n_383),
.B2(n_385),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_1884),
.Y(n_2359)
);

AO31x2_ASAP7_75t_L g2360 ( 
.A1(n_2100),
.A2(n_390),
.A3(n_388),
.B(n_389),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1915),
.Y(n_2361)
);

AOI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2101),
.A2(n_392),
.B(n_393),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_1823),
.B(n_394),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_1883),
.B(n_395),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_1801),
.B(n_396),
.Y(n_2365)
);

NAND3xp33_ASAP7_75t_SL g2366 ( 
.A(n_1931),
.B(n_397),
.C(n_398),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_1942),
.B(n_399),
.Y(n_2367)
);

OAI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_1958),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_2368)
);

INVx1_ASAP7_75t_SL g2369 ( 
.A(n_1826),
.Y(n_2369)
);

NOR2x1_ASAP7_75t_SL g2370 ( 
.A(n_1960),
.B(n_404),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2007),
.B(n_405),
.Y(n_2371)
);

BUFx2_ASAP7_75t_L g2372 ( 
.A(n_2101),
.Y(n_2372)
);

AND2x4_ASAP7_75t_L g2373 ( 
.A(n_1946),
.B(n_407),
.Y(n_2373)
);

OR2x2_ASAP7_75t_L g2374 ( 
.A(n_1866),
.B(n_409),
.Y(n_2374)
);

OAI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2009),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_2375)
);

OAI21xp5_ASAP7_75t_SL g2376 ( 
.A1(n_1886),
.A2(n_412),
.B(n_413),
.Y(n_2376)
);

OAI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_1936),
.A2(n_412),
.B(n_413),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_1813),
.Y(n_2378)
);

OAI21xp33_ASAP7_75t_L g2379 ( 
.A1(n_1881),
.A2(n_414),
.B(n_415),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_1873),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2107),
.A2(n_416),
.B(n_417),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_1814),
.B(n_418),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_SL g2383 ( 
.A(n_2111),
.B(n_418),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1937),
.Y(n_2384)
);

AOI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2124),
.A2(n_420),
.B(n_421),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2127),
.B(n_420),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_SL g2387 ( 
.A1(n_1952),
.A2(n_421),
.B(n_422),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_1849),
.B(n_422),
.Y(n_2388)
);

OA21x2_ASAP7_75t_L g2389 ( 
.A1(n_1901),
.A2(n_423),
.B(n_424),
.Y(n_2389)
);

AO31x2_ASAP7_75t_L g2390 ( 
.A1(n_2134),
.A2(n_427),
.A3(n_425),
.B(n_426),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_1879),
.B(n_427),
.Y(n_2391)
);

INVx6_ASAP7_75t_L g2392 ( 
.A(n_1871),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_1844),
.B(n_428),
.Y(n_2393)
);

A2O1A1Ixp33_ASAP7_75t_L g2394 ( 
.A1(n_2013),
.A2(n_433),
.B(n_431),
.C(n_432),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_1845),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2014),
.B(n_2015),
.Y(n_2396)
);

AOI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2018),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2029),
.A2(n_438),
.B(n_440),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_1815),
.B(n_441),
.Y(n_2399)
);

OA21x2_ASAP7_75t_L g2400 ( 
.A1(n_1906),
.A2(n_442),
.B(n_443),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2016),
.B(n_444),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_1905),
.Y(n_2402)
);

NAND3xp33_ASAP7_75t_L g2403 ( 
.A(n_1947),
.B(n_445),
.C(n_446),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2020),
.B(n_447),
.Y(n_2404)
);

INVx4_ASAP7_75t_L g2405 ( 
.A(n_1944),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2021),
.B(n_448),
.Y(n_2406)
);

OAI21xp33_ASAP7_75t_L g2407 ( 
.A1(n_2022),
.A2(n_449),
.B(n_450),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_1920),
.B(n_450),
.Y(n_2408)
);

BUFx2_ASAP7_75t_L g2409 ( 
.A(n_2031),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2137),
.Y(n_2410)
);

BUFx10_ASAP7_75t_L g2411 ( 
.A(n_2042),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2023),
.B(n_2025),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2026),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2136),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_1905),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2027),
.B(n_2028),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2135),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2030),
.B(n_2032),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2049),
.A2(n_458),
.B(n_459),
.Y(n_2419)
);

INVx5_ASAP7_75t_L g2420 ( 
.A(n_1947),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2033),
.Y(n_2421)
);

AOI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2062),
.A2(n_459),
.B(n_460),
.Y(n_2422)
);

BUFx2_ASAP7_75t_L g2423 ( 
.A(n_2065),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_SL g2424 ( 
.A1(n_2034),
.A2(n_461),
.B(n_463),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2035),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2036),
.B(n_461),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1925),
.Y(n_2427)
);

NOR2xp67_ASAP7_75t_SL g2428 ( 
.A(n_2038),
.B(n_463),
.Y(n_2428)
);

NAND2x1p5_ASAP7_75t_L g2429 ( 
.A(n_1919),
.B(n_464),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2040),
.B(n_466),
.Y(n_2430)
);

CKINVDCx20_ASAP7_75t_R g2431 ( 
.A(n_1811),
.Y(n_2431)
);

NAND3xp33_ASAP7_75t_L g2432 ( 
.A(n_1925),
.B(n_466),
.C(n_467),
.Y(n_2432)
);

AOI221xp5_ASAP7_75t_L g2433 ( 
.A1(n_1877),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.C(n_471),
.Y(n_2433)
);

AO31x2_ASAP7_75t_L g2434 ( 
.A1(n_1953),
.A2(n_472),
.A3(n_470),
.B(n_471),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_1817),
.A2(n_472),
.B(n_473),
.Y(n_2435)
);

OAI22x1_ASAP7_75t_L g2436 ( 
.A1(n_2041),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2133),
.Y(n_2437)
);

INVxp67_ASAP7_75t_SL g2438 ( 
.A(n_2043),
.Y(n_2438)
);

NAND2xp33_ASAP7_75t_SL g2439 ( 
.A(n_2045),
.B(n_477),
.Y(n_2439)
);

OAI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_2046),
.A2(n_478),
.B(n_479),
.Y(n_2440)
);

AOI21xp33_ASAP7_75t_L g2441 ( 
.A1(n_1808),
.A2(n_478),
.B(n_479),
.Y(n_2441)
);

BUFx3_ASAP7_75t_L g2442 ( 
.A(n_1932),
.Y(n_2442)
);

NAND3xp33_ASAP7_75t_L g2443 ( 
.A(n_1932),
.B(n_481),
.C(n_483),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2132),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2047),
.B(n_484),
.Y(n_2445)
);

A2O1A1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2048),
.A2(n_2053),
.B(n_2054),
.C(n_2051),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2131),
.Y(n_2447)
);

INVx5_ASAP7_75t_L g2448 ( 
.A(n_1852),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2055),
.A2(n_485),
.B(n_486),
.Y(n_2449)
);

NOR2x1_ASAP7_75t_L g2450 ( 
.A(n_2057),
.B(n_487),
.Y(n_2450)
);

OAI21x1_ASAP7_75t_L g2451 ( 
.A1(n_2059),
.A2(n_489),
.B(n_490),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2201),
.A2(n_2061),
.B(n_2060),
.Y(n_2452)
);

O2A1O1Ixp33_ASAP7_75t_L g2453 ( 
.A1(n_2446),
.A2(n_1892),
.B(n_2064),
.C(n_2063),
.Y(n_2453)
);

OA21x2_ASAP7_75t_L g2454 ( 
.A1(n_2234),
.A2(n_2069),
.B(n_2067),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2142),
.Y(n_2455)
);

AOI222xp33_ASAP7_75t_SL g2456 ( 
.A1(n_2185),
.A2(n_493),
.B1(n_495),
.B2(n_491),
.C1(n_492),
.C2(n_494),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2141),
.B(n_2146),
.Y(n_2457)
);

AOI22xp33_ASAP7_75t_SL g2458 ( 
.A1(n_2207),
.A2(n_2072),
.B1(n_2073),
.B2(n_2071),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2259),
.B(n_1926),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2290),
.B(n_2074),
.Y(n_2460)
);

O2A1O1Ixp33_ASAP7_75t_L g2461 ( 
.A1(n_2262),
.A2(n_2075),
.B(n_2077),
.C(n_2076),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2215),
.B(n_1804),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2290),
.B(n_2078),
.Y(n_2463)
);

INVx1_ASAP7_75t_SL g2464 ( 
.A(n_2284),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2216),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2216),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2176),
.A2(n_2087),
.B1(n_2088),
.B2(n_2086),
.Y(n_2467)
);

OAI21x1_ASAP7_75t_L g2468 ( 
.A1(n_2427),
.A2(n_2090),
.B(n_2089),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2290),
.B(n_2091),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2163),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2178),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2264),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2155),
.B(n_2092),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2187),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2165),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_2176),
.A2(n_2096),
.B1(n_2097),
.B2(n_2094),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_SL g2477 ( 
.A(n_2405),
.B(n_1851),
.Y(n_2477)
);

OA21x2_ASAP7_75t_L g2478 ( 
.A1(n_2291),
.A2(n_2102),
.B(n_2098),
.Y(n_2478)
);

HB1xp67_ASAP7_75t_L g2479 ( 
.A(n_2155),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2144),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2232),
.B(n_2103),
.Y(n_2481)
);

OA21x2_ASAP7_75t_L g2482 ( 
.A1(n_2307),
.A2(n_2108),
.B(n_2104),
.Y(n_2482)
);

BUFx3_ASAP7_75t_L g2483 ( 
.A(n_2144),
.Y(n_2483)
);

HB1xp67_ASAP7_75t_L g2484 ( 
.A(n_2286),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2274),
.B(n_2293),
.Y(n_2485)
);

AOI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_2197),
.A2(n_2110),
.B1(n_2112),
.B2(n_2109),
.Y(n_2486)
);

NAND2x1p5_ASAP7_75t_L g2487 ( 
.A(n_2259),
.B(n_1927),
.Y(n_2487)
);

OR2x6_ASAP7_75t_L g2488 ( 
.A(n_2247),
.B(n_2114),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2259),
.B(n_2115),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2209),
.B(n_1853),
.Y(n_2490)
);

O2A1O1Ixp33_ASAP7_75t_L g2491 ( 
.A1(n_2269),
.A2(n_2118),
.B(n_2120),
.C(n_2116),
.Y(n_2491)
);

OA21x2_ASAP7_75t_L g2492 ( 
.A1(n_2312),
.A2(n_2123),
.B(n_2122),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2264),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_2154),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2217),
.Y(n_2495)
);

INVx2_ASAP7_75t_SL g2496 ( 
.A(n_2336),
.Y(n_2496)
);

OR2x6_ASAP7_75t_L g2497 ( 
.A(n_2263),
.B(n_2125),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2278),
.B(n_2130),
.Y(n_2498)
);

AO31x2_ASAP7_75t_L g2499 ( 
.A1(n_2255),
.A2(n_496),
.A3(n_491),
.B(n_492),
.Y(n_2499)
);

OAI21x1_ASAP7_75t_L g2500 ( 
.A1(n_2318),
.A2(n_1800),
.B(n_1799),
.Y(n_2500)
);

OR2x6_ASAP7_75t_L g2501 ( 
.A(n_2405),
.B(n_499),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2197),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2285),
.B(n_502),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2288),
.B(n_503),
.Y(n_2504)
);

AOI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_2192),
.A2(n_503),
.B(n_504),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2336),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2160),
.Y(n_2507)
);

O2A1O1Ixp33_ASAP7_75t_L g2508 ( 
.A1(n_2272),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_2305),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2261),
.A2(n_505),
.B(n_506),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2249),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2208),
.Y(n_2512)
);

OAI221xp5_ASAP7_75t_L g2513 ( 
.A1(n_2189),
.A2(n_802),
.B1(n_511),
.B2(n_509),
.C(n_510),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2167),
.B(n_512),
.Y(n_2514)
);

CKINVDCx16_ASAP7_75t_R g2515 ( 
.A(n_2346),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2147),
.B(n_514),
.Y(n_2516)
);

NAND2x1p5_ASAP7_75t_L g2517 ( 
.A(n_2171),
.B(n_801),
.Y(n_2517)
);

OR2x2_ASAP7_75t_L g2518 ( 
.A(n_2184),
.B(n_515),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2235),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2420),
.B(n_516),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2177),
.A2(n_520),
.B1(n_517),
.B2(n_519),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2249),
.Y(n_2522)
);

HB1xp67_ASAP7_75t_L g2523 ( 
.A(n_2170),
.Y(n_2523)
);

CKINVDCx20_ASAP7_75t_R g2524 ( 
.A(n_2431),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2256),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2147),
.B(n_2219),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2256),
.Y(n_2527)
);

HB1xp67_ASAP7_75t_L g2528 ( 
.A(n_2170),
.Y(n_2528)
);

A2O1A1Ixp33_ASAP7_75t_L g2529 ( 
.A1(n_2383),
.A2(n_523),
.B(n_521),
.C(n_522),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2219),
.B(n_522),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2208),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2145),
.B(n_524),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2256),
.Y(n_2533)
);

AND2x4_ASAP7_75t_L g2534 ( 
.A(n_2420),
.B(n_2139),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2208),
.Y(n_2535)
);

NAND2x1p5_ASAP7_75t_L g2536 ( 
.A(n_2420),
.B(n_526),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2208),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2328),
.B(n_527),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_2139),
.B(n_528),
.Y(n_2539)
);

BUFx4f_ASAP7_75t_SL g2540 ( 
.A(n_2181),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2181),
.Y(n_2541)
);

NAND2x1p5_ASAP7_75t_L g2542 ( 
.A(n_2204),
.B(n_800),
.Y(n_2542)
);

OAI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2173),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2214),
.B(n_529),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2202),
.Y(n_2545)
);

HB1xp67_ASAP7_75t_L g2546 ( 
.A(n_2309),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2202),
.Y(n_2547)
);

O2A1O1Ixp5_ASAP7_75t_L g2548 ( 
.A1(n_2386),
.A2(n_533),
.B(n_530),
.C(n_532),
.Y(n_2548)
);

OAI21xp5_ASAP7_75t_L g2549 ( 
.A1(n_2248),
.A2(n_534),
.B(n_535),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2196),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2202),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2229),
.B(n_539),
.Y(n_2552)
);

NAND3x1_ASAP7_75t_L g2553 ( 
.A(n_2330),
.B(n_541),
.C(n_542),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2239),
.B(n_543),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2204),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2372),
.A2(n_547),
.B(n_549),
.Y(n_2556)
);

O2A1O1Ixp33_ASAP7_75t_SL g2557 ( 
.A1(n_2218),
.A2(n_552),
.B(n_550),
.C(n_551),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2341),
.Y(n_2558)
);

OAI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2175),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_2559)
);

INVxp67_ASAP7_75t_L g2560 ( 
.A(n_2235),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2221),
.B(n_555),
.Y(n_2561)
);

AO21x2_ASAP7_75t_L g2562 ( 
.A1(n_2303),
.A2(n_800),
.B(n_556),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2199),
.A2(n_558),
.B(n_559),
.Y(n_2563)
);

AO31x2_ASAP7_75t_L g2564 ( 
.A1(n_2335),
.A2(n_562),
.A3(n_560),
.B(n_561),
.Y(n_2564)
);

OAI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2273),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_2565)
);

INVx3_ASAP7_75t_SL g2566 ( 
.A(n_2346),
.Y(n_2566)
);

AOI21xp33_ASAP7_75t_L g2567 ( 
.A1(n_2321),
.A2(n_565),
.B(n_566),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2162),
.B(n_566),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2231),
.Y(n_2569)
);

AOI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2235),
.A2(n_570),
.B1(n_567),
.B2(n_568),
.Y(n_2570)
);

AOI22xp33_ASAP7_75t_SL g2571 ( 
.A1(n_2235),
.A2(n_575),
.B1(n_571),
.B2(n_574),
.Y(n_2571)
);

NAND2x1_ASAP7_75t_L g2572 ( 
.A(n_2183),
.B(n_574),
.Y(n_2572)
);

CKINVDCx20_ASAP7_75t_R g2573 ( 
.A(n_2378),
.Y(n_2573)
);

OAI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2280),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2190),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2138),
.A2(n_580),
.B1(n_577),
.B2(n_578),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2302),
.B(n_580),
.Y(n_2577)
);

INVx1_ASAP7_75t_SL g2578 ( 
.A(n_2252),
.Y(n_2578)
);

OAI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2169),
.A2(n_581),
.B(n_582),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2359),
.B(n_581),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2260),
.A2(n_585),
.B(n_586),
.Y(n_2581)
);

BUFx3_ASAP7_75t_L g2582 ( 
.A(n_2231),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2354),
.B(n_585),
.Y(n_2583)
);

INVx5_ASAP7_75t_L g2584 ( 
.A(n_2231),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_L g2585 ( 
.A(n_2355),
.B(n_588),
.Y(n_2585)
);

OAI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2270),
.A2(n_2297),
.B(n_2271),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2364),
.B(n_589),
.Y(n_2587)
);

NAND2x1p5_ASAP7_75t_L g2588 ( 
.A(n_2183),
.B(n_589),
.Y(n_2588)
);

NAND2x1p5_ASAP7_75t_L g2589 ( 
.A(n_2183),
.B(n_799),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2166),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2341),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2157),
.Y(n_2592)
);

BUFx2_ASAP7_75t_R g2593 ( 
.A(n_2143),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2203),
.A2(n_590),
.B(n_591),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2166),
.Y(n_2595)
);

CKINVDCx11_ASAP7_75t_R g2596 ( 
.A(n_2411),
.Y(n_2596)
);

BUFx2_ASAP7_75t_SL g2597 ( 
.A(n_2317),
.Y(n_2597)
);

AOI21x1_ASAP7_75t_L g2598 ( 
.A1(n_2409),
.A2(n_591),
.B(n_592),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_2402),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2226),
.A2(n_593),
.B(n_594),
.Y(n_2600)
);

AO21x2_ASAP7_75t_L g2601 ( 
.A1(n_2195),
.A2(n_595),
.B(n_596),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2239),
.B(n_596),
.Y(n_2602)
);

BUFx3_ASAP7_75t_L g2603 ( 
.A(n_2357),
.Y(n_2603)
);

AOI21xp33_ASAP7_75t_L g2604 ( 
.A1(n_2331),
.A2(n_597),
.B(n_598),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2353),
.Y(n_2605)
);

NAND2x1p5_ASAP7_75t_L g2606 ( 
.A(n_2395),
.B(n_597),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2242),
.Y(n_2607)
);

CKINVDCx20_ASAP7_75t_R g2608 ( 
.A(n_2392),
.Y(n_2608)
);

OA21x2_ASAP7_75t_L g2609 ( 
.A1(n_2148),
.A2(n_600),
.B(n_601),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2242),
.Y(n_2610)
);

BUFx4_ASAP7_75t_SL g2611 ( 
.A(n_2415),
.Y(n_2611)
);

AO21x2_ASAP7_75t_L g2612 ( 
.A1(n_2200),
.A2(n_798),
.B(n_600),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_SL g2613 ( 
.A1(n_2380),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2164),
.B(n_604),
.Y(n_2614)
);

BUFx6f_ASAP7_75t_L g2615 ( 
.A(n_2338),
.Y(n_2615)
);

OR2x6_ASAP7_75t_SL g2616 ( 
.A(n_2254),
.B(n_606),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2243),
.B(n_606),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_2352),
.Y(n_2618)
);

BUFx2_ASAP7_75t_L g2619 ( 
.A(n_2392),
.Y(n_2619)
);

INVx5_ASAP7_75t_L g2620 ( 
.A(n_2411),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2238),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2423),
.A2(n_2289),
.B1(n_2366),
.B2(n_2439),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2353),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2243),
.B(n_607),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2353),
.Y(n_2625)
);

CKINVDCx11_ASAP7_75t_R g2626 ( 
.A(n_2369),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2360),
.Y(n_2627)
);

INVx3_ASAP7_75t_L g2628 ( 
.A(n_2442),
.Y(n_2628)
);

NAND2x1p5_ASAP7_75t_L g2629 ( 
.A(n_2428),
.B(n_609),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2360),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2360),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2390),
.Y(n_2632)
);

INVx1_ASAP7_75t_SL g2633 ( 
.A(n_2332),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2390),
.Y(n_2634)
);

AOI21xp5_ASAP7_75t_L g2635 ( 
.A1(n_2152),
.A2(n_609),
.B(n_611),
.Y(n_2635)
);

OAI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2298),
.A2(n_611),
.B(n_612),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2246),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2246),
.B(n_612),
.Y(n_2638)
);

CKINVDCx20_ASAP7_75t_R g2639 ( 
.A(n_2224),
.Y(n_2639)
);

NAND2x1p5_ASAP7_75t_L g2640 ( 
.A(n_2448),
.B(n_797),
.Y(n_2640)
);

OR2x6_ASAP7_75t_L g2641 ( 
.A(n_2153),
.B(n_613),
.Y(n_2641)
);

BUFx10_ASAP7_75t_L g2642 ( 
.A(n_2367),
.Y(n_2642)
);

INVx2_ASAP7_75t_SL g2643 ( 
.A(n_2158),
.Y(n_2643)
);

NAND2x1p5_ASAP7_75t_L g2644 ( 
.A(n_2448),
.B(n_616),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2179),
.B(n_2186),
.Y(n_2645)
);

AOI221xp5_ASAP7_75t_L g2646 ( 
.A1(n_2140),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.C(n_622),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2391),
.B(n_621),
.Y(n_2647)
);

NAND2xp33_ASAP7_75t_SL g2648 ( 
.A(n_2161),
.B(n_624),
.Y(n_2648)
);

BUFx12f_ASAP7_75t_L g2649 ( 
.A(n_2228),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2180),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_2650)
);

BUFx8_ASAP7_75t_SL g2651 ( 
.A(n_2367),
.Y(n_2651)
);

AO31x2_ASAP7_75t_L g2652 ( 
.A1(n_2156),
.A2(n_628),
.A3(n_625),
.B(n_626),
.Y(n_2652)
);

OAI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2267),
.A2(n_629),
.B(n_632),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2206),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2324),
.B(n_629),
.Y(n_2655)
);

AND2x4_ASAP7_75t_L g2656 ( 
.A(n_2172),
.B(n_633),
.Y(n_2656)
);

OAI221xp5_ASAP7_75t_L g2657 ( 
.A1(n_2168),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.C(n_637),
.Y(n_2657)
);

BUFx2_ASAP7_75t_L g2658 ( 
.A(n_2332),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2374),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2408),
.Y(n_2660)
);

BUFx3_ASAP7_75t_L g2661 ( 
.A(n_2338),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2338),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2257),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2276),
.Y(n_2664)
);

OR2x2_ASAP7_75t_L g2665 ( 
.A(n_2211),
.B(n_638),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2213),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2233),
.Y(n_2667)
);

INVx3_ASAP7_75t_L g2668 ( 
.A(n_2332),
.Y(n_2668)
);

AO21x2_ASAP7_75t_L g2669 ( 
.A1(n_2150),
.A2(n_797),
.B(n_639),
.Y(n_2669)
);

NAND2x1p5_ASAP7_75t_L g2670 ( 
.A(n_2448),
.B(n_2227),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2332),
.B(n_641),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_2361),
.B(n_643),
.Y(n_2672)
);

CKINVDCx20_ASAP7_75t_R g2673 ( 
.A(n_2349),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2351),
.A2(n_643),
.B(n_644),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2332),
.B(n_645),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2418),
.B(n_647),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2373),
.A2(n_648),
.B1(n_649),
.B2(n_650),
.Y(n_2677)
);

OAI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2174),
.A2(n_651),
.B(n_652),
.Y(n_2678)
);

BUFx3_ASAP7_75t_L g2679 ( 
.A(n_2323),
.Y(n_2679)
);

AO21x2_ASAP7_75t_L g2680 ( 
.A1(n_2188),
.A2(n_651),
.B(n_652),
.Y(n_2680)
);

OAI21xp5_ASAP7_75t_SL g2681 ( 
.A1(n_2376),
.A2(n_655),
.B(n_656),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2323),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2304),
.B(n_655),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2434),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2373),
.A2(n_657),
.B1(n_658),
.B2(n_659),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2345),
.B(n_659),
.Y(n_2686)
);

OAI21xp5_ASAP7_75t_L g2687 ( 
.A1(n_2326),
.A2(n_660),
.B(n_661),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2191),
.B(n_660),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2325),
.B(n_2334),
.Y(n_2689)
);

INVx1_ASAP7_75t_SL g2690 ( 
.A(n_2323),
.Y(n_2690)
);

A2O1A1Ixp33_ASAP7_75t_SL g2691 ( 
.A1(n_2393),
.A2(n_2382),
.B(n_2365),
.C(n_2193),
.Y(n_2691)
);

OA21x2_ASAP7_75t_L g2692 ( 
.A1(n_2337),
.A2(n_662),
.B(n_663),
.Y(n_2692)
);

HB1xp67_ASAP7_75t_L g2693 ( 
.A(n_2220),
.Y(n_2693)
);

CKINVDCx11_ASAP7_75t_R g2694 ( 
.A(n_2410),
.Y(n_2694)
);

BUFx2_ASAP7_75t_L g2695 ( 
.A(n_2241),
.Y(n_2695)
);

BUFx6f_ASAP7_75t_L g2696 ( 
.A(n_2333),
.Y(n_2696)
);

AOI21xp33_ASAP7_75t_SL g2697 ( 
.A1(n_2358),
.A2(n_665),
.B(n_666),
.Y(n_2697)
);

OAI21x1_ASAP7_75t_SL g2698 ( 
.A1(n_2370),
.A2(n_666),
.B(n_667),
.Y(n_2698)
);

BUFx2_ASAP7_75t_L g2699 ( 
.A(n_2429),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2436),
.Y(n_2700)
);

OA21x2_ASAP7_75t_L g2701 ( 
.A1(n_2198),
.A2(n_671),
.B(n_672),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2434),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2314),
.Y(n_2703)
);

OA21x2_ASAP7_75t_L g2704 ( 
.A1(n_2205),
.A2(n_672),
.B(n_673),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2343),
.B(n_675),
.Y(n_2705)
);

OR2x6_ASAP7_75t_L g2706 ( 
.A(n_2149),
.B(n_675),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2245),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_R g2708 ( 
.A1(n_2311),
.A2(n_676),
.B(n_677),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2182),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2449),
.Y(n_2710)
);

OR2x6_ASAP7_75t_L g2711 ( 
.A(n_2151),
.B(n_678),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_2275),
.Y(n_2712)
);

BUFx2_ASAP7_75t_L g2713 ( 
.A(n_2245),
.Y(n_2713)
);

OAI21x1_ASAP7_75t_SL g2714 ( 
.A1(n_2320),
.A2(n_679),
.B(n_680),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2222),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2194),
.B(n_681),
.Y(n_2716)
);

BUFx10_ASAP7_75t_L g2717 ( 
.A(n_2363),
.Y(n_2717)
);

BUFx12f_ASAP7_75t_L g2718 ( 
.A(n_2387),
.Y(n_2718)
);

OAI211xp5_ASAP7_75t_L g2719 ( 
.A1(n_2433),
.A2(n_681),
.B(n_682),
.C(n_683),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2225),
.B(n_684),
.Y(n_2720)
);

OA21x2_ASAP7_75t_L g2721 ( 
.A1(n_2212),
.A2(n_684),
.B(n_685),
.Y(n_2721)
);

OAI22xp5_ASAP7_75t_L g2722 ( 
.A1(n_2236),
.A2(n_687),
.B1(n_689),
.B2(n_690),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2244),
.A2(n_692),
.B1(n_693),
.B2(n_695),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2384),
.B(n_2299),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2451),
.Y(n_2725)
);

NAND3x1_ASAP7_75t_L g2726 ( 
.A(n_2450),
.B(n_692),
.C(n_693),
.Y(n_2726)
);

CKINVDCx6p67_ASAP7_75t_R g2727 ( 
.A(n_2210),
.Y(n_2727)
);

OAI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2159),
.A2(n_696),
.B(n_697),
.Y(n_2728)
);

OA21x2_ASAP7_75t_L g2729 ( 
.A1(n_2237),
.A2(n_698),
.B(n_700),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2251),
.Y(n_2730)
);

O2A1O1Ixp33_ASAP7_75t_L g2731 ( 
.A1(n_2329),
.A2(n_701),
.B(n_702),
.C(n_703),
.Y(n_2731)
);

AO31x2_ASAP7_75t_L g2732 ( 
.A1(n_2306),
.A2(n_701),
.A3(n_702),
.B(n_704),
.Y(n_2732)
);

CKINVDCx20_ASAP7_75t_R g2733 ( 
.A(n_2397),
.Y(n_2733)
);

AO31x2_ASAP7_75t_L g2734 ( 
.A1(n_2310),
.A2(n_705),
.A3(n_706),
.B(n_707),
.Y(n_2734)
);

OAI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2347),
.A2(n_705),
.B1(n_706),
.B2(n_707),
.Y(n_2735)
);

INVx6_ASAP7_75t_L g2736 ( 
.A(n_2424),
.Y(n_2736)
);

AND2x6_ASAP7_75t_L g2737 ( 
.A(n_2223),
.B(n_796),
.Y(n_2737)
);

OR2x6_ASAP7_75t_L g2738 ( 
.A(n_2342),
.B(n_709),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2308),
.Y(n_2739)
);

BUFx3_ASAP7_75t_L g2740 ( 
.A(n_2400),
.Y(n_2740)
);

OAI221xp5_ASAP7_75t_L g2741 ( 
.A1(n_2282),
.A2(n_794),
.B1(n_711),
.B2(n_712),
.C(n_713),
.Y(n_2741)
);

OAI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2350),
.A2(n_710),
.B1(n_711),
.B2(n_712),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2344),
.Y(n_2743)
);

NOR2xp67_ASAP7_75t_L g2744 ( 
.A(n_2403),
.B(n_710),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2344),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2230),
.Y(n_2746)
);

AOI221xp5_ASAP7_75t_L g2747 ( 
.A1(n_2250),
.A2(n_713),
.B1(n_714),
.B2(n_716),
.C(n_717),
.Y(n_2747)
);

AO21x2_ASAP7_75t_L g2748 ( 
.A1(n_2348),
.A2(n_716),
.B(n_718),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2240),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_2546),
.Y(n_2750)
);

INVx1_ASAP7_75t_SL g2751 ( 
.A(n_2599),
.Y(n_2751)
);

BUFx2_ASAP7_75t_L g2752 ( 
.A(n_2480),
.Y(n_2752)
);

CKINVDCx20_ASAP7_75t_R g2753 ( 
.A(n_2524),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2663),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_SL g2755 ( 
.A1(n_2501),
.A2(n_2394),
.B(n_2240),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2457),
.B(n_2344),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2607),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2664),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2610),
.Y(n_2759)
);

INVx5_ASAP7_75t_L g2760 ( 
.A(n_2501),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2534),
.Y(n_2761)
);

BUFx6f_ASAP7_75t_L g2762 ( 
.A(n_2483),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2455),
.Y(n_2763)
);

HB1xp67_ASAP7_75t_L g2764 ( 
.A(n_2658),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2474),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2637),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2526),
.Y(n_2767)
);

INVx3_ASAP7_75t_L g2768 ( 
.A(n_2534),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2516),
.Y(n_2769)
);

OR2x2_ASAP7_75t_L g2770 ( 
.A(n_2485),
.B(n_2281),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2516),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2530),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2727),
.A2(n_2414),
.B1(n_2421),
.B2(n_2417),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2530),
.Y(n_2774)
);

INVxp67_ASAP7_75t_L g2775 ( 
.A(n_2695),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2554),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2554),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2602),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2645),
.B(n_2532),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_SL g2780 ( 
.A1(n_2515),
.A2(n_2443),
.B1(n_2432),
.B2(n_2301),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2602),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_2670),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2617),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2501),
.A2(n_2362),
.B1(n_2385),
.B2(n_2381),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2617),
.Y(n_2785)
);

OR2x2_ASAP7_75t_L g2786 ( 
.A(n_2479),
.B(n_2258),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2624),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2624),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_2633),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2676),
.B(n_2356),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_L g2791 ( 
.A1(n_2737),
.A2(n_2425),
.B1(n_2444),
.B2(n_2437),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2670),
.Y(n_2792)
);

INVx3_ASAP7_75t_L g2793 ( 
.A(n_2620),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2638),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2620),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2560),
.B(n_2447),
.Y(n_2796)
);

BUFx3_ASAP7_75t_L g2797 ( 
.A(n_2471),
.Y(n_2797)
);

OR2x2_ASAP7_75t_L g2798 ( 
.A(n_2514),
.B(n_2265),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2460),
.B(n_2438),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2638),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2659),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2660),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_L g2803 ( 
.A(n_2733),
.B(n_2616),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_2651),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2583),
.B(n_2356),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2503),
.Y(n_2806)
);

INVx1_ASAP7_75t_SL g2807 ( 
.A(n_2599),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2503),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2587),
.B(n_2356),
.Y(n_2809)
);

INVxp33_ASAP7_75t_L g2810 ( 
.A(n_2626),
.Y(n_2810)
);

OR2x2_ASAP7_75t_L g2811 ( 
.A(n_2518),
.B(n_2266),
.Y(n_2811)
);

BUFx2_ASAP7_75t_L g2812 ( 
.A(n_2608),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_2596),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2647),
.B(n_2295),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2504),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2504),
.Y(n_2816)
);

HB1xp67_ASAP7_75t_L g2817 ( 
.A(n_2633),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2689),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2689),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2705),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2519),
.A2(n_2398),
.B1(n_2419),
.B2(n_2422),
.Y(n_2821)
);

BUFx2_ASAP7_75t_L g2822 ( 
.A(n_2495),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2705),
.Y(n_2823)
);

OR2x6_ASAP7_75t_L g2824 ( 
.A(n_2536),
.B(n_2283),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2460),
.B(n_2315),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2667),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2499),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2620),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_2573),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2655),
.B(n_2295),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2737),
.A2(n_2566),
.B1(n_2513),
.B2(n_2657),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2499),
.Y(n_2832)
);

O2A1O1Ixp33_ASAP7_75t_L g2833 ( 
.A1(n_2691),
.A2(n_2279),
.B(n_2416),
.C(n_2396),
.Y(n_2833)
);

INVx2_ASAP7_75t_SL g2834 ( 
.A(n_2611),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2481),
.B(n_2295),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2561),
.B(n_2313),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2584),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2499),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2538),
.B(n_2313),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2683),
.Y(n_2840)
);

INVx1_ASAP7_75t_SL g2841 ( 
.A(n_2628),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2584),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2470),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2688),
.B(n_2313),
.Y(n_2844)
);

BUFx2_ASAP7_75t_SL g2845 ( 
.A(n_2475),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2509),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2584),
.Y(n_2847)
);

AND2x4_ASAP7_75t_L g2848 ( 
.A(n_2520),
.B(n_2316),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2656),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2656),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2590),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2595),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2716),
.B(n_719),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2477),
.B(n_2440),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2746),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2749),
.Y(n_2856)
);

BUFx2_ASAP7_75t_SL g2857 ( 
.A(n_2496),
.Y(n_2857)
);

BUFx6f_ASAP7_75t_L g2858 ( 
.A(n_2582),
.Y(n_2858)
);

INVx1_ASAP7_75t_SL g2859 ( 
.A(n_2628),
.Y(n_2859)
);

BUFx6f_ASAP7_75t_L g2860 ( 
.A(n_2615),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2672),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2672),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2724),
.Y(n_2863)
);

INVx3_ASAP7_75t_SL g2864 ( 
.A(n_2507),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2463),
.B(n_2322),
.Y(n_2865)
);

AND2x4_ASAP7_75t_L g2866 ( 
.A(n_2520),
.B(n_2287),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2493),
.B(n_720),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2539),
.Y(n_2868)
);

BUFx3_ASAP7_75t_L g2869 ( 
.A(n_2540),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2724),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2539),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2465),
.Y(n_2872)
);

HB1xp67_ASAP7_75t_L g2873 ( 
.A(n_2668),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2466),
.Y(n_2874)
);

AOI22xp33_ASAP7_75t_L g2875 ( 
.A1(n_2737),
.A2(n_2407),
.B1(n_2327),
.B2(n_2319),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2472),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2739),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2671),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_L g2879 ( 
.A1(n_2737),
.A2(n_2379),
.B1(n_2377),
.B2(n_2388),
.Y(n_2879)
);

NOR2x1_ASAP7_75t_R g2880 ( 
.A(n_2494),
.B(n_2412),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2473),
.B(n_720),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2519),
.A2(n_2400),
.B1(n_2268),
.B2(n_2277),
.Y(n_2882)
);

AO22x1_ASAP7_75t_L g2883 ( 
.A1(n_2700),
.A2(n_2368),
.B1(n_2375),
.B2(n_2413),
.Y(n_2883)
);

BUFx3_ASAP7_75t_L g2884 ( 
.A(n_2592),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2671),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2619),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2464),
.B(n_2253),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2598),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2720),
.B(n_721),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2642),
.Y(n_2890)
);

BUFx6f_ASAP7_75t_L g2891 ( 
.A(n_2615),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2523),
.B(n_721),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2558),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2528),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2591),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2464),
.A2(n_2389),
.B1(n_2300),
.B2(n_2340),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2605),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2649),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2623),
.Y(n_2899)
);

INVx4_ASAP7_75t_L g2900 ( 
.A(n_2642),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2625),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2627),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2630),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2631),
.Y(n_2904)
);

HB1xp67_ASAP7_75t_L g2905 ( 
.A(n_2463),
.Y(n_2905)
);

INVx3_ASAP7_75t_L g2906 ( 
.A(n_2506),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2632),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2634),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_2694),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2498),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2654),
.B(n_722),
.Y(n_2911)
);

HB1xp67_ASAP7_75t_L g2912 ( 
.A(n_2469),
.Y(n_2912)
);

BUFx2_ASAP7_75t_L g2913 ( 
.A(n_2661),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_2603),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2666),
.B(n_722),
.Y(n_2915)
);

BUFx2_ASAP7_75t_L g2916 ( 
.A(n_2484),
.Y(n_2916)
);

INVx3_ASAP7_75t_L g2917 ( 
.A(n_2736),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2498),
.Y(n_2918)
);

CKINVDCx6p67_ASAP7_75t_R g2919 ( 
.A(n_2597),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2732),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2693),
.B(n_723),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2469),
.B(n_2339),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2541),
.Y(n_2923)
);

INVx6_ASAP7_75t_L g2924 ( 
.A(n_2718),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2732),
.Y(n_2925)
);

OAI21x1_ASAP7_75t_SL g2926 ( 
.A1(n_2681),
.A2(n_2435),
.B(n_2445),
.Y(n_2926)
);

BUFx3_ASAP7_75t_L g2927 ( 
.A(n_2673),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2732),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2734),
.Y(n_2929)
);

INVx3_ASAP7_75t_L g2930 ( 
.A(n_2736),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2734),
.Y(n_2931)
);

INVx2_ASAP7_75t_SL g2932 ( 
.A(n_2606),
.Y(n_2932)
);

BUFx2_ASAP7_75t_L g2933 ( 
.A(n_2679),
.Y(n_2933)
);

AOI22xp33_ASAP7_75t_L g2934 ( 
.A1(n_2513),
.A2(n_2292),
.B1(n_2294),
.B2(n_2296),
.Y(n_2934)
);

OR2x6_ASAP7_75t_L g2935 ( 
.A(n_2640),
.B(n_2245),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2712),
.B(n_723),
.Y(n_2936)
);

BUFx2_ASAP7_75t_L g2937 ( 
.A(n_2682),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2730),
.B(n_2743),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2585),
.B(n_724),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2709),
.Y(n_2940)
);

BUFx2_ASAP7_75t_L g2941 ( 
.A(n_2639),
.Y(n_2941)
);

INVx4_ASAP7_75t_L g2942 ( 
.A(n_2644),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2684),
.Y(n_2943)
);

AND2x4_ASAP7_75t_L g2944 ( 
.A(n_2555),
.B(n_2371),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_SL g2945 ( 
.A1(n_2618),
.A2(n_2399),
.B1(n_2430),
.B2(n_2426),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_SL g2946 ( 
.A1(n_2613),
.A2(n_2406),
.B1(n_2404),
.B2(n_2401),
.Y(n_2946)
);

INVx2_ASAP7_75t_SL g2947 ( 
.A(n_2699),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2702),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2652),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2745),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2652),
.Y(n_2951)
);

AND2x4_ASAP7_75t_L g2952 ( 
.A(n_2569),
.B(n_724),
.Y(n_2952)
);

BUFx2_ASAP7_75t_L g2953 ( 
.A(n_2662),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2517),
.Y(n_2954)
);

AO21x1_ASAP7_75t_SL g2955 ( 
.A1(n_2622),
.A2(n_2441),
.B(n_726),
.Y(n_2955)
);

BUFx3_ASAP7_75t_L g2956 ( 
.A(n_2569),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2568),
.B(n_792),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2652),
.Y(n_2958)
);

INVx1_ASAP7_75t_SL g2959 ( 
.A(n_2550),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2703),
.Y(n_2960)
);

INVx2_ASAP7_75t_SL g2961 ( 
.A(n_2488),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2511),
.B(n_725),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2614),
.B(n_727),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2657),
.A2(n_727),
.B1(n_728),
.B2(n_730),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2565),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2522),
.B(n_731),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2512),
.B(n_2531),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2565),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2574),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2715),
.B(n_2650),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2650),
.B(n_792),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2574),
.Y(n_2972)
);

INVx3_ASAP7_75t_L g2973 ( 
.A(n_2662),
.Y(n_2973)
);

OAI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2681),
.A2(n_731),
.B1(n_732),
.B2(n_733),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2748),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2488),
.Y(n_2976)
);

AO21x2_ASAP7_75t_L g2977 ( 
.A1(n_2710),
.A2(n_733),
.B(n_734),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2748),
.Y(n_2978)
);

AO21x2_ASAP7_75t_L g2979 ( 
.A1(n_2725),
.A2(n_734),
.B(n_735),
.Y(n_2979)
);

INVx3_ASAP7_75t_L g2980 ( 
.A(n_2542),
.Y(n_2980)
);

BUFx2_ASAP7_75t_SL g2981 ( 
.A(n_2643),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2669),
.Y(n_2982)
);

OAI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2708),
.A2(n_735),
.B1(n_736),
.B2(n_737),
.Y(n_2983)
);

INVx3_ASAP7_75t_L g2984 ( 
.A(n_2588),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2747),
.A2(n_2741),
.B1(n_2648),
.B2(n_2735),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2577),
.B(n_2576),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2459),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2576),
.B(n_791),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2544),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2571),
.B(n_791),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2552),
.Y(n_2991)
);

BUFx3_ASAP7_75t_L g2992 ( 
.A(n_2535),
.Y(n_2992)
);

OAI211xp5_ASAP7_75t_L g2993 ( 
.A1(n_2697),
.A2(n_738),
.B(n_740),
.C(n_741),
.Y(n_2993)
);

CKINVDCx20_ASAP7_75t_R g2994 ( 
.A(n_2621),
.Y(n_2994)
);

INVx3_ASAP7_75t_L g2995 ( 
.A(n_2589),
.Y(n_2995)
);

INVx3_ASAP7_75t_L g2996 ( 
.A(n_2537),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2564),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2525),
.B(n_743),
.Y(n_2998)
);

CKINVDCx12_ASAP7_75t_R g2999 ( 
.A(n_2613),
.Y(n_2999)
);

INVxp67_ASAP7_75t_L g3000 ( 
.A(n_2750),
.Y(n_3000)
);

INVxp67_ASAP7_75t_L g3001 ( 
.A(n_2752),
.Y(n_3001)
);

INVxp67_ASAP7_75t_L g3002 ( 
.A(n_2822),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_R g3003 ( 
.A(n_2898),
.B(n_2580),
.Y(n_3003)
);

XNOR2xp5_ASAP7_75t_L g3004 ( 
.A(n_2813),
.B(n_2804),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2760),
.B(n_2697),
.Y(n_3005)
);

NAND2xp33_ASAP7_75t_R g3006 ( 
.A(n_2804),
.B(n_2488),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2779),
.B(n_2550),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_R g3008 ( 
.A(n_2898),
.B(n_2462),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2801),
.Y(n_3009)
);

NAND2xp33_ASAP7_75t_R g3010 ( 
.A(n_2909),
.B(n_2497),
.Y(n_3010)
);

INVxp67_ASAP7_75t_L g3011 ( 
.A(n_2880),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_R g3012 ( 
.A(n_2753),
.B(n_2717),
.Y(n_3012)
);

XNOR2xp5_ASAP7_75t_L g3013 ( 
.A(n_2813),
.B(n_2726),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_R g3014 ( 
.A(n_2753),
.B(n_2717),
.Y(n_3014)
);

XNOR2xp5_ASAP7_75t_L g3015 ( 
.A(n_2843),
.B(n_2559),
.Y(n_3015)
);

NAND2xp33_ASAP7_75t_R g3016 ( 
.A(n_2909),
.B(n_2497),
.Y(n_3016)
);

OR2x4_ASAP7_75t_L g3017 ( 
.A(n_2803),
.B(n_2686),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_2762),
.Y(n_3018)
);

BUFx12f_ASAP7_75t_L g3019 ( 
.A(n_2834),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2802),
.B(n_2578),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_R g3021 ( 
.A(n_2994),
.B(n_744),
.Y(n_3021)
);

NAND2xp33_ASAP7_75t_R g3022 ( 
.A(n_2803),
.B(n_2497),
.Y(n_3022)
);

AND2x4_ASAP7_75t_L g3023 ( 
.A(n_2760),
.B(n_2578),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2881),
.B(n_2707),
.Y(n_3024)
);

INVxp67_ASAP7_75t_L g3025 ( 
.A(n_2880),
.Y(n_3025)
);

NAND2xp33_ASAP7_75t_R g3026 ( 
.A(n_2793),
.B(n_2701),
.Y(n_3026)
);

INVxp67_ASAP7_75t_L g3027 ( 
.A(n_2981),
.Y(n_3027)
);

NAND2xp33_ASAP7_75t_R g3028 ( 
.A(n_2793),
.B(n_2701),
.Y(n_3028)
);

NAND2xp33_ASAP7_75t_R g3029 ( 
.A(n_2795),
.B(n_2704),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2959),
.B(n_2713),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2959),
.B(n_2690),
.Y(n_3031)
);

NAND2xp33_ASAP7_75t_R g3032 ( 
.A(n_2795),
.B(n_2704),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2754),
.B(n_2747),
.Y(n_3033)
);

BUFx3_ASAP7_75t_L g3034 ( 
.A(n_2797),
.Y(n_3034)
);

AND2x4_ASAP7_75t_L g3035 ( 
.A(n_2761),
.B(n_2575),
.Y(n_3035)
);

CKINVDCx12_ASAP7_75t_R g3036 ( 
.A(n_2935),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_2758),
.B(n_2690),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_2900),
.B(n_2556),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2877),
.B(n_2527),
.Y(n_3039)
);

NOR2xp33_ASAP7_75t_R g3040 ( 
.A(n_2994),
.B(n_744),
.Y(n_3040)
);

XNOR2xp5_ASAP7_75t_L g3041 ( 
.A(n_2810),
.B(n_2559),
.Y(n_3041)
);

BUFx6f_ASAP7_75t_L g3042 ( 
.A(n_2762),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2960),
.B(n_2533),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_R g3044 ( 
.A(n_2869),
.B(n_2919),
.Y(n_3044)
);

NAND2xp33_ASAP7_75t_R g3045 ( 
.A(n_2828),
.B(n_2721),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_R g3046 ( 
.A(n_2762),
.B(n_745),
.Y(n_3046)
);

NAND2xp33_ASAP7_75t_R g3047 ( 
.A(n_2828),
.B(n_2721),
.Y(n_3047)
);

AND2x4_ASAP7_75t_L g3048 ( 
.A(n_2935),
.B(n_2545),
.Y(n_3048)
);

AND2x4_ASAP7_75t_L g3049 ( 
.A(n_2935),
.B(n_2547),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2900),
.B(n_2556),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_R g3051 ( 
.A(n_2864),
.B(n_745),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2894),
.B(n_2562),
.Y(n_3052)
);

AND2x4_ASAP7_75t_L g3053 ( 
.A(n_2768),
.B(n_2913),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2927),
.B(n_2593),
.Y(n_3054)
);

BUFx3_ASAP7_75t_L g3055 ( 
.A(n_2884),
.Y(n_3055)
);

NAND2xp33_ASAP7_75t_R g3056 ( 
.A(n_2812),
.B(n_2729),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2763),
.Y(n_3057)
);

OR2x6_ASAP7_75t_L g3058 ( 
.A(n_2924),
.B(n_2857),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2766),
.Y(n_3059)
);

XNOR2xp5_ASAP7_75t_L g3060 ( 
.A(n_2810),
.B(n_2553),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2970),
.B(n_2562),
.Y(n_3061)
);

NAND2xp33_ASAP7_75t_R g3062 ( 
.A(n_2941),
.B(n_2729),
.Y(n_3062)
);

AND2x4_ASAP7_75t_L g3063 ( 
.A(n_2764),
.B(n_2863),
.Y(n_3063)
);

AND2x4_ASAP7_75t_L g3064 ( 
.A(n_2764),
.B(n_2551),
.Y(n_3064)
);

NAND2xp33_ASAP7_75t_R g3065 ( 
.A(n_2890),
.B(n_2692),
.Y(n_3065)
);

AND2x4_ASAP7_75t_L g3066 ( 
.A(n_2870),
.B(n_2740),
.Y(n_3066)
);

NAND2xp33_ASAP7_75t_R g3067 ( 
.A(n_2890),
.B(n_2692),
.Y(n_3067)
);

NAND2xp33_ASAP7_75t_R g3068 ( 
.A(n_2837),
.B(n_2842),
.Y(n_3068)
);

NAND2xp33_ASAP7_75t_R g3069 ( 
.A(n_2837),
.B(n_2609),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_2835),
.B(n_2586),
.Y(n_3070)
);

CKINVDCx11_ASAP7_75t_R g3071 ( 
.A(n_2864),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_R g3072 ( 
.A(n_2765),
.B(n_746),
.Y(n_3072)
);

OR2x2_ASAP7_75t_L g3073 ( 
.A(n_2767),
.B(n_2665),
.Y(n_3073)
);

NAND2xp33_ASAP7_75t_R g3074 ( 
.A(n_2842),
.B(n_2609),
.Y(n_3074)
);

AND2x4_ASAP7_75t_L g3075 ( 
.A(n_2933),
.B(n_2459),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_R g3076 ( 
.A(n_2829),
.B(n_746),
.Y(n_3076)
);

OR2x4_ASAP7_75t_L g3077 ( 
.A(n_2770),
.B(n_2456),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2872),
.Y(n_3078)
);

NAND2xp33_ASAP7_75t_R g3079 ( 
.A(n_2847),
.B(n_2641),
.Y(n_3079)
);

XOR2xp5_ASAP7_75t_L g3080 ( 
.A(n_2845),
.B(n_2593),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_R g3081 ( 
.A(n_2846),
.B(n_747),
.Y(n_3081)
);

AND2x4_ASAP7_75t_L g3082 ( 
.A(n_2937),
.B(n_2886),
.Y(n_3082)
);

CKINVDCx5p33_ASAP7_75t_R g3083 ( 
.A(n_2924),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2874),
.Y(n_3084)
);

NAND2xp33_ASAP7_75t_R g3085 ( 
.A(n_2847),
.B(n_2641),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_2924),
.Y(n_3086)
);

NAND2xp33_ASAP7_75t_R g3087 ( 
.A(n_2906),
.B(n_2641),
.Y(n_3087)
);

BUFx3_ASAP7_75t_L g3088 ( 
.A(n_2914),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2876),
.Y(n_3089)
);

CKINVDCx11_ASAP7_75t_R g3090 ( 
.A(n_2916),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2756),
.B(n_2454),
.Y(n_3091)
);

AND2x4_ASAP7_75t_L g3092 ( 
.A(n_2961),
.B(n_2489),
.Y(n_3092)
);

AND2x4_ASAP7_75t_L g3093 ( 
.A(n_2976),
.B(n_2489),
.Y(n_3093)
);

OR2x4_ASAP7_75t_L g3094 ( 
.A(n_2999),
.B(n_2826),
.Y(n_3094)
);

OR2x4_ASAP7_75t_L g3095 ( 
.A(n_2786),
.B(n_2456),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_R g3096 ( 
.A(n_2782),
.B(n_748),
.Y(n_3096)
);

NAND2xp33_ASAP7_75t_R g3097 ( 
.A(n_2906),
.B(n_2706),
.Y(n_3097)
);

NAND2xp33_ASAP7_75t_R g3098 ( 
.A(n_2782),
.B(n_2792),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2989),
.B(n_2454),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2806),
.B(n_2674),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_2792),
.B(n_2706),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_R g3102 ( 
.A(n_2942),
.B(n_749),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2808),
.B(n_2646),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2815),
.B(n_2646),
.Y(n_3104)
);

INVxp67_ASAP7_75t_L g3105 ( 
.A(n_2923),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_R g3106 ( 
.A(n_2942),
.B(n_749),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2757),
.Y(n_3107)
);

AND2x4_ASAP7_75t_L g3108 ( 
.A(n_2858),
.B(n_2706),
.Y(n_3108)
);

CKINVDCx8_ASAP7_75t_R g3109 ( 
.A(n_2858),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2991),
.B(n_2478),
.Y(n_3110)
);

BUFx3_ASAP7_75t_L g3111 ( 
.A(n_2858),
.Y(n_3111)
);

INVxp67_ASAP7_75t_L g3112 ( 
.A(n_2936),
.Y(n_3112)
);

NAND2xp33_ASAP7_75t_R g3113 ( 
.A(n_2971),
.B(n_2711),
.Y(n_3113)
);

INVxp67_ASAP7_75t_L g3114 ( 
.A(n_2911),
.Y(n_3114)
);

NAND2xp33_ASAP7_75t_SL g3115 ( 
.A(n_2831),
.B(n_2570),
.Y(n_3115)
);

OR2x6_ASAP7_75t_L g3116 ( 
.A(n_2932),
.B(n_2711),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2759),
.Y(n_3117)
);

NAND2xp33_ASAP7_75t_R g3118 ( 
.A(n_2988),
.B(n_2711),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2816),
.B(n_2521),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2818),
.Y(n_3120)
);

XNOR2xp5_ASAP7_75t_L g3121 ( 
.A(n_2945),
.B(n_2629),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2819),
.Y(n_3122)
);

NOR2xp33_ASAP7_75t_L g3123 ( 
.A(n_2947),
.B(n_2458),
.Y(n_3123)
);

BUFx2_ASAP7_75t_SL g3124 ( 
.A(n_2954),
.Y(n_3124)
);

OR2x6_ASAP7_75t_L g3125 ( 
.A(n_2755),
.B(n_2738),
.Y(n_3125)
);

OR2x2_ASAP7_75t_L g3126 ( 
.A(n_2910),
.B(n_2741),
.Y(n_3126)
);

BUFx24_ASAP7_75t_SL g3127 ( 
.A(n_2945),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2992),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2938),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2751),
.B(n_2478),
.Y(n_3130)
);

NAND2xp33_ASAP7_75t_SL g3131 ( 
.A(n_2831),
.B(n_2680),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_2974),
.B(n_2773),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2952),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_R g3134 ( 
.A(n_2980),
.B(n_750),
.Y(n_3134)
);

NAND2xp33_ASAP7_75t_R g3135 ( 
.A(n_2866),
.B(n_2738),
.Y(n_3135)
);

NAND2xp33_ASAP7_75t_R g3136 ( 
.A(n_2866),
.B(n_2738),
.Y(n_3136)
);

XNOR2xp5_ASAP7_75t_L g3137 ( 
.A(n_2853),
.B(n_2543),
.Y(n_3137)
);

NAND2xp33_ASAP7_75t_R g3138 ( 
.A(n_2990),
.B(n_751),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2751),
.B(n_2482),
.Y(n_3139)
);

NAND2xp33_ASAP7_75t_R g3140 ( 
.A(n_2939),
.B(n_751),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_R g3141 ( 
.A(n_2980),
.B(n_752),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2938),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_2889),
.B(n_2487),
.Y(n_3143)
);

AND2x4_ASAP7_75t_L g3144 ( 
.A(n_2956),
.B(n_2500),
.Y(n_3144)
);

INVxp67_ASAP7_75t_L g3145 ( 
.A(n_2915),
.Y(n_3145)
);

NAND2xp33_ASAP7_75t_R g3146 ( 
.A(n_2921),
.B(n_753),
.Y(n_3146)
);

BUFx4f_ASAP7_75t_L g3147 ( 
.A(n_2952),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_2807),
.B(n_2675),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_R g3149 ( 
.A(n_2984),
.B(n_754),
.Y(n_3149)
);

CKINVDCx20_ASAP7_75t_R g3150 ( 
.A(n_2775),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2998),
.Y(n_3151)
);

BUFx3_ASAP7_75t_L g3152 ( 
.A(n_2953),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_2775),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_2807),
.B(n_2490),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2855),
.Y(n_3155)
);

NAND2xp33_ASAP7_75t_R g3156 ( 
.A(n_2957),
.B(n_754),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2841),
.B(n_2482),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2841),
.B(n_2492),
.Y(n_3158)
);

NAND2xp33_ASAP7_75t_R g3159 ( 
.A(n_2963),
.B(n_755),
.Y(n_3159)
);

AND2x4_ASAP7_75t_L g3160 ( 
.A(n_2859),
.B(n_2579),
.Y(n_3160)
);

BUFx24_ASAP7_75t_SL g3161 ( 
.A(n_2946),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2962),
.Y(n_3162)
);

NAND2xp33_ASAP7_75t_R g3163 ( 
.A(n_2984),
.B(n_755),
.Y(n_3163)
);

NAND2xp33_ASAP7_75t_R g3164 ( 
.A(n_2995),
.B(n_756),
.Y(n_3164)
);

CKINVDCx12_ASAP7_75t_R g3165 ( 
.A(n_2887),
.Y(n_3165)
);

BUFx3_ASAP7_75t_L g3166 ( 
.A(n_2987),
.Y(n_3166)
);

INVxp67_ASAP7_75t_L g3167 ( 
.A(n_2955),
.Y(n_3167)
);

OR2x4_ASAP7_75t_L g3168 ( 
.A(n_2965),
.B(n_2696),
.Y(n_3168)
);

OR2x2_ASAP7_75t_L g3169 ( 
.A(n_2918),
.B(n_2579),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_2859),
.B(n_2744),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_R g3171 ( 
.A(n_2995),
.B(n_756),
.Y(n_3171)
);

BUFx3_ASAP7_75t_L g3172 ( 
.A(n_2987),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_2849),
.B(n_2744),
.Y(n_3173)
);

OR2x2_ASAP7_75t_L g3174 ( 
.A(n_2885),
.B(n_2505),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_2805),
.B(n_2492),
.Y(n_3175)
);

NAND2xp33_ASAP7_75t_R g3176 ( 
.A(n_2917),
.B(n_757),
.Y(n_3176)
);

NAND2xp33_ASAP7_75t_SL g3177 ( 
.A(n_2791),
.B(n_2773),
.Y(n_3177)
);

AND2x4_ASAP7_75t_L g3178 ( 
.A(n_2850),
.B(n_2505),
.Y(n_3178)
);

AND2x4_ASAP7_75t_L g3179 ( 
.A(n_2868),
.B(n_2563),
.Y(n_3179)
);

INVxp67_ASAP7_75t_L g3180 ( 
.A(n_2892),
.Y(n_3180)
);

AND2x4_ASAP7_75t_L g3181 ( 
.A(n_2871),
.B(n_2563),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_2987),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_2917),
.B(n_2529),
.Y(n_3183)
);

BUFx3_ASAP7_75t_L g3184 ( 
.A(n_2973),
.Y(n_3184)
);

AND2x4_ASAP7_75t_L g3185 ( 
.A(n_2930),
.B(n_2796),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2998),
.Y(n_3186)
);

NAND2xp33_ASAP7_75t_R g3187 ( 
.A(n_2930),
.B(n_2986),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2769),
.B(n_2771),
.Y(n_3188)
);

NAND2xp33_ASAP7_75t_R g3189 ( 
.A(n_2839),
.B(n_758),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2856),
.Y(n_3190)
);

INVxp67_ASAP7_75t_L g3191 ( 
.A(n_2867),
.Y(n_3191)
);

OR2x2_ASAP7_75t_L g3192 ( 
.A(n_2878),
.B(n_2564),
.Y(n_3192)
);

XNOR2xp5_ASAP7_75t_L g3193 ( 
.A(n_2974),
.B(n_2723),
.Y(n_3193)
);

OR2x6_ASAP7_75t_L g3194 ( 
.A(n_2824),
.B(n_2698),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_R g3195 ( 
.A(n_2973),
.B(n_759),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2809),
.B(n_2601),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_R g3197 ( 
.A(n_2791),
.B(n_759),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_SL g3198 ( 
.A(n_2946),
.B(n_2567),
.Y(n_3198)
);

XNOR2xp5_ASAP7_75t_L g3199 ( 
.A(n_2883),
.B(n_2723),
.Y(n_3199)
);

NAND2xp33_ASAP7_75t_SL g3200 ( 
.A(n_2985),
.B(n_2680),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_2985),
.B(n_2567),
.Y(n_3201)
);

AND2x4_ASAP7_75t_L g3202 ( 
.A(n_2796),
.B(n_2468),
.Y(n_3202)
);

NAND2xp33_ASAP7_75t_R g3203 ( 
.A(n_2814),
.B(n_760),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2851),
.Y(n_3204)
);

CKINVDCx12_ASAP7_75t_R g3205 ( 
.A(n_2824),
.Y(n_3205)
);

INVxp67_ASAP7_75t_L g3206 ( 
.A(n_2873),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2772),
.B(n_2677),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_R g3208 ( 
.A(n_2860),
.B(n_760),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2774),
.B(n_2685),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2962),
.Y(n_3210)
);

XOR2x2_ASAP7_75t_SL g3211 ( 
.A(n_2983),
.B(n_2735),
.Y(n_3211)
);

INVxp67_ASAP7_75t_L g3212 ( 
.A(n_2798),
.Y(n_3212)
);

XNOR2xp5_ASAP7_75t_L g3213 ( 
.A(n_2844),
.B(n_2742),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_2830),
.B(n_2601),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2852),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2966),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_R g3217 ( 
.A(n_2860),
.B(n_761),
.Y(n_3217)
);

BUFx3_ASAP7_75t_L g3218 ( 
.A(n_2860),
.Y(n_3218)
);

CKINVDCx20_ASAP7_75t_R g3219 ( 
.A(n_2811),
.Y(n_3219)
);

XNOR2xp5_ASAP7_75t_L g3220 ( 
.A(n_2983),
.B(n_2742),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_R g3221 ( 
.A(n_2891),
.B(n_761),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2776),
.B(n_2604),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_R g3223 ( 
.A(n_2891),
.B(n_762),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2777),
.B(n_2604),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_2789),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_2836),
.B(n_2612),
.Y(n_3226)
);

AND2x2_ASAP7_75t_SL g3227 ( 
.A(n_3147),
.B(n_2789),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_3115),
.A2(n_2878),
.B1(n_2969),
.B2(n_2968),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3099),
.B(n_2827),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3155),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3057),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3009),
.Y(n_3232)
);

OR2x2_ASAP7_75t_L g3233 ( 
.A(n_3007),
.B(n_2799),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3078),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3084),
.Y(n_3235)
);

BUFx2_ASAP7_75t_SL g3236 ( 
.A(n_3034),
.Y(n_3236)
);

AOI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_3113),
.A2(n_2972),
.B1(n_2879),
.B2(n_2964),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3190),
.Y(n_3238)
);

AND2x4_ASAP7_75t_L g3239 ( 
.A(n_3048),
.B(n_2940),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3089),
.Y(n_3240)
);

BUFx3_ASAP7_75t_L g3241 ( 
.A(n_3058),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3031),
.B(n_2817),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3110),
.B(n_2832),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3024),
.B(n_2817),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3059),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3129),
.B(n_2838),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3188),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_3048),
.B(n_2940),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3120),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_SL g3250 ( 
.A1(n_3096),
.A2(n_2790),
.B1(n_2993),
.B2(n_2778),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_3020),
.B(n_2905),
.Y(n_3251)
);

INVx3_ASAP7_75t_L g3252 ( 
.A(n_3058),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_3112),
.B(n_2905),
.Y(n_3253)
);

INVx3_ASAP7_75t_L g3254 ( 
.A(n_3125),
.Y(n_3254)
);

OR2x2_ASAP7_75t_L g3255 ( 
.A(n_3212),
.B(n_2799),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3000),
.B(n_2912),
.Y(n_3256)
);

INVxp67_ASAP7_75t_SL g3257 ( 
.A(n_3225),
.Y(n_3257)
);

CKINVDCx11_ASAP7_75t_R g3258 ( 
.A(n_3019),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3193),
.A2(n_2934),
.B1(n_2964),
.B2(n_2879),
.Y(n_3259)
);

INVx3_ASAP7_75t_L g3260 ( 
.A(n_3125),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_3049),
.B(n_2897),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3122),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3117),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3142),
.B(n_2949),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3128),
.B(n_2912),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3061),
.B(n_2951),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3204),
.Y(n_3267)
);

BUFx3_ASAP7_75t_L g3268 ( 
.A(n_3018),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3039),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3030),
.B(n_2996),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3215),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3107),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3082),
.B(n_2996),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3001),
.B(n_2967),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3091),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_3063),
.B(n_2967),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_3199),
.A2(n_2934),
.B1(n_2875),
.B2(n_2780),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3063),
.B(n_2950),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3175),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_3002),
.B(n_2861),
.Y(n_3280)
);

INVxp67_ASAP7_75t_L g3281 ( 
.A(n_3069),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3043),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3165),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3052),
.B(n_2958),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3037),
.B(n_3053),
.Y(n_3285)
);

OR2x2_ASAP7_75t_L g3286 ( 
.A(n_3206),
.B(n_3073),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3151),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3070),
.B(n_2862),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3162),
.Y(n_3289)
);

OAI21xp33_ASAP7_75t_L g3290 ( 
.A1(n_3021),
.A2(n_2780),
.B(n_2875),
.Y(n_3290)
);

AND2x6_ASAP7_75t_SL g3291 ( 
.A(n_3054),
.B(n_2824),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3114),
.B(n_2893),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3145),
.B(n_2895),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3152),
.B(n_2901),
.Y(n_3294)
);

OR2x2_ASAP7_75t_L g3295 ( 
.A(n_3186),
.B(n_2825),
.Y(n_3295)
);

BUFx2_ASAP7_75t_L g3296 ( 
.A(n_3111),
.Y(n_3296)
);

OR2x2_ASAP7_75t_L g3297 ( 
.A(n_3210),
.B(n_2825),
.Y(n_3297)
);

BUFx2_ASAP7_75t_L g3298 ( 
.A(n_3018),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3216),
.Y(n_3299)
);

OR2x2_ASAP7_75t_L g3300 ( 
.A(n_3192),
.B(n_2865),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3116),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3116),
.Y(n_3302)
);

OR2x2_ASAP7_75t_L g3303 ( 
.A(n_3174),
.B(n_2865),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3180),
.B(n_3191),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3049),
.B(n_2902),
.Y(n_3305)
);

INVxp67_ASAP7_75t_L g3306 ( 
.A(n_3074),
.Y(n_3306)
);

OR2x2_ASAP7_75t_L g3307 ( 
.A(n_3226),
.B(n_2922),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3075),
.B(n_2904),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_3105),
.B(n_2943),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3196),
.B(n_2948),
.Y(n_3310)
);

AOI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_3132),
.A2(n_2823),
.B1(n_2820),
.B2(n_2926),
.Y(n_3311)
);

INVx4_ASAP7_75t_R g3312 ( 
.A(n_3055),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3139),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3157),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3214),
.B(n_2920),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3064),
.B(n_2899),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_3131),
.B(n_2896),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_3064),
.B(n_2903),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3092),
.B(n_2907),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3158),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3100),
.B(n_2925),
.Y(n_3321)
);

HB1xp67_ASAP7_75t_L g3322 ( 
.A(n_3130),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3088),
.B(n_2922),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3066),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3093),
.B(n_2908),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3222),
.Y(n_3326)
);

BUFx2_ASAP7_75t_SL g3327 ( 
.A(n_3109),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3066),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3202),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3185),
.B(n_3133),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3285),
.B(n_3153),
.Y(n_3331)
);

NAND3xp33_ASAP7_75t_SL g3332 ( 
.A(n_3290),
.B(n_3040),
.C(n_3072),
.Y(n_3332)
);

AOI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_3277),
.A2(n_3118),
.B1(n_3136),
.B2(n_3135),
.Y(n_3333)
);

AO21x2_ASAP7_75t_L g3334 ( 
.A1(n_3317),
.A2(n_3198),
.B(n_2888),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3301),
.B(n_3090),
.Y(n_3335)
);

INVx1_ASAP7_75t_SL g3336 ( 
.A(n_3236),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3231),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3230),
.Y(n_3338)
);

AND2x2_ASAP7_75t_L g3339 ( 
.A(n_3302),
.B(n_3276),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3326),
.B(n_2975),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_3277),
.A2(n_3177),
.B1(n_3259),
.B2(n_3250),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_3244),
.B(n_3150),
.Y(n_3342)
);

OR2x6_ASAP7_75t_L g3343 ( 
.A(n_3254),
.B(n_3194),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_3312),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3242),
.B(n_3011),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3230),
.Y(n_3346)
);

OAI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3237),
.A2(n_3077),
.B1(n_3095),
.B2(n_3220),
.Y(n_3347)
);

HB1xp67_ASAP7_75t_L g3348 ( 
.A(n_3322),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3274),
.B(n_3025),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3273),
.B(n_3154),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3259),
.A2(n_3201),
.B1(n_3200),
.B2(n_3127),
.Y(n_3351)
);

BUFx2_ASAP7_75t_L g3352 ( 
.A(n_3241),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3232),
.Y(n_3353)
);

BUFx3_ASAP7_75t_L g3354 ( 
.A(n_3258),
.Y(n_3354)
);

NAND3xp33_ASAP7_75t_L g3355 ( 
.A(n_3317),
.B(n_3062),
.C(n_3056),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3330),
.B(n_3170),
.Y(n_3356)
);

OAI31xp33_ASAP7_75t_L g3357 ( 
.A1(n_3281),
.A2(n_3121),
.A3(n_3041),
.B(n_3060),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3238),
.Y(n_3358)
);

OR2x6_ASAP7_75t_L g3359 ( 
.A(n_3254),
.B(n_3194),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3234),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3269),
.B(n_2978),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3270),
.B(n_3023),
.Y(n_3362)
);

OAI21xp33_ASAP7_75t_L g3363 ( 
.A1(n_3281),
.A2(n_3051),
.B(n_3081),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3279),
.B(n_3144),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3235),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3240),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3279),
.B(n_3108),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_3322),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3282),
.B(n_3247),
.Y(n_3369)
);

AND2x4_ASAP7_75t_SL g3370 ( 
.A(n_3252),
.B(n_3042),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3287),
.B(n_2928),
.Y(n_3371)
);

AOI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3250),
.A2(n_3187),
.B1(n_3138),
.B2(n_3189),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3245),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3289),
.B(n_2929),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3249),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3251),
.B(n_3160),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_3239),
.B(n_3179),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3288),
.B(n_3173),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3299),
.B(n_2931),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_3257),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3262),
.Y(n_3381)
);

INVx3_ASAP7_75t_L g3382 ( 
.A(n_3241),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_3283),
.B(n_3017),
.Y(n_3383)
);

AO21x2_ASAP7_75t_L g3384 ( 
.A1(n_3306),
.A2(n_2982),
.B(n_2966),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3263),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3323),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3255),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3238),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3286),
.Y(n_3389)
);

OAI31xp33_ASAP7_75t_SL g3390 ( 
.A1(n_3239),
.A2(n_3015),
.A3(n_3101),
.B(n_3213),
.Y(n_3390)
);

INVx4_ASAP7_75t_L g3391 ( 
.A(n_3258),
.Y(n_3391)
);

AOI31xp33_ASAP7_75t_L g3392 ( 
.A1(n_3306),
.A2(n_3098),
.A3(n_3097),
.B(n_3087),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3257),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3253),
.B(n_3181),
.Y(n_3394)
);

NOR3xp33_ASAP7_75t_L g3395 ( 
.A(n_3252),
.B(n_2993),
.C(n_2833),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_3327),
.B(n_3094),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3275),
.B(n_3178),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3271),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3256),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3275),
.B(n_3027),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3227),
.A2(n_3050),
.B(n_3038),
.Y(n_3401)
);

NAND2x1_ASAP7_75t_L g3402 ( 
.A(n_3260),
.B(n_3042),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3271),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3233),
.Y(n_3404)
);

HB1xp67_ASAP7_75t_L g3405 ( 
.A(n_3313),
.Y(n_3405)
);

INVxp67_ASAP7_75t_L g3406 ( 
.A(n_3296),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_3309),
.B(n_3166),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3272),
.Y(n_3408)
);

OR2x2_ASAP7_75t_L g3409 ( 
.A(n_3307),
.B(n_2997),
.Y(n_3409)
);

HB1xp67_ASAP7_75t_L g3410 ( 
.A(n_3313),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3308),
.B(n_3172),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3305),
.B(n_3124),
.Y(n_3412)
);

HB1xp67_ASAP7_75t_L g3413 ( 
.A(n_3314),
.Y(n_3413)
);

CKINVDCx20_ASAP7_75t_R g3414 ( 
.A(n_3354),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3387),
.B(n_3228),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_SL g3416 ( 
.A(n_3390),
.B(n_3227),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3369),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3340),
.B(n_3315),
.Y(n_3418)
);

OR2x2_ASAP7_75t_L g3419 ( 
.A(n_3348),
.B(n_3315),
.Y(n_3419)
);

OR2x2_ASAP7_75t_L g3420 ( 
.A(n_3348),
.B(n_3266),
.Y(n_3420)
);

OR2x2_ASAP7_75t_L g3421 ( 
.A(n_3368),
.B(n_3266),
.Y(n_3421)
);

AND2x4_ASAP7_75t_SL g3422 ( 
.A(n_3391),
.B(n_3294),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3350),
.B(n_3248),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3356),
.B(n_3248),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3393),
.B(n_3284),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3369),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3337),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3376),
.B(n_3304),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3353),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3386),
.B(n_3284),
.Y(n_3430)
);

INVx1_ASAP7_75t_SL g3431 ( 
.A(n_3336),
.Y(n_3431)
);

INVx4_ASAP7_75t_L g3432 ( 
.A(n_3391),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3340),
.B(n_3321),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3336),
.B(n_3071),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3389),
.B(n_3229),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3394),
.B(n_3260),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3343),
.B(n_3261),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_3378),
.B(n_3292),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3360),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3368),
.Y(n_3440)
);

HB1xp67_ASAP7_75t_L g3441 ( 
.A(n_3380),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3362),
.B(n_3293),
.Y(n_3442)
);

BUFx2_ASAP7_75t_SL g3443 ( 
.A(n_3344),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3365),
.Y(n_3444)
);

AOI22xp33_ASAP7_75t_L g3445 ( 
.A1(n_3347),
.A2(n_3311),
.B1(n_3161),
.B2(n_3183),
.Y(n_3445)
);

AND2x4_ASAP7_75t_L g3446 ( 
.A(n_3343),
.B(n_3261),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3361),
.B(n_3321),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3404),
.B(n_3229),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3399),
.B(n_3243),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3366),
.Y(n_3450)
);

INVxp67_ASAP7_75t_L g3451 ( 
.A(n_3352),
.Y(n_3451)
);

HB1xp67_ASAP7_75t_L g3452 ( 
.A(n_3405),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3361),
.B(n_3243),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3405),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3373),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3375),
.Y(n_3456)
);

HB1xp67_ASAP7_75t_L g3457 ( 
.A(n_3410),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3409),
.B(n_3310),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3381),
.B(n_3300),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3410),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3377),
.B(n_3324),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3385),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3371),
.Y(n_3463)
);

OR2x2_ASAP7_75t_L g3464 ( 
.A(n_3413),
.B(n_3314),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3371),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3374),
.Y(n_3466)
);

NAND2x1p5_ASAP7_75t_L g3467 ( 
.A(n_3402),
.B(n_3268),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3341),
.B(n_3311),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3374),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3413),
.Y(n_3470)
);

OR2x2_ASAP7_75t_L g3471 ( 
.A(n_3338),
.B(n_3320),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3351),
.B(n_3265),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3377),
.B(n_3324),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3347),
.B(n_3400),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3379),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3379),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3334),
.B(n_3246),
.Y(n_3477)
);

INVxp67_ASAP7_75t_SL g3478 ( 
.A(n_3406),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_3383),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3346),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3358),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3407),
.B(n_3328),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3345),
.B(n_3328),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3388),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_3416),
.B(n_3390),
.Y(n_3485)
);

NAND2xp33_ASAP7_75t_SL g3486 ( 
.A(n_3432),
.B(n_3044),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3417),
.B(n_3334),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3426),
.B(n_3333),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3419),
.B(n_3406),
.Y(n_3489)
);

AO221x2_ASAP7_75t_L g3490 ( 
.A1(n_3474),
.A2(n_3080),
.B1(n_3355),
.B2(n_3392),
.C(n_3022),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_3414),
.Y(n_3491)
);

OR2x2_ASAP7_75t_L g3492 ( 
.A(n_3420),
.B(n_3320),
.Y(n_3492)
);

NOR2x1_ASAP7_75t_L g3493 ( 
.A(n_3432),
.B(n_3332),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3463),
.B(n_3401),
.Y(n_3494)
);

INVxp67_ASAP7_75t_L g3495 ( 
.A(n_3431),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3465),
.B(n_3401),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3466),
.B(n_3384),
.Y(n_3497)
);

CKINVDCx5p33_ASAP7_75t_R g3498 ( 
.A(n_3443),
.Y(n_3498)
);

NAND2xp33_ASAP7_75t_R g3499 ( 
.A(n_3437),
.B(n_3102),
.Y(n_3499)
);

NOR2x1_ASAP7_75t_L g3500 ( 
.A(n_3431),
.B(n_3332),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3469),
.B(n_3384),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3421),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_3434),
.B(n_3396),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3475),
.B(n_3395),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3437),
.B(n_3349),
.Y(n_3505)
);

AND2x4_ASAP7_75t_L g3506 ( 
.A(n_3422),
.B(n_3343),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3476),
.B(n_3395),
.Y(n_3507)
);

AO221x2_ASAP7_75t_L g3508 ( 
.A1(n_3468),
.A2(n_3392),
.B1(n_3357),
.B2(n_3016),
.C(n_3010),
.Y(n_3508)
);

NAND2xp33_ASAP7_75t_SL g3509 ( 
.A(n_3446),
.B(n_3106),
.Y(n_3509)
);

AO221x2_ASAP7_75t_L g3510 ( 
.A1(n_3472),
.A2(n_3006),
.B1(n_3446),
.B2(n_3363),
.C(n_3415),
.Y(n_3510)
);

AO221x2_ASAP7_75t_L g3511 ( 
.A1(n_3477),
.A2(n_3291),
.B1(n_3012),
.B2(n_3014),
.C(n_3372),
.Y(n_3511)
);

BUFx2_ASAP7_75t_L g3512 ( 
.A(n_3441),
.Y(n_3512)
);

NAND2xp33_ASAP7_75t_SL g3513 ( 
.A(n_3452),
.B(n_3068),
.Y(n_3513)
);

OAI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3478),
.A2(n_3359),
.B1(n_3382),
.B2(n_3085),
.Y(n_3514)
);

NAND2xp33_ASAP7_75t_SL g3515 ( 
.A(n_3457),
.B(n_3046),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_R g3516 ( 
.A(n_3479),
.B(n_3163),
.Y(n_3516)
);

BUFx2_ASAP7_75t_L g3517 ( 
.A(n_3467),
.Y(n_3517)
);

AO221x2_ASAP7_75t_L g3518 ( 
.A1(n_3477),
.A2(n_3458),
.B1(n_3036),
.B2(n_3140),
.C(n_3454),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_3451),
.Y(n_3519)
);

NAND2xp33_ASAP7_75t_SL g3520 ( 
.A(n_3440),
.B(n_3412),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3433),
.B(n_3397),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3433),
.B(n_3280),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3447),
.B(n_3278),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_SL g3524 ( 
.A(n_3467),
.B(n_3083),
.Y(n_3524)
);

CKINVDCx5p33_ASAP7_75t_R g3525 ( 
.A(n_3436),
.Y(n_3525)
);

OAI221xp5_ASAP7_75t_L g3526 ( 
.A1(n_3445),
.A2(n_3164),
.B1(n_3359),
.B2(n_3176),
.C(n_3382),
.Y(n_3526)
);

NOR2x1_ASAP7_75t_L g3527 ( 
.A(n_3460),
.B(n_3359),
.Y(n_3527)
);

OAI221xp5_ASAP7_75t_L g3528 ( 
.A1(n_3447),
.A2(n_3167),
.B1(n_3013),
.B2(n_3156),
.C(n_3159),
.Y(n_3528)
);

HB1xp67_ASAP7_75t_L g3529 ( 
.A(n_3470),
.Y(n_3529)
);

AO221x2_ASAP7_75t_L g3530 ( 
.A1(n_3448),
.A2(n_3008),
.B1(n_3146),
.B2(n_3086),
.C(n_3003),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_3459),
.B(n_3335),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3424),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3418),
.B(n_3339),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3512),
.Y(n_3534)
);

NOR2x1_ASAP7_75t_L g3535 ( 
.A(n_3493),
.B(n_3004),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3489),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3495),
.Y(n_3537)
);

AOI22xp33_ASAP7_75t_L g3538 ( 
.A1(n_3508),
.A2(n_3123),
.B1(n_3435),
.B2(n_3076),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3511),
.B(n_3490),
.Y(n_3539)
);

AOI22xp33_ASAP7_75t_SL g3540 ( 
.A1(n_3530),
.A2(n_3141),
.B1(n_3149),
.B2(n_3134),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_3508),
.A2(n_3430),
.B1(n_3449),
.B2(n_3418),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3502),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3504),
.B(n_3453),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3492),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3507),
.B(n_3427),
.Y(n_3545)
);

CKINVDCx16_ASAP7_75t_R g3546 ( 
.A(n_3486),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_3494),
.B(n_3425),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3490),
.A2(n_3485),
.B1(n_3511),
.B2(n_3518),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3518),
.A2(n_3459),
.B1(n_3473),
.B2(n_3461),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3523),
.Y(n_3550)
);

OAI21x1_ASAP7_75t_L g3551 ( 
.A1(n_3527),
.A2(n_3464),
.B(n_3439),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3529),
.Y(n_3552)
);

INVxp67_ASAP7_75t_L g3553 ( 
.A(n_3500),
.Y(n_3553)
);

HB1xp67_ASAP7_75t_L g3554 ( 
.A(n_3496),
.Y(n_3554)
);

CKINVDCx16_ASAP7_75t_R g3555 ( 
.A(n_3499),
.Y(n_3555)
);

AND3x1_ASAP7_75t_L g3556 ( 
.A(n_3524),
.B(n_3342),
.C(n_3331),
.Y(n_3556)
);

OAI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3487),
.A2(n_3444),
.B(n_3429),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3510),
.A2(n_3195),
.B1(n_3217),
.B2(n_3208),
.Y(n_3558)
);

BUFx3_ASAP7_75t_L g3559 ( 
.A(n_3491),
.Y(n_3559)
);

OR2x2_ASAP7_75t_L g3560 ( 
.A(n_3520),
.B(n_3488),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3517),
.B(n_3423),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3497),
.B(n_3450),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3521),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3501),
.B(n_3455),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3510),
.A2(n_3223),
.B1(n_3221),
.B2(n_3303),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3506),
.B(n_3428),
.Y(n_3566)
);

OR2x2_ASAP7_75t_L g3567 ( 
.A(n_3522),
.B(n_3471),
.Y(n_3567)
);

OR2x2_ASAP7_75t_L g3568 ( 
.A(n_3533),
.B(n_3480),
.Y(n_3568)
);

AND2x2_ASAP7_75t_L g3569 ( 
.A(n_3505),
.B(n_3482),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3498),
.Y(n_3570)
);

NAND3xp33_ASAP7_75t_L g3571 ( 
.A(n_3509),
.B(n_3203),
.C(n_3456),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3519),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3531),
.B(n_3462),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3503),
.B(n_3438),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3532),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3530),
.B(n_3483),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3514),
.B(n_3481),
.Y(n_3577)
);

NOR2x1_ASAP7_75t_L g3578 ( 
.A(n_3526),
.B(n_3219),
.Y(n_3578)
);

OR2x2_ASAP7_75t_L g3579 ( 
.A(n_3513),
.B(n_3484),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_3515),
.A2(n_3411),
.B1(n_3367),
.B2(n_3318),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3525),
.Y(n_3581)
);

HB1xp67_ASAP7_75t_L g3582 ( 
.A(n_3516),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3528),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3511),
.B(n_3442),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3504),
.B(n_3398),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3554),
.B(n_3316),
.Y(n_3586)
);

OAI322xp33_ASAP7_75t_L g3587 ( 
.A1(n_3553),
.A2(n_3297),
.A3(n_3295),
.B1(n_3137),
.B2(n_3126),
.C1(n_3079),
.C2(n_3104),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3554),
.B(n_3319),
.Y(n_3588)
);

AOI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_3539),
.A2(n_3205),
.B1(n_3143),
.B2(n_3026),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3534),
.B(n_3325),
.Y(n_3590)
);

OA211x2_ASAP7_75t_L g3591 ( 
.A1(n_3548),
.A2(n_3565),
.B(n_3571),
.C(n_3538),
.Y(n_3591)
);

INVx3_ASAP7_75t_L g3592 ( 
.A(n_3556),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_L g3593 ( 
.A(n_3555),
.B(n_3370),
.Y(n_3593)
);

AOI32xp33_ASAP7_75t_L g3594 ( 
.A1(n_3578),
.A2(n_3364),
.A3(n_3005),
.B1(n_3211),
.B2(n_2784),
.Y(n_3594)
);

OAI322xp33_ASAP7_75t_L g3595 ( 
.A1(n_3553),
.A2(n_3103),
.A3(n_3033),
.B1(n_3224),
.B2(n_3032),
.C1(n_3029),
.C2(n_3028),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3546),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3583),
.B(n_3403),
.Y(n_3597)
);

OAI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3549),
.A2(n_3541),
.B1(n_3558),
.B2(n_3540),
.Y(n_3598)
);

OAI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3582),
.A2(n_2854),
.B(n_2833),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3559),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3584),
.B(n_3298),
.Y(n_3601)
);

OR2x2_ASAP7_75t_L g3602 ( 
.A(n_3543),
.B(n_3408),
.Y(n_3602)
);

AOI221xp5_ASAP7_75t_L g3603 ( 
.A1(n_3582),
.A2(n_3171),
.B1(n_2784),
.B2(n_2508),
.C(n_3197),
.Y(n_3603)
);

AOI221xp5_ASAP7_75t_L g3604 ( 
.A1(n_3537),
.A2(n_3246),
.B1(n_2821),
.B2(n_3264),
.C(n_2781),
.Y(n_3604)
);

OAI22xp33_ASAP7_75t_L g3605 ( 
.A1(n_3560),
.A2(n_3168),
.B1(n_3047),
.B2(n_3045),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3536),
.Y(n_3606)
);

AOI32xp33_ASAP7_75t_L g3607 ( 
.A1(n_3540),
.A2(n_2848),
.A3(n_3329),
.B1(n_3148),
.B2(n_2821),
.Y(n_3607)
);

AOI211xp5_ASAP7_75t_L g3608 ( 
.A1(n_3576),
.A2(n_2882),
.B(n_2854),
.C(n_2722),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3585),
.Y(n_3609)
);

NOR3xp33_ASAP7_75t_L g3610 ( 
.A(n_3535),
.B(n_2719),
.C(n_2722),
.Y(n_3610)
);

OAI32xp33_ASAP7_75t_L g3611 ( 
.A1(n_3577),
.A2(n_3067),
.A3(n_3065),
.B1(n_3268),
.B2(n_3169),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3585),
.Y(n_3612)
);

AOI221xp5_ASAP7_75t_L g3613 ( 
.A1(n_3545),
.A2(n_3264),
.B1(n_2785),
.B2(n_2788),
.C(n_2787),
.Y(n_3613)
);

OAI211xp5_ASAP7_75t_SL g3614 ( 
.A1(n_3572),
.A2(n_3581),
.B(n_3570),
.C(n_3575),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3563),
.B(n_3267),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3568),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_3572),
.B(n_3566),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3561),
.B(n_3329),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3600),
.B(n_3545),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3596),
.B(n_3574),
.Y(n_3620)
);

NAND3x1_ASAP7_75t_L g3621 ( 
.A(n_3592),
.B(n_3573),
.C(n_3542),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3616),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3597),
.Y(n_3623)
);

OR2x2_ASAP7_75t_L g3624 ( 
.A(n_3609),
.B(n_3612),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3592),
.A2(n_3547),
.B1(n_3550),
.B2(n_3552),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3617),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3599),
.B(n_3573),
.Y(n_3627)
);

NOR2x1_ASAP7_75t_L g3628 ( 
.A(n_3614),
.B(n_3579),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3586),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3615),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3606),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3604),
.B(n_3562),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3588),
.Y(n_3633)
);

AND2x4_ASAP7_75t_SL g3634 ( 
.A(n_3593),
.B(n_3580),
.Y(n_3634)
);

INVx2_ASAP7_75t_SL g3635 ( 
.A(n_3601),
.Y(n_3635)
);

AND2x2_ASAP7_75t_L g3636 ( 
.A(n_3618),
.B(n_3569),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3602),
.Y(n_3637)
);

OR2x2_ASAP7_75t_L g3638 ( 
.A(n_3598),
.B(n_3562),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3590),
.Y(n_3639)
);

INVx3_ASAP7_75t_L g3640 ( 
.A(n_3591),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3587),
.Y(n_3641)
);

AND2x4_ASAP7_75t_L g3642 ( 
.A(n_3589),
.B(n_3551),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3613),
.Y(n_3643)
);

INVx1_ASAP7_75t_SL g3644 ( 
.A(n_3607),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3637),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3619),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3637),
.Y(n_3647)
);

HB1xp67_ASAP7_75t_SL g3648 ( 
.A(n_3626),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3624),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3623),
.Y(n_3650)
);

BUFx4f_ASAP7_75t_SL g3651 ( 
.A(n_3640),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3630),
.Y(n_3652)
);

INVxp33_ASAP7_75t_L g3653 ( 
.A(n_3620),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3622),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3631),
.Y(n_3655)
);

CKINVDCx5p33_ASAP7_75t_R g3656 ( 
.A(n_3640),
.Y(n_3656)
);

BUFx8_ASAP7_75t_SL g3657 ( 
.A(n_3633),
.Y(n_3657)
);

CKINVDCx20_ASAP7_75t_R g3658 ( 
.A(n_3634),
.Y(n_3658)
);

INVx1_ASAP7_75t_SL g3659 ( 
.A(n_3621),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3629),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3639),
.Y(n_3661)
);

BUFx4f_ASAP7_75t_SL g3662 ( 
.A(n_3638),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3635),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3627),
.Y(n_3664)
);

XOR2x2_ASAP7_75t_L g3665 ( 
.A(n_3641),
.B(n_3610),
.Y(n_3665)
);

INVxp33_ASAP7_75t_SL g3666 ( 
.A(n_3625),
.Y(n_3666)
);

NAND3xp33_ASAP7_75t_SL g3667 ( 
.A(n_3656),
.B(n_3644),
.C(n_3594),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3666),
.A2(n_3628),
.B(n_3632),
.Y(n_3668)
);

NOR2xp67_ASAP7_75t_SL g3669 ( 
.A(n_3651),
.B(n_3643),
.Y(n_3669)
);

AOI221xp5_ASAP7_75t_L g3670 ( 
.A1(n_3653),
.A2(n_3642),
.B1(n_3611),
.B2(n_3595),
.C(n_3603),
.Y(n_3670)
);

INVxp67_ASAP7_75t_L g3671 ( 
.A(n_3648),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3648),
.Y(n_3672)
);

NAND4xp25_ASAP7_75t_L g3673 ( 
.A(n_3663),
.B(n_3642),
.C(n_3608),
.D(n_3636),
.Y(n_3673)
);

OAI221xp5_ASAP7_75t_L g3674 ( 
.A1(n_3659),
.A2(n_3564),
.B1(n_2502),
.B2(n_3544),
.C(n_3567),
.Y(n_3674)
);

OAI211xp5_ASAP7_75t_L g3675 ( 
.A1(n_3658),
.A2(n_3564),
.B(n_2476),
.C(n_2486),
.Y(n_3675)
);

NOR3x1_ASAP7_75t_L g3676 ( 
.A(n_3646),
.B(n_3557),
.C(n_2719),
.Y(n_3676)
);

AOI311xp33_ASAP7_75t_L g3677 ( 
.A1(n_3664),
.A2(n_3605),
.A3(n_2581),
.B(n_2635),
.C(n_2794),
.Y(n_3677)
);

NOR4xp25_ASAP7_75t_L g3678 ( 
.A(n_3650),
.B(n_2731),
.C(n_2491),
.D(n_2461),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_3665),
.A2(n_3645),
.B(n_3647),
.Y(n_3679)
);

NOR2xp67_ASAP7_75t_L g3680 ( 
.A(n_3649),
.B(n_763),
.Y(n_3680)
);

NAND4xp25_ASAP7_75t_L g3681 ( 
.A(n_3668),
.B(n_3660),
.C(n_3661),
.D(n_3652),
.Y(n_3681)
);

XNOR2xp5_ASAP7_75t_L g3682 ( 
.A(n_3667),
.B(n_3654),
.Y(n_3682)
);

OAI211xp5_ASAP7_75t_SL g3683 ( 
.A1(n_3671),
.A2(n_3655),
.B(n_3662),
.C(n_3657),
.Y(n_3683)
);

NAND4xp25_ASAP7_75t_L g3684 ( 
.A(n_3672),
.B(n_3662),
.C(n_2467),
.D(n_2581),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_L g3685 ( 
.A1(n_3669),
.A2(n_3184),
.B1(n_3182),
.B2(n_2848),
.Y(n_3685)
);

AOI211xp5_ASAP7_75t_L g3686 ( 
.A1(n_3679),
.A2(n_2678),
.B(n_2687),
.C(n_2728),
.Y(n_3686)
);

OAI211xp5_ASAP7_75t_SL g3687 ( 
.A1(n_3670),
.A2(n_2678),
.B(n_2728),
.C(n_2687),
.Y(n_3687)
);

AOI22xp5_ASAP7_75t_SL g3688 ( 
.A1(n_3676),
.A2(n_2549),
.B1(n_2653),
.B2(n_2636),
.Y(n_3688)
);

AOI22xp5_ASAP7_75t_L g3689 ( 
.A1(n_3673),
.A2(n_3119),
.B1(n_3209),
.B2(n_3207),
.Y(n_3689)
);

NAND3xp33_ASAP7_75t_L g3690 ( 
.A(n_3680),
.B(n_3677),
.C(n_3674),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3675),
.Y(n_3691)
);

XNOR2xp5_ASAP7_75t_L g3692 ( 
.A(n_3678),
.B(n_763),
.Y(n_3692)
);

BUFx2_ASAP7_75t_L g3693 ( 
.A(n_3692),
.Y(n_3693)
);

XOR2x2_ASAP7_75t_L g3694 ( 
.A(n_3682),
.B(n_3690),
.Y(n_3694)
);

AO22x1_ASAP7_75t_L g3695 ( 
.A1(n_3691),
.A2(n_2549),
.B1(n_2653),
.B2(n_2636),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3683),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3689),
.Y(n_3697)
);

XNOR2xp5_ASAP7_75t_L g3698 ( 
.A(n_3684),
.B(n_764),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3687),
.A2(n_3218),
.B1(n_2944),
.B2(n_3035),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3688),
.B(n_2548),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_R g3701 ( 
.A(n_3696),
.B(n_764),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_R g3702 ( 
.A(n_3698),
.B(n_765),
.Y(n_3702)
);

NOR2xp33_ASAP7_75t_R g3703 ( 
.A(n_3693),
.B(n_3697),
.Y(n_3703)
);

OAI221xp5_ASAP7_75t_L g3704 ( 
.A1(n_3703),
.A2(n_3681),
.B1(n_3700),
.B2(n_3694),
.C(n_3686),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3702),
.B(n_3685),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3701),
.Y(n_3706)
);

OAI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3704),
.A2(n_3699),
.B1(n_3695),
.B2(n_2840),
.Y(n_3707)
);

OAI22xp5_ASAP7_75t_SL g3708 ( 
.A1(n_3707),
.A2(n_3706),
.B1(n_3705),
.B2(n_2572),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_L g3709 ( 
.A1(n_3708),
.A2(n_2944),
.B1(n_2979),
.B2(n_2977),
.Y(n_3709)
);

OAI322xp33_ASAP7_75t_L g3710 ( 
.A1(n_3709),
.A2(n_2594),
.A3(n_2600),
.B1(n_2510),
.B2(n_2635),
.C1(n_2453),
.C2(n_2452),
.Y(n_3710)
);

AO221x1_ASAP7_75t_L g3711 ( 
.A1(n_3710),
.A2(n_2714),
.B1(n_2882),
.B2(n_2800),
.C(n_2783),
.Y(n_3711)
);

INVxp67_ASAP7_75t_SL g3712 ( 
.A(n_3711),
.Y(n_3712)
);

OAI221xp5_ASAP7_75t_R g3713 ( 
.A1(n_3712),
.A2(n_765),
.B1(n_766),
.B2(n_767),
.C(n_768),
.Y(n_3713)
);

AOI211xp5_ASAP7_75t_L g3714 ( 
.A1(n_3713),
.A2(n_2557),
.B(n_2600),
.C(n_2594),
.Y(n_3714)
);


endmodule