module fake_jpeg_4048_n_43 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_22),
.B(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_19),
.B(n_23),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_31),
.B1(n_29),
.B2(n_22),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_21),
.B(n_25),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_26),
.Y(n_36)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_29),
.B1(n_24),
.B2(n_17),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_33),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_10),
.B(n_17),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_6),
.Y(n_38)
);

OAI21x1_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_6),
.B(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

AOI321xp33_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_10),
.A3(n_13),
.B1(n_7),
.B2(n_9),
.C(n_4),
.Y(n_42)
);

OAI31xp33_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.A3(n_9),
.B(n_0),
.Y(n_43)
);


endmodule