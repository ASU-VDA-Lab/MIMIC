module real_aes_1511_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g517 ( .A(n_0), .B(n_214), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_1), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g148 ( .A(n_2), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_3), .B(n_520), .Y(n_539) );
NAND2xp33_ASAP7_75t_SL g510 ( .A(n_4), .B(n_169), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_5), .B(n_182), .Y(n_205) );
INVx1_ASAP7_75t_L g502 ( .A(n_6), .Y(n_502) );
INVx1_ASAP7_75t_L g239 ( .A(n_7), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g794 ( .A(n_8), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_9), .Y(n_256) );
AND2x2_ASAP7_75t_L g537 ( .A(n_10), .B(n_138), .Y(n_537) );
INVx2_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g215 ( .A(n_13), .Y(n_215) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_14), .A2(n_105), .B1(n_787), .B2(n_798), .C(n_805), .Y(n_104) );
AOI221x1_ASAP7_75t_L g505 ( .A1(n_14), .A2(n_171), .B1(n_506), .B2(n_508), .C(n_509), .Y(n_505) );
OAI22xp5_ASAP7_75t_SL g807 ( .A1(n_14), .A2(n_58), .B1(n_808), .B2(n_809), .Y(n_807) );
INVxp67_ASAP7_75t_L g809 ( .A(n_14), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_15), .B(n_520), .Y(n_573) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVx1_ASAP7_75t_L g212 ( .A(n_17), .Y(n_212) );
INVx1_ASAP7_75t_SL g160 ( .A(n_18), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_19), .B(n_163), .Y(n_185) );
AOI33xp33_ASAP7_75t_L g230 ( .A1(n_20), .A2(n_48), .A3(n_145), .B1(n_156), .B2(n_231), .B3(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_508), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_22), .B(n_214), .Y(n_542) );
AOI221xp5_ASAP7_75t_SL g582 ( .A1(n_23), .A2(n_39), .B1(n_508), .B2(n_520), .C(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g249 ( .A(n_24), .Y(n_249) );
OR2x2_ASAP7_75t_L g140 ( .A(n_25), .B(n_92), .Y(n_140) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_25), .A2(n_92), .B(n_139), .Y(n_173) );
INVxp67_ASAP7_75t_L g504 ( .A(n_26), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_27), .B(n_217), .Y(n_577) );
AND2x2_ASAP7_75t_L g531 ( .A(n_28), .B(n_137), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_29), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_30), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_31), .A2(n_508), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_32), .B(n_217), .Y(n_584) );
AND2x2_ASAP7_75t_L g150 ( .A(n_33), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g155 ( .A(n_33), .Y(n_155) );
AND2x2_ASAP7_75t_L g169 ( .A(n_33), .B(n_148), .Y(n_169) );
OR2x6_ASAP7_75t_L g111 ( .A(n_34), .B(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_35), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_36), .B(n_143), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_37), .A2(n_172), .B1(n_178), .B2(n_182), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_38), .B(n_187), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_40), .A2(n_84), .B1(n_153), .B2(n_508), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_41), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_42), .B(n_214), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_43), .B(n_189), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_44), .B(n_163), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_45), .Y(n_181) );
AND2x2_ASAP7_75t_L g521 ( .A(n_46), .B(n_137), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_47), .B(n_137), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_49), .B(n_163), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_50), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_50), .A2(n_63), .B1(n_428), .B2(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_51), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g146 ( .A(n_52), .Y(n_146) );
INVx1_ASAP7_75t_L g165 ( .A(n_52), .Y(n_165) );
AOI22x1_ASAP7_75t_L g118 ( .A1(n_53), .A2(n_119), .B1(n_120), .B2(n_121), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_53), .Y(n_119) );
AND2x2_ASAP7_75t_L g281 ( .A(n_54), .B(n_137), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g237 ( .A1(n_55), .A2(n_77), .B1(n_143), .B2(n_153), .C(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_56), .B(n_143), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_57), .B(n_520), .Y(n_530) );
INVx1_ASAP7_75t_L g808 ( .A(n_58), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_59), .B(n_172), .Y(n_258) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_60), .A2(n_153), .B(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g558 ( .A(n_61), .B(n_137), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_62), .B(n_217), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_63), .Y(n_820) );
INVx1_ASAP7_75t_L g208 ( .A(n_64), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_65), .B(n_214), .Y(n_556) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_66), .B(n_138), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_67), .A2(n_508), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g279 ( .A(n_68), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_69), .B(n_217), .Y(n_543) );
AND2x2_ASAP7_75t_SL g550 ( .A(n_70), .B(n_189), .Y(n_550) );
XOR2xp5_ASAP7_75t_L g117 ( .A(n_71), .B(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_72), .A2(n_103), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_72), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_73), .A2(n_153), .B(n_278), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_74), .A2(n_818), .B1(n_819), .B2(n_821), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_74), .Y(n_818) );
INVx1_ASAP7_75t_L g151 ( .A(n_75), .Y(n_151) );
INVx1_ASAP7_75t_L g167 ( .A(n_75), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_76), .B(n_143), .Y(n_233) );
AND2x2_ASAP7_75t_L g170 ( .A(n_78), .B(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g209 ( .A(n_79), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_80), .A2(n_153), .B(n_159), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_81), .A2(n_153), .B(n_184), .C(n_188), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_82), .A2(n_87), .B1(n_143), .B2(n_520), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_83), .B(n_520), .Y(n_557) );
INVx1_ASAP7_75t_L g114 ( .A(n_85), .Y(n_114) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_86), .B(n_171), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_88), .A2(n_153), .B1(n_228), .B2(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_89), .B(n_214), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_90), .B(n_214), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_91), .A2(n_508), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g196 ( .A(n_93), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_94), .B(n_217), .Y(n_555) );
AND2x2_ASAP7_75t_L g234 ( .A(n_95), .B(n_171), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_96), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
INVxp67_ASAP7_75t_L g507 ( .A(n_97), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_98), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_99), .B(n_217), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_100), .A2(n_508), .B(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g795 ( .A(n_101), .Y(n_795) );
BUFx2_ASAP7_75t_SL g802 ( .A(n_101), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_102), .B(n_163), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_103), .Y(n_123) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_115), .Y(n_106) );
INVx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x6_ASAP7_75t_SL g492 ( .A(n_110), .B(n_111), .Y(n_492) );
OR2x6_ASAP7_75t_SL g783 ( .A(n_110), .B(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_110), .B(n_784), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_111), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B1(n_124), .B2(n_785), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_491), .B1(n_493), .B2(n_781), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_126), .A2(n_491), .B1(n_494), .B2(n_786), .Y(n_785) );
AND3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_485), .C(n_488), .Y(n_126) );
NAND5xp2_ASAP7_75t_L g127 ( .A(n_128), .B(n_385), .C(n_415), .D(n_429), .E(n_455), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_129), .A2(n_428), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g814 ( .A(n_129), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_334), .Y(n_129) );
NOR3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_282), .C(n_316), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_199), .B(n_221), .C(n_260), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_174), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_134), .B(n_272), .Y(n_337) );
AND2x2_ASAP7_75t_L g424 ( .A(n_134), .B(n_202), .Y(n_424) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g220 ( .A(n_135), .B(n_191), .Y(n_220) );
INVx1_ASAP7_75t_L g262 ( .A(n_135), .Y(n_262) );
INVx2_ASAP7_75t_L g267 ( .A(n_135), .Y(n_267) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_135), .Y(n_295) );
INVx1_ASAP7_75t_L g309 ( .A(n_135), .Y(n_309) );
AND2x2_ASAP7_75t_L g313 ( .A(n_135), .B(n_204), .Y(n_313) );
AND2x2_ASAP7_75t_L g394 ( .A(n_135), .B(n_203), .Y(n_394) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .B(n_170), .Y(n_135) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_136), .A2(n_525), .B(n_531), .Y(n_524) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_136), .A2(n_552), .B(n_558), .Y(n_551) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_136), .A2(n_525), .B(n_531), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_137), .Y(n_136) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_137), .A2(n_582), .B(n_586), .Y(n_581) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g182 ( .A(n_139), .B(n_140), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_152), .Y(n_141) );
INVx1_ASAP7_75t_L g259 ( .A(n_143), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_143), .A2(n_153), .B1(n_501), .B2(n_503), .Y(n_500) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
OR2x6_ASAP7_75t_L g161 ( .A(n_145), .B(n_157), .Y(n_161) );
INVxp33_ASAP7_75t_L g231 ( .A(n_145), .Y(n_231) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g158 ( .A(n_146), .B(n_148), .Y(n_158) );
AND2x4_ASAP7_75t_L g217 ( .A(n_146), .B(n_166), .Y(n_217) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g508 ( .A(n_150), .B(n_158), .Y(n_508) );
INVx2_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
AND2x6_ASAP7_75t_L g214 ( .A(n_151), .B(n_164), .Y(n_214) );
INVxp67_ASAP7_75t_L g257 ( .A(n_153), .Y(n_257) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_158), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g232 ( .A(n_156), .Y(n_232) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g159 ( .A1(n_160), .A2(n_161), .B(n_162), .C(n_168), .Y(n_159) );
INVx2_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_168), .B(n_196), .C(n_197), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_161), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_161), .A2(n_168), .B(n_239), .C(n_240), .Y(n_238) );
INVxp67_ASAP7_75t_L g247 ( .A(n_161), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_161), .A2(n_168), .B(n_279), .C(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
AND2x4_ASAP7_75t_L g520 ( .A(n_163), .B(n_169), .Y(n_520) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_166), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_168), .A2(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_168), .B(n_182), .Y(n_218) );
INVx1_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_168), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_168), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_168), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_168), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_168), .A2(n_576), .B(n_577), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_168), .A2(n_584), .B(n_585), .Y(n_583) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_171), .A2(n_246), .B1(n_251), .B2(n_252), .Y(n_245) );
INVx3_ASAP7_75t_L g252 ( .A(n_171), .Y(n_252) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_172), .B(n_255), .Y(n_254) );
AOI21x1_ASAP7_75t_L g513 ( .A1(n_172), .A2(n_514), .B(n_521), .Y(n_513) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_173), .Y(n_189) );
AND2x4_ASAP7_75t_SL g174 ( .A(n_175), .B(n_190), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g219 ( .A(n_176), .Y(n_219) );
AND2x2_ASAP7_75t_L g263 ( .A(n_176), .B(n_204), .Y(n_263) );
AND2x2_ASAP7_75t_L g284 ( .A(n_176), .B(n_191), .Y(n_284) );
INVx1_ASAP7_75t_L g307 ( .A(n_176), .Y(n_307) );
AND2x4_ASAP7_75t_L g374 ( .A(n_176), .B(n_203), .Y(n_374) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_183), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .C(n_181), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_182), .A2(n_194), .B(n_198), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_182), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_182), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_182), .B(n_507), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_182), .B(n_210), .C(n_510), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_182), .A2(n_539), .B(n_540), .Y(n_538) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_188), .A2(n_226), .B(n_234), .Y(n_225) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_188), .A2(n_226), .B(n_234), .Y(n_289) );
AOI21x1_ASAP7_75t_L g546 ( .A1(n_188), .A2(n_547), .B(n_550), .Y(n_546) );
INVx2_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_189), .A2(n_237), .B(n_241), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_189), .A2(n_573), .B(n_574), .Y(n_572) );
AND2x4_ASAP7_75t_L g390 ( .A(n_190), .B(n_307), .Y(n_390) );
OR2x2_ASAP7_75t_L g431 ( .A(n_190), .B(n_432), .Y(n_431) );
NOR2xp67_ASAP7_75t_SL g450 ( .A(n_190), .B(n_323), .Y(n_450) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_190), .B(n_382), .Y(n_468) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2x1_ASAP7_75t_SL g268 ( .A(n_191), .B(n_204), .Y(n_268) );
AND2x4_ASAP7_75t_L g306 ( .A(n_191), .B(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_191), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_191), .B(n_266), .Y(n_344) );
INVx2_ASAP7_75t_L g358 ( .A(n_191), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_191), .B(n_310), .Y(n_380) );
AND2x2_ASAP7_75t_L g472 ( .A(n_191), .B(n_330), .Y(n_472) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2x1_ASAP7_75t_L g200 ( .A(n_201), .B(n_220), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_202), .B(n_309), .Y(n_323) );
AND2x2_ASAP7_75t_SL g332 ( .A(n_202), .B(n_312), .Y(n_332) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_219), .Y(n_202) );
INVx1_ASAP7_75t_L g310 ( .A(n_203), .Y(n_310) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g330 ( .A(n_204), .Y(n_330) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_211), .B(n_218), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_210), .B(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B1(n_215), .B2(n_216), .Y(n_211) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g363 ( .A(n_219), .Y(n_363) );
INVx2_ASAP7_75t_SL g408 ( .A(n_220), .Y(n_408) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_242), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_223), .B(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g354 ( .A(n_223), .Y(n_354) );
AND2x2_ASAP7_75t_L g478 ( .A(n_223), .B(n_303), .Y(n_478) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_235), .Y(n_223) );
AND2x4_ASAP7_75t_L g291 ( .A(n_224), .B(n_273), .Y(n_291) );
INVx1_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
AND2x2_ASAP7_75t_L g333 ( .A(n_224), .B(n_288), .Y(n_333) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_225), .B(n_236), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_225), .B(n_274), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_227), .B(n_233), .Y(n_226) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVxp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g271 ( .A(n_236), .Y(n_271) );
AND2x4_ASAP7_75t_L g339 ( .A(n_236), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g351 ( .A(n_236), .Y(n_351) );
INVx1_ASAP7_75t_L g393 ( .A(n_236), .Y(n_393) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_236), .Y(n_405) );
AND2x2_ASAP7_75t_L g421 ( .A(n_236), .B(n_244), .Y(n_421) );
BUFx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g368 ( .A(n_243), .B(n_326), .Y(n_368) );
INVx1_ASAP7_75t_SL g370 ( .A(n_243), .Y(n_370) );
AND2x2_ASAP7_75t_L g391 ( .A(n_243), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x4_ASAP7_75t_L g270 ( .A(n_244), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g298 ( .A(n_244), .Y(n_298) );
INVx2_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_244), .B(n_274), .Y(n_319) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_253), .Y(n_244) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_275), .B(n_281), .Y(n_274) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_252), .A2(n_275), .B(n_281), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_257), .B1(n_258), .B2(n_259), .Y(n_253) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B(n_269), .Y(n_260) );
INVx1_ASAP7_75t_L g400 ( .A(n_261), .Y(n_400) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g320 ( .A(n_263), .Y(n_320) );
AND2x2_ASAP7_75t_L g376 ( .A(n_263), .B(n_312), .Y(n_376) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_265), .B(n_306), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_265), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g397 ( .A(n_265), .B(n_390), .Y(n_397) );
AND2x2_ASAP7_75t_L g471 ( .A(n_265), .B(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_266), .Y(n_459) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_267), .Y(n_379) );
AND2x2_ASAP7_75t_L g292 ( .A(n_268), .B(n_293), .Y(n_292) );
OAI21xp33_ASAP7_75t_L g480 ( .A1(n_268), .A2(n_481), .B(n_483), .Y(n_480) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx3_ASAP7_75t_L g366 ( .A(n_270), .Y(n_366) );
NAND2x1_ASAP7_75t_SL g410 ( .A(n_270), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g413 ( .A(n_270), .B(n_291), .Y(n_413) );
AND2x2_ASAP7_75t_L g325 ( .A(n_272), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g462 ( .A(n_272), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g473 ( .A(n_272), .B(n_421), .Y(n_473) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_273), .B(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g404 ( .A(n_274), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_296), .B(n_299), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_291), .B2(n_292), .Y(n_283) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_290), .Y(n_285) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g420 ( .A(n_286), .B(n_421), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_286), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_286), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_288), .B(n_304), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_288), .B(n_304), .Y(n_384) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_288), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g340 ( .A(n_289), .Y(n_340) );
AND2x2_ASAP7_75t_L g348 ( .A(n_289), .B(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g411 ( .A(n_289), .Y(n_411) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_294), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g441 ( .A(n_297), .B(n_326), .Y(n_441) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
AND2x2_ASAP7_75t_L g338 ( .A(n_298), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g426 ( .A(n_298), .B(n_333), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_305), .B1(n_311), .B2(n_314), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g434 ( .A(n_301), .B(n_435), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g464 ( .A(n_304), .B(n_351), .Y(n_464) );
AND2x2_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx2_ASAP7_75t_L g331 ( .A(n_306), .Y(n_331) );
OAI21xp33_ASAP7_75t_SL g477 ( .A1(n_306), .A2(n_478), .B(n_479), .Y(n_477) );
AND2x4_ASAP7_75t_SL g308 ( .A(n_309), .B(n_310), .Y(n_308) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_309), .Y(n_467) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_SL g409 ( .A1(n_312), .A2(n_410), .B(n_412), .C(n_414), .Y(n_409) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_313), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g414 ( .A(n_313), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_313), .B(n_390), .Y(n_454) );
INVx1_ASAP7_75t_SL g321 ( .A(n_314), .Y(n_321) );
AND2x2_ASAP7_75t_L g402 ( .A(n_315), .B(n_339), .Y(n_402) );
INVx1_ASAP7_75t_L g447 ( .A(n_315), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B1(n_321), .B2(n_322), .C(n_324), .Y(n_316) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_317), .Y(n_436) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g484 ( .A(n_319), .B(n_327), .Y(n_484) );
OR2x2_ASAP7_75t_L g343 ( .A(n_320), .B(n_344), .Y(n_343) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_320), .B(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_320), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g482 ( .A(n_320), .B(n_379), .Y(n_482) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI32xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .A3(n_331), .B1(n_332), .B2(n_333), .Y(n_324) );
INVx1_ASAP7_75t_L g345 ( .A(n_326), .Y(n_345) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_328), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g440 ( .A(n_329), .Y(n_440) );
OAI22xp33_ASAP7_75t_SL g422 ( .A1(n_331), .A2(n_423), .B1(n_425), .B2(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g453 ( .A(n_332), .Y(n_453) );
AOI211x1_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_341), .B(n_342), .C(n_359), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_336), .B(n_421), .Y(n_427) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g383 ( .A(n_339), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g449 ( .A(n_339), .Y(n_449) );
OAI222xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B1(n_346), .B2(n_352), .C1(n_353), .C2(n_355), .Y(n_342) );
INVxp67_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_347), .B(n_432), .Y(n_479) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g395 ( .A(n_348), .B(n_392), .Y(n_395) );
INVx3_ASAP7_75t_L g435 ( .A(n_350), .Y(n_435) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g373 ( .A(n_358), .B(n_374), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B1(n_367), .B2(n_372), .C(n_375), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_361), .A2(n_418), .B(n_420), .Y(n_417) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g371 ( .A(n_365), .Y(n_371) );
OR2x2_ASAP7_75t_L g475 ( .A(n_366), .B(n_411), .Y(n_475) );
NOR2xp67_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_369), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_372), .A2(n_401), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_373), .A2(n_445), .B(n_452), .Y(n_451) );
INVx4_ASAP7_75t_L g382 ( .A(n_374), .Y(n_382) );
OAI31xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .A3(n_381), .B(n_383), .Y(n_375) );
INVx1_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_398), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_386), .B(n_398), .C(n_417), .D(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_396), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_391), .B1(n_394), .B2(n_395), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g458 ( .A(n_390), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_391), .B(n_411), .Y(n_419) );
INVx1_ASAP7_75t_SL g432 ( .A(n_394), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_409), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_403), .B2(n_406), .Y(n_399) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_408), .A2(n_471), .B1(n_473), .B2(n_474), .Y(n_470) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_422), .C(n_428), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g487 ( .A(n_422), .Y(n_487) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_428), .A2(n_489), .B(n_490), .Y(n_488) );
INVxp33_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
AND2x2_ASAP7_75t_L g813 ( .A(n_429), .B(n_455), .Y(n_813) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_430), .B(n_437), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_434), .B2(n_436), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_434), .A2(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g444 ( .A(n_435), .Y(n_444) );
NAND3xp33_ASAP7_75t_SL g437 ( .A(n_438), .B(n_442), .C(n_451), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_445), .B1(n_448), .B2(n_450), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVxp33_ASAP7_75t_SL g490 ( .A(n_455), .Y(n_490) );
NOR3x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_469), .C(n_476), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_477), .B(n_480), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g815 ( .A(n_486), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_658), .Y(n_494) );
NOR4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_601), .C(n_640), .D(n_647), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_522), .B1(n_559), .B2(n_568), .C(n_587), .Y(n_496) );
OR2x2_ASAP7_75t_L g731 ( .A(n_497), .B(n_593), .Y(n_731) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g646 ( .A(n_498), .B(n_571), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_498), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_498), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_511), .Y(n_498) );
AND2x4_ASAP7_75t_SL g570 ( .A(n_499), .B(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g592 ( .A(n_499), .Y(n_592) );
AND2x2_ASAP7_75t_L g627 ( .A(n_499), .B(n_600), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_499), .B(n_512), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_499), .B(n_594), .Y(n_679) );
OR2x2_ASAP7_75t_L g757 ( .A(n_499), .B(n_571), .Y(n_757) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .Y(n_499) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g579 ( .A(n_512), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_512), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g605 ( .A(n_512), .Y(n_605) );
OR2x2_ASAP7_75t_L g610 ( .A(n_512), .B(n_594), .Y(n_610) );
AND2x2_ASAP7_75t_L g623 ( .A(n_512), .B(n_581), .Y(n_623) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_512), .Y(n_626) );
INVx1_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_512), .B(n_592), .Y(n_703) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_532), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g567 ( .A(n_524), .B(n_551), .Y(n_567) );
AND2x4_ASAP7_75t_L g597 ( .A(n_524), .B(n_536), .Y(n_597) );
INVx2_ASAP7_75t_L g631 ( .A(n_524), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_524), .B(n_551), .Y(n_689) );
AND2x2_ASAP7_75t_L g736 ( .A(n_524), .B(n_565), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
AOI222xp33_ASAP7_75t_L g724 ( .A1(n_532), .A2(n_596), .B1(n_639), .B2(n_699), .C1(n_725), .C2(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_544), .Y(n_533) );
AND2x2_ASAP7_75t_L g643 ( .A(n_534), .B(n_563), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_534), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g772 ( .A(n_534), .B(n_612), .Y(n_772) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_535), .A2(n_603), .B(n_607), .Y(n_602) );
AND2x2_ASAP7_75t_L g683 ( .A(n_535), .B(n_566), .Y(n_683) );
OR2x2_ASAP7_75t_L g708 ( .A(n_535), .B(n_567), .Y(n_708) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx5_ASAP7_75t_L g562 ( .A(n_536), .Y(n_562) );
AND2x2_ASAP7_75t_L g649 ( .A(n_536), .B(n_631), .Y(n_649) );
AND2x2_ASAP7_75t_L g675 ( .A(n_536), .B(n_551), .Y(n_675) );
OR2x2_ASAP7_75t_L g678 ( .A(n_536), .B(n_565), .Y(n_678) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_536), .Y(n_696) );
AND2x4_ASAP7_75t_SL g753 ( .A(n_536), .B(n_630), .Y(n_753) );
OR2x2_ASAP7_75t_L g762 ( .A(n_536), .B(n_589), .Y(n_762) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
AOI221xp5_ASAP7_75t_SL g713 ( .A1(n_544), .A2(n_597), .B1(n_714), .B2(n_716), .C(n_717), .Y(n_713) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_551), .Y(n_544) );
OR2x2_ASAP7_75t_L g652 ( .A(n_545), .B(n_622), .Y(n_652) );
OR2x2_ASAP7_75t_L g662 ( .A(n_545), .B(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g688 ( .A(n_545), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g694 ( .A(n_545), .B(n_613), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_545), .B(n_677), .Y(n_706) );
INVx2_ASAP7_75t_L g719 ( .A(n_545), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_545), .B(n_597), .Y(n_740) );
AND2x2_ASAP7_75t_L g744 ( .A(n_545), .B(n_566), .Y(n_744) );
AND2x2_ASAP7_75t_L g752 ( .A(n_545), .B(n_753), .Y(n_752) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g565 ( .A(n_546), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_551), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g596 ( .A(n_551), .B(n_565), .Y(n_596) );
INVx2_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
AND2x4_ASAP7_75t_L g630 ( .A(n_551), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_551), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g742 ( .A(n_561), .B(n_564), .Y(n_742) );
AND2x4_ASAP7_75t_L g588 ( .A(n_562), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g629 ( .A(n_562), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g656 ( .A(n_562), .B(n_596), .Y(n_656) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
AND2x2_ASAP7_75t_L g760 ( .A(n_564), .B(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g612 ( .A(n_565), .B(n_613), .Y(n_612) );
OAI21xp5_ASAP7_75t_SL g632 ( .A1(n_566), .A2(n_633), .B(n_639), .Y(n_632) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_579), .Y(n_569) );
INVx1_ASAP7_75t_SL g686 ( .A(n_570), .Y(n_686) );
AND2x2_ASAP7_75t_L g716 ( .A(n_570), .B(n_626), .Y(n_716) );
AND2x4_ASAP7_75t_L g727 ( .A(n_570), .B(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g593 ( .A(n_571), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g600 ( .A(n_571), .Y(n_600) );
AND2x4_ASAP7_75t_L g606 ( .A(n_571), .B(n_592), .Y(n_606) );
INVx2_ASAP7_75t_L g617 ( .A(n_571), .Y(n_617) );
INVx1_ASAP7_75t_L g666 ( .A(n_571), .Y(n_666) );
OR2x2_ASAP7_75t_L g687 ( .A(n_571), .B(n_671), .Y(n_687) );
OR2x2_ASAP7_75t_L g701 ( .A(n_571), .B(n_581), .Y(n_701) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_571), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_571), .B(n_623), .Y(n_773) );
OR2x6_ASAP7_75t_L g571 ( .A(n_572), .B(n_578), .Y(n_571) );
INVx1_ASAP7_75t_L g618 ( .A(n_579), .Y(n_618) );
AND2x2_ASAP7_75t_L g751 ( .A(n_579), .B(n_617), .Y(n_751) );
AND2x2_ASAP7_75t_L g776 ( .A(n_579), .B(n_606), .Y(n_776) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g594 ( .A(n_581), .Y(n_594) );
BUFx3_ASAP7_75t_L g636 ( .A(n_581), .Y(n_636) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_581), .Y(n_663) );
INVx1_ASAP7_75t_L g672 ( .A(n_581), .Y(n_672) );
AOI33xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_590), .A3(n_595), .B1(n_596), .B2(n_597), .B3(n_598), .Y(n_587) );
AOI21x1_ASAP7_75t_SL g690 ( .A1(n_588), .A2(n_612), .B(n_674), .Y(n_690) );
INVx2_ASAP7_75t_L g720 ( .A(n_588), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_588), .B(n_719), .Y(n_726) );
AND2x2_ASAP7_75t_L g674 ( .A(n_589), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g637 ( .A(n_592), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g738 ( .A(n_593), .Y(n_738) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_594), .Y(n_728) );
OAI32xp33_ASAP7_75t_L g777 ( .A1(n_595), .A2(n_597), .A3(n_773), .B1(n_778), .B2(n_780), .Y(n_777) );
AND2x2_ASAP7_75t_L g695 ( .A(n_596), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_SL g685 ( .A(n_597), .Y(n_685) );
AND2x2_ASAP7_75t_L g750 ( .A(n_597), .B(n_694), .Y(n_750) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_611), .B1(n_614), .B2(n_628), .C(n_632), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_605), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_606), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_606), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_606), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g655 ( .A(n_610), .Y(n_655) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .C(n_624), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_616), .A2(n_678), .B1(n_718), .B2(n_721), .Y(n_717) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g621 ( .A(n_617), .Y(n_621) );
NOR2x1p5_ASAP7_75t_L g635 ( .A(n_617), .B(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI322xp33_ASAP7_75t_L g684 ( .A1(n_620), .A2(n_662), .A3(n_685), .B1(n_686), .B2(n_687), .C1(n_688), .C2(n_690), .Y(n_684) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_622), .A2(n_641), .B(n_642), .C(n_644), .Y(n_640) );
OR2x2_ASAP7_75t_L g732 ( .A(n_622), .B(n_686), .Y(n_732) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g639 ( .A(n_623), .B(n_627), .Y(n_639) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g645 ( .A(n_629), .B(n_646), .Y(n_645) );
INVx3_ASAP7_75t_SL g677 ( .A(n_630), .Y(n_677) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_634), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_SL g681 ( .A(n_637), .Y(n_681) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_638), .Y(n_723) );
OR2x6_ASAP7_75t_SL g778 ( .A(n_641), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI211xp5_ASAP7_75t_L g768 ( .A1(n_646), .A2(n_769), .B(n_770), .C(n_777), .Y(n_768) );
O2A1O1Ixp33_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_650), .B(n_653), .C(n_657), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_648), .A2(n_660), .B(n_667), .C(n_691), .Y(n_659) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_704), .C(n_748), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_663), .Y(n_755) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g710 ( .A(n_666), .Y(n_710) );
NOR3xp33_ASAP7_75t_SL g667 ( .A(n_668), .B(n_680), .C(n_684), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_673), .B1(n_676), .B2(n_679), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g712 ( .A(n_672), .Y(n_712) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_672), .Y(n_779) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_SL g765 ( .A(n_678), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
OR2x2_ASAP7_75t_L g715 ( .A(n_681), .B(n_701), .Y(n_715) );
OR2x2_ASAP7_75t_L g766 ( .A(n_681), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g764 ( .A(n_689), .Y(n_764) );
OR2x2_ASAP7_75t_L g780 ( .A(n_689), .B(n_719), .Y(n_780) );
OAI21xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B(n_697), .Y(n_691) );
OAI31xp33_ASAP7_75t_L g705 ( .A1(n_692), .A2(n_706), .A3(n_707), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g737 ( .A(n_702), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND4xp25_ASAP7_75t_SL g704 ( .A(n_705), .B(n_713), .C(n_724), .D(n_729), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_712), .Y(n_747) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_733), .B1(n_737), .B2(n_739), .C(n_741), .Y(n_729) );
NAND2xp33_ASAP7_75t_SL g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g774 ( .A(n_733), .Y(n_774) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g769 ( .A(n_743), .Y(n_769) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_749), .B(n_768), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B1(n_752), .B2(n_754), .C(n_758), .Y(n_749) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_763), .B(n_766), .Y(n_758) );
INVxp33_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_773), .B1(n_774), .B2(n_775), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_782), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_796), .Y(n_789) );
INVxp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_792), .B(n_795), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_793), .A2(n_800), .B(n_803), .Y(n_799) );
OR2x2_ASAP7_75t_SL g831 ( .A(n_793), .B(n_795), .Y(n_831) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_L g804 ( .A(n_797), .Y(n_804) );
BUFx3_ASAP7_75t_L g825 ( .A(n_797), .Y(n_825) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
CKINVDCx11_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
CKINVDCx8_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_826), .B(n_829), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_810), .B(n_822), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_807), .A2(n_823), .B(n_824), .Y(n_822) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g823 ( .A(n_811), .Y(n_823) );
XNOR2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_816), .Y(n_811) );
NAND3x1_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .C(n_815), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g821 ( .A(n_819), .Y(n_821) );
CKINVDCx11_ASAP7_75t_R g828 ( .A(n_824), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
endmodule