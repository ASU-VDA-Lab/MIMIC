module real_aes_8915_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_34;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_9;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
INVx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
OAI221xp5_ASAP7_75t_L g22 ( .A1(n_1), .A2(n_3), .B1(n_7), .B2(n_23), .C(n_24), .Y(n_22) );
INVxp67_ASAP7_75t_L g25 ( .A(n_1), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
INVxp67_ASAP7_75t_L g26 ( .A(n_3), .Y(n_26) );
AND2x6_ASAP7_75t_L g18 ( .A(n_4), .B(n_19), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_4), .B(n_21), .Y(n_20) );
INVx1_ASAP7_75t_L g31 ( .A(n_4), .Y(n_31) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
INVx1_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_SL g8 ( .A1(n_9), .A2(n_20), .B(n_27), .C(n_32), .Y(n_8) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_14), .B(n_18), .Y(n_13) );
OA21x2_ASAP7_75t_L g27 ( .A1(n_14), .A2(n_28), .B(n_30), .Y(n_27) );
AND2x2_ASAP7_75t_L g14 ( .A(n_15), .B(n_17), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_19), .Y(n_29) );
INVxp67_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_25), .B(n_26), .Y(n_24) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_27), .Y(n_34) );
INVx1_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
NAND2xp5_ASAP7_75t_SL g30 ( .A(n_29), .B(n_31), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_31), .B(n_33), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
endmodule