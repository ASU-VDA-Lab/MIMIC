module real_jpeg_17875_n_22 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_100, n_11, n_14, n_7, n_18, n_3, n_99, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_22);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_100;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_99;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_22;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

OAI221xp5_ASAP7_75t_L g23 ( 
.A1(n_2),
.A2(n_11),
.B1(n_24),
.B2(n_29),
.C(n_30),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_17),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_18),
.B(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_6),
.B(n_51),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_6),
.C(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_4),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_7),
.B(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_8),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_8),
.B(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_13),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_25),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_16),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_86),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_62),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_93),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_24),
.A2(n_38),
.B(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_96),
.Y(n_97)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_47),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_68),
.C(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_87),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_39),
.B(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_31),
.A2(n_39),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_95),
.B(n_97),
.Y(n_32)
);

OAI311xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.A3(n_36),
.B1(n_89),
.C1(n_91),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.C(n_42),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_85),
.B(n_88),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_81),
.B(n_84),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_80),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_76),
.B(n_79),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_71),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_65),
.B(n_70),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_61),
.B(n_64),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B(n_69),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_99),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_100),
.Y(n_63)
);


endmodule