module fake_jpeg_3459_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_44),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_45),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_110)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_21),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_28),
.B1(n_32),
.B2(n_30),
.Y(n_96)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_60),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_39),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_4),
.B(n_5),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_73),
.Y(n_106)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_26),
.A2(n_7),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_22),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_76),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_86),
.B(n_93),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_88),
.B(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_91),
.B(n_92),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_37),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_110),
.B1(n_90),
.B2(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_50),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_29),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_107),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_47),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_37),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_41),
.B(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_105),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_36),
.B1(n_48),
.B2(n_59),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_77),
.B1(n_98),
.B2(n_79),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_117),
.B(n_129),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_66),
.B(n_41),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_135),
.B(n_113),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_120),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_46),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_51),
.B1(n_53),
.B2(n_72),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx24_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_134),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_85),
.B(n_104),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_87),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_89),
.B1(n_79),
.B2(n_90),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_132),
.B1(n_118),
.B2(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_95),
.B1(n_103),
.B2(n_112),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_104),
.C(n_85),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_119),
.C(n_134),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_149),
.Y(n_152)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_146),
.Y(n_153)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

CKINVDCx12_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_150),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_105),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_167),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_140),
.B1(n_127),
.B2(n_139),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_128),
.Y(n_164)
);

XNOR2x2_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_120),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_168),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_133),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_164),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_144),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_174),
.C(n_155),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_170),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_141),
.B(n_150),
.C(n_159),
.D(n_166),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_172),
.B1(n_162),
.B2(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_168),
.B1(n_152),
.B2(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_175),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_152),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_186),
.C(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_209),
.B1(n_195),
.B2(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_176),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_192),
.C(n_178),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_176),
.B1(n_153),
.B2(n_165),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_173),
.B(n_177),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_207),
.B1(n_204),
.B2(n_198),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_219),
.Y(n_225)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_186),
.C(n_200),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_189),
.B1(n_195),
.B2(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_205),
.B1(n_209),
.B2(n_203),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_223),
.Y(n_233)
);

AOI321xp33_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_201),
.A3(n_184),
.B1(n_198),
.B2(n_202),
.C(n_206),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_197),
.B(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_223),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_156),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_231),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_230),
.A2(n_228),
.B1(n_211),
.B2(n_225),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_184),
.C(n_214),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_180),
.B1(n_215),
.B2(n_213),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_239),
.A3(n_173),
.B1(n_232),
.B2(n_231),
.C1(n_161),
.C2(n_158),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_215),
.B1(n_153),
.B2(n_165),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_158),
.A3(n_161),
.B1(n_233),
.B2(n_221),
.C1(n_234),
.C2(n_201),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_238),
.C(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_244),
.B(n_240),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);


endmodule