module fake_jpeg_16019_n_192 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_37),
.B(n_42),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_23),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_6),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_43),
.B(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_16),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_10),
.B1(n_28),
.B2(n_35),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_28),
.B1(n_34),
.B2(n_31),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_16),
.B(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_17),
.A2(n_29),
.B1(n_21),
.B2(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_95)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_22),
.Y(n_66)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_66),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_85),
.B1(n_88),
.B2(n_67),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_17),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_34),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_85),
.Y(n_96)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_90),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_21),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_82),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_30),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_83),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_32),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_25),
.C(n_38),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_40),
.B1(n_65),
.B2(n_23),
.Y(n_121)
);

NAND2x1_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_44),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_104),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_77),
.B(n_68),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_107),
.B(n_108),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_121),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_84),
.B1(n_62),
.B2(n_75),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_106),
.B1(n_111),
.B2(n_114),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_65),
.B1(n_76),
.B2(n_87),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_63),
.B(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_89),
.B1(n_75),
.B2(n_70),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_82),
.B(n_71),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_68),
.B1(n_73),
.B2(n_80),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_79),
.B1(n_74),
.B2(n_78),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_61),
.A2(n_86),
.B1(n_77),
.B2(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_78),
.B1(n_82),
.B2(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_96),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_107),
.C(n_101),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_137),
.C(n_133),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_112),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_139),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_100),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_99),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_110),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_105),
.C(n_114),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_156),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_106),
.B1(n_111),
.B2(n_119),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_157),
.B1(n_126),
.B2(n_125),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_131),
.C(n_127),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_141),
.C(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_115),
.B1(n_116),
.B2(n_103),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_134),
.B(n_143),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_142),
.B(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_162),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_143),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_132),
.B1(n_123),
.B2(n_124),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_178),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_147),
.A3(n_156),
.B1(n_146),
.B2(n_153),
.C1(n_115),
.C2(n_145),
.Y(n_177)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_148),
.C(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_160),
.B1(n_164),
.B2(n_159),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_155),
.B(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_168),
.B1(n_163),
.B2(n_126),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_162),
.B(n_165),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_178),
.C(n_169),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_180),
.CI(n_179),
.CON(n_189),
.SN(n_189)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_169),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_185),
.A2(n_183),
.B(n_174),
.C(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_175),
.B1(n_186),
.B2(n_187),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_175),
.C(n_172),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_191),
.Y(n_192)
);


endmodule