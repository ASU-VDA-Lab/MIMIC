module fake_jpeg_24019_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_18),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_44),
.CON(n_61),
.SN(n_61)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_1),
.C(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_63),
.B1(n_69),
.B2(n_19),
.Y(n_90)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_64),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_22),
.B1(n_28),
.B2(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_32),
.B1(n_22),
.B2(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_76),
.Y(n_103)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_78),
.Y(n_111)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_49),
.Y(n_101)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_43),
.B1(n_37),
.B2(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_87),
.B1(n_57),
.B2(n_62),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_89),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_43),
.B1(n_37),
.B2(n_40),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_40),
.B(n_44),
.C(n_45),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_90),
.B1(n_98),
.B2(n_20),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_48),
.B1(n_47),
.B2(n_34),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_50),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_48),
.C(n_49),
.Y(n_104)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_52),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_106),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_73),
.B(n_83),
.Y(n_124)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_109),
.B1(n_93),
.B2(n_47),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_57),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_56),
.B1(n_45),
.B2(n_62),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_79),
.B(n_82),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_29),
.B1(n_26),
.B2(n_18),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_23),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_114),
.A2(n_94),
.B(n_47),
.C(n_33),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_74),
.B(n_15),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_15),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_75),
.Y(n_136)
);

NOR4xp25_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_77),
.C(n_87),
.D(n_85),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_125),
.B(n_114),
.C(n_119),
.D(n_106),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_140),
.B(n_118),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_82),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_94),
.C(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_138),
.Y(n_149)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_78),
.B1(n_84),
.B2(n_81),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_137),
.B1(n_142),
.B2(n_143),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_95),
.B1(n_70),
.B2(n_34),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_141),
.B1(n_105),
.B2(n_115),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_2),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_33),
.B1(n_29),
.B2(n_26),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_33),
.B1(n_29),
.B2(n_26),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_110),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_148),
.C(n_153),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_111),
.B(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_120),
.C(n_102),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_114),
.B(n_107),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_157),
.B1(n_123),
.B2(n_8),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_126),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_143),
.B1(n_126),
.B2(n_131),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_158),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_159),
.C(n_150),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_102),
.B1(n_115),
.B2(n_121),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_117),
.C(n_99),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_2),
.B(n_3),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_6),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_153),
.B(n_151),
.C(n_156),
.D(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_164),
.C(n_173),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_129),
.B(n_140),
.C(n_143),
.D(n_128),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_161),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_165),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_146),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_145),
.C(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_146),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_166),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_152),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_164),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_172),
.B(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_163),
.C(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_181),
.C(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_9),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_190),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_194),
.B(n_184),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_10),
.B(n_12),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_199),
.B(n_12),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_12),
.Y(n_202)
);


endmodule