module fake_aes_12153_n_17 (n_1, n_2, n_4, n_3, n_0, n_17);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
CKINVDCx20_ASAP7_75t_R g5 ( .A(n_1), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
BUFx6f_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
INVxp67_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_9), .B(n_5), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
AOI22xp33_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_11), .Y(n_13) );
INVx3_ASAP7_75t_SL g14 ( .A(n_13), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_13), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
OAI22xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_14), .B1(n_15), .B2(n_12), .Y(n_17) );
endmodule