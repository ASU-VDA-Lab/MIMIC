module fake_jpeg_207_n_518 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_518);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_518;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_58),
.B(n_60),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_0),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_0),
.C(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_65),
.Y(n_104)
);

NAND2x1_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_96),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_1),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_92),
.Y(n_100)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g125 ( 
.A(n_69),
.Y(n_125)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_2),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_19),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_84),
.Y(n_115)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_2),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_28),
.B(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_28),
.B(n_3),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_99),
.B(n_116),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_47),
.B1(n_30),
.B2(n_48),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_103),
.A2(n_113),
.B1(n_119),
.B2(n_123),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_85),
.B1(n_73),
.B2(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_108),
.A2(n_121),
.B1(n_14),
.B2(n_15),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_31),
.B1(n_48),
.B2(n_42),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_31),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_56),
.A2(n_48),
.B1(n_44),
.B2(n_42),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_44),
.B1(n_33),
.B2(n_32),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_141),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_19),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_132),
.B(n_136),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_74),
.A2(n_27),
.B1(n_29),
.B2(n_94),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_133),
.A2(n_135),
.B1(n_140),
.B2(n_110),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_95),
.A2(n_27),
.B1(n_26),
.B2(n_6),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_55),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_26),
.B1(n_5),
.B2(n_8),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_57),
.B(n_59),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_145),
.B(n_125),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_5),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_159),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_5),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_153),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_71),
.B(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_10),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_9),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_129),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_160),
.B(n_197),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_172),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_98),
.B1(n_96),
.B2(n_87),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_120),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_80),
.B1(n_72),
.B2(n_77),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_99),
.A2(n_26),
.B1(n_11),
.B2(n_12),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_169),
.B(n_183),
.Y(n_230)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_101),
.B(n_11),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_173),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_174),
.B(n_204),
.Y(n_257)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_176),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_107),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_104),
.B(n_11),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_178),
.B(n_182),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_101),
.A2(n_26),
.B(n_12),
.C(n_13),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_179),
.A2(n_180),
.B(n_196),
.C(n_183),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_101),
.A2(n_11),
.B(n_12),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_187),
.C(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_13),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_13),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_14),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_194),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_126),
.B(n_14),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_189),
.A2(n_216),
.B1(n_144),
.B2(n_137),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_106),
.B(n_17),
.C(n_15),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_15),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_113),
.A2(n_16),
.B1(n_131),
.B2(n_124),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_195),
.A2(n_215),
.B1(n_209),
.B2(n_160),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_16),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_196),
.Y(n_256)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_130),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_106),
.B(n_118),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_207),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_152),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_201),
.B(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_118),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_130),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_125),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_125),
.B(n_138),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_210),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_102),
.B(n_112),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx4_ASAP7_75t_SL g214 ( 
.A(n_137),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_218),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_131),
.A2(n_143),
.B1(n_124),
.B2(n_128),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_110),
.A2(n_151),
.B1(n_157),
.B2(n_148),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_225),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_239),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_164),
.B(n_112),
.C(n_122),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_186),
.C(n_191),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_151),
.B1(n_109),
.B2(n_128),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_235),
.A2(n_241),
.B(n_264),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_179),
.A2(n_129),
.B(n_157),
.C(n_144),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_237),
.A2(n_184),
.B(n_170),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_174),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_178),
.A2(n_150),
.B(n_137),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_109),
.B1(n_120),
.B2(n_139),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_245),
.A2(n_266),
.B1(n_217),
.B2(n_176),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_195),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_207),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_175),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_206),
.A2(n_143),
.B1(n_139),
.B2(n_146),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g299 ( 
.A1(n_253),
.A2(n_219),
.B(n_245),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_164),
.A2(n_146),
.B1(n_155),
.B2(n_144),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_203),
.B1(n_214),
.B2(n_210),
.Y(n_273)
);

OR2x2_ASAP7_75t_SL g264 ( 
.A(n_208),
.B(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_267),
.B(n_264),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_203),
.A2(n_196),
.B1(n_188),
.B2(n_181),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_194),
.B(n_182),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_211),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_273),
.A2(n_253),
.B1(n_247),
.B2(n_248),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_274),
.A2(n_275),
.B1(n_287),
.B2(n_292),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_185),
.B1(n_169),
.B2(n_200),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_275),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_279),
.B(n_294),
.Y(n_321)
);

INVx11_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_284),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_225),
.B(n_165),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_167),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_286),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_192),
.B(n_198),
.C(n_213),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_229),
.B(n_166),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_289),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_229),
.B(n_218),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_290),
.A2(n_305),
.B(n_307),
.Y(n_319)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_171),
.B1(n_246),
.B2(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_230),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_234),
.A2(n_266),
.B1(n_259),
.B2(n_219),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_295),
.A2(n_299),
.B1(n_315),
.B2(n_318),
.Y(n_354)
);

OR2x4_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_249),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_312),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_233),
.B(n_224),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_230),
.B(n_256),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_228),
.B(n_239),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_301),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_242),
.B(n_261),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_270),
.B(n_242),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_302),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_259),
.A2(n_236),
.B1(n_252),
.B2(n_241),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_221),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_257),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_236),
.A2(n_252),
.B(n_244),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_312),
.A2(n_223),
.B(n_240),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_227),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_316),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_236),
.B(n_257),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_262),
.B(n_223),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_235),
.A2(n_253),
.B1(n_220),
.B2(n_226),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_221),
.B(n_222),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_253),
.A2(n_226),
.B1(n_244),
.B2(n_265),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_271),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_320),
.B(n_346),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_322),
.A2(n_342),
.B(n_344),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_247),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_326),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_325),
.A2(n_274),
.B1(n_308),
.B2(n_311),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_231),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_358),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_231),
.C(n_232),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_347),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_290),
.A2(n_232),
.B(n_238),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_337),
.A2(n_351),
.B(n_286),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_292),
.B(n_296),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_341),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_272),
.Y(n_343)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_305),
.A2(n_240),
.B(n_293),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_271),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_298),
.C(n_307),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_272),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_349),
.B(n_310),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_296),
.A2(n_317),
.B(n_293),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_353),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_314),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_288),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_283),
.B(n_284),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_359),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_300),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_279),
.Y(n_366)
);

AO22x1_ASAP7_75t_SL g362 ( 
.A1(n_341),
.A2(n_318),
.B1(n_315),
.B2(n_295),
.Y(n_362)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_348),
.Y(n_365)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_369),
.B1(n_371),
.B2(n_378),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_354),
.A2(n_299),
.B1(n_286),
.B2(n_287),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_360),
.B1(n_332),
.B2(n_343),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_370),
.B(n_377),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_348),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_373),
.A2(n_375),
.B1(n_384),
.B2(n_387),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_353),
.B(n_319),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_354),
.A2(n_274),
.B1(n_294),
.B2(n_285),
.Y(n_375)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_320),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_383),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_352),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_327),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_382),
.C(n_389),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_SL g404 ( 
.A(n_380),
.B(n_359),
.C(n_332),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_302),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_327),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_334),
.A2(n_304),
.B1(n_281),
.B2(n_299),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_313),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_386),
.B(n_393),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_334),
.A2(n_304),
.B1(n_299),
.B2(n_273),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_SL g388 ( 
.A(n_341),
.B(n_280),
.C(n_291),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_344),
.C(n_351),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_276),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_323),
.B(n_282),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_336),
.C(n_322),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_324),
.B(n_277),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_363),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_340),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_406),
.Y(n_439)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_399),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_381),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_394),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_340),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_408),
.A2(n_413),
.B(n_422),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_381),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_410),
.B(n_321),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_361),
.B(n_352),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_414),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_326),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_417),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_339),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_420),
.C(n_423),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_364),
.B(n_391),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_387),
.A2(n_346),
.B1(n_349),
.B2(n_338),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_418),
.A2(n_368),
.B1(n_378),
.B2(n_365),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_364),
.B(n_385),
.C(n_339),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_392),
.B(n_367),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_341),
.C(n_321),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_422),
.A2(n_353),
.B(n_374),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_432),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_414),
.C(n_417),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_429),
.C(n_430),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_390),
.C(n_371),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_390),
.C(n_372),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_413),
.A2(n_395),
.B(n_319),
.Y(n_432)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_372),
.C(n_383),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_435),
.B(n_423),
.Y(n_455)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_400),
.B1(n_384),
.B2(n_373),
.Y(n_459)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_409),
.Y(n_442)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_335),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_443),
.B(n_424),
.Y(n_460)
);

INVx11_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_444),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_398),
.B(n_375),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_448),
.Y(n_463)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_447),
.B(n_331),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_420),
.B(n_395),
.Y(n_448)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_446),
.B(n_416),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_407),
.Y(n_454)
);

OAI321xp33_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_437),
.A3(n_444),
.B1(n_328),
.B2(n_333),
.C(n_345),
.Y(n_478)
);

OAI221xp5_ASAP7_75t_L g477 ( 
.A1(n_455),
.A2(n_462),
.B1(n_439),
.B2(n_431),
.C(n_425),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_419),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_456),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_400),
.B1(n_418),
.B2(n_412),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_461),
.B1(n_449),
.B2(n_435),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_464),
.B1(n_466),
.B2(n_350),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_399),
.B1(n_325),
.B2(n_337),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_331),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_441),
.A2(n_362),
.B1(n_388),
.B2(n_403),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_426),
.A2(n_362),
.B1(n_356),
.B2(n_304),
.Y(n_466)
);

FAx1_ASAP7_75t_SL g467 ( 
.A(n_440),
.B(n_362),
.CI(n_356),
.CON(n_467),
.SN(n_467)
);

FAx1_ASAP7_75t_SL g472 ( 
.A(n_467),
.B(n_430),
.CI(n_445),
.CON(n_472),
.SN(n_472)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_428),
.B(n_432),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_470),
.B(n_471),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_473),
.C(n_483),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_SL g473 ( 
.A1(n_453),
.A2(n_449),
.B(n_330),
.C(n_448),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_431),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_465),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_446),
.C(n_427),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_467),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_464),
.B(n_454),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_476),
.A2(n_477),
.B(n_303),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_478),
.A2(n_481),
.B1(n_482),
.B2(n_456),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_458),
.A2(n_425),
.B1(n_439),
.B2(n_328),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_463),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_468),
.A2(n_333),
.B1(n_345),
.B2(n_350),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_466),
.A2(n_330),
.B(n_280),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_485),
.B(n_469),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_486),
.B(n_490),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_493),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_482),
.A2(n_456),
.B1(n_467),
.B2(n_459),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_488),
.A2(n_492),
.B1(n_479),
.B2(n_473),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_451),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_463),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_491),
.B(n_494),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_480),
.B(n_451),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_495),
.B(n_472),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_483),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_471),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_500),
.B(n_501),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_474),
.C(n_470),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_489),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_488),
.C(n_481),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_506),
.B(n_507),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_508),
.A2(n_510),
.B(n_473),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_501),
.A2(n_489),
.B(n_473),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_499),
.C(n_505),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_512),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_513),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_511),
.B1(n_498),
.B2(n_472),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_514),
.B(n_330),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_303),
.Y(n_518)
);


endmodule