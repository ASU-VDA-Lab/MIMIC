module real_jpeg_19863_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_269, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_269;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_0),
.A2(n_3),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_42),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_0),
.A2(n_42),
.B1(n_62),
.B2(n_63),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_0),
.A2(n_9),
.B(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_0),
.B(n_52),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_0),
.A2(n_10),
.B(n_63),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_0),
.A2(n_27),
.B(n_28),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_3),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_38),
.B1(n_62),
.B2(n_63),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_3),
.B1(n_37),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_49),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_35),
.B(n_42),
.C(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_4),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_4),
.A2(n_19),
.B1(n_62),
.B2(n_63),
.Y(n_95)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

BUFx3_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_83),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_82),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_65),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_16),
.B(n_65),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_16),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_33),
.CI(n_46),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_18),
.A2(n_24),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_20),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_20),
.A2(n_29),
.B(n_42),
.C(n_208),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_25),
.B(n_28),
.C(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_23),
.B(n_81),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_24),
.A2(n_80),
.B(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_25),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_25),
.A2(n_31),
.B1(n_81),
.B2(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_25),
.B(n_42),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_27),
.A2(n_42),
.B(n_60),
.C(n_185),
.Y(n_184)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_31),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B(n_39),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_37),
.B(n_44),
.C(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_34),
.B(n_43),
.Y(n_97)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_44),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_48),
.B(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_42),
.B(n_93),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_42),
.B(n_61),
.Y(n_191)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.C(n_55),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_113),
.C(n_118),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_47),
.A2(n_68),
.B1(n_106),
.B2(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_47),
.B(n_152),
.C(n_153),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_47),
.A2(n_68),
.B1(n_118),
.B2(n_163),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_55),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_55),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_57),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_58),
.A2(n_61),
.B1(n_64),
.B2(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_61),
.B1(n_104),
.B2(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_62),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_73),
.C(n_75),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.C(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_74),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_73),
.A2(n_74),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_73),
.A2(n_74),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_118),
.C(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_74),
.B(n_240),
.C(n_242),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_127),
.A3(n_131),
.B1(n_265),
.B2(n_266),
.C(n_269),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_119),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_85),
.B(n_119),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_105),
.C(n_111),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_86),
.B(n_105),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_99),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_98),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_88),
.A2(n_89),
.B1(n_100),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_96),
.B(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_91),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_92),
.A2(n_93),
.B1(n_146),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_93),
.A2(n_115),
.B(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_96),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_100),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_110),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_109),
.Y(n_110)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_169),
.C(n_171),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_106),
.A2(n_152),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_121),
.C(n_124),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_111),
.A2(n_112),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_113),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_114),
.A2(n_116),
.B1(n_200),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_114),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_116),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_157),
.C(n_199),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_116),
.A2(n_200),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_116),
.B(n_218),
.C(n_223),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_148),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_118),
.A2(n_138),
.B1(n_139),
.B2(n_163),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_118),
.B(n_139),
.C(n_206),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_128),
.B(n_129),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_259),
.B(n_264),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_247),
.B(n_258),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_175),
.B(n_232),
.C(n_246),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_159),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_135),
.B(n_159),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_150),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_147),
.C(n_150),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_139),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_138),
.B(n_143),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_184),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_191),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_167),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.C(n_168),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_160),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_168),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_231),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_225),
.B(n_230),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_215),
.B(n_224),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_203),
.B(n_214),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_194),
.B(n_202),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_193),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B(n_192),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_212),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_244),
.B2(n_245),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_239),
.C(n_245),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);


endmodule