module real_jpeg_26212_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_72),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_64),
.B1(n_67),
.B2(n_72),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_36),
.B1(n_64),
.B2(n_67),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_4),
.A2(n_36),
.B1(n_59),
.B2(n_169),
.Y(n_349)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_5),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_6),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_6),
.B(n_63),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_6),
.A2(n_67),
.B(n_81),
.C(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_6),
.A2(n_64),
.B1(n_67),
.B2(n_170),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_6),
.B(n_29),
.C(n_45),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_170),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_6),
.A2(n_26),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_6),
.B(n_124),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_61),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_61),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_8),
.A2(n_64),
.B1(n_67),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_8),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_160),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_160),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_160),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_50),
.B1(n_64),
.B2(n_67),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_9),
.A2(n_50),
.B1(n_57),
.B2(n_60),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_12),
.A2(n_64),
.B1(n_67),
.B2(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_12),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_85),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_60),
.B1(n_85),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_85),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_13),
.A2(n_60),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_13),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_108),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_108),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_108),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_14),
.A2(n_40),
.B1(n_64),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_40),
.B1(n_73),
.B2(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_16),
.A2(n_27),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_16),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_16),
.A2(n_27),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_352),
.B(n_355),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_347),
.B(n_351),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_334),
.B(n_346),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_135),
.A3(n_149),
.B(n_331),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_113),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_22),
.B(n_113),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.C(n_92),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_23),
.A2(n_76),
.B1(n_77),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_23),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_52),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_24),
.A2(n_25),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_25),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_53),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_26),
.A2(n_35),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_26),
.A2(n_177),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_26),
.A2(n_97),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_26),
.A2(n_260),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_27),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_29),
.B1(n_45),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_28),
.B(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_39),
.A2(n_43),
.B1(n_51),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_42),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_41),
.B(n_252),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_42),
.A2(n_82),
.B(n_170),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_43),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_43),
.A2(n_51),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_43),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_43),
.A2(n_51),
.B1(n_227),
.B2(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_48),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_48),
.A2(n_88),
.B1(n_102),
.B2(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_48),
.B(n_170),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_48),
.A2(n_165),
.B(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_51),
.B(n_166),
.Y(n_228)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_56),
.A2(n_62),
.B1(n_110),
.B2(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_57),
.Y(n_169)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_68),
.Y(n_75)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_62),
.A2(n_110),
.B1(n_132),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_62),
.A2(n_69),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_63),
.A2(n_74),
.B1(n_107),
.B2(n_201),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_63),
.A2(n_74),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_63),
.A2(n_74),
.B1(n_342),
.B2(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_63),
.A2(n_74),
.B(n_349),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g67 ( 
.A(n_64),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_67),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_64),
.A2(n_68),
.B(n_171),
.C(n_181),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_SL g181 ( 
.A(n_66),
.B(n_67),
.C(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_73),
.B(n_170),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_74),
.A2(n_112),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_87),
.B(n_91),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_79),
.A2(n_80),
.B1(n_126),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_79),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_79),
.A2(n_198),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_80),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_80),
.A2(n_104),
.B(n_186),
.Y(n_310)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_88),
.A2(n_226),
.B(n_228),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_88),
.A2(n_228),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_92),
.A2(n_93),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_105),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_94),
.A2(n_95),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_96),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_98),
.B(n_170),
.Y(n_264)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_98),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_98),
.A2(n_234),
.B(n_258),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_103),
.B(n_105),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_110),
.B(n_111),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.C(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_131),
.B2(n_134),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_128),
.C(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_123),
.A2(n_124),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_124),
.B(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_128),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_128),
.B(n_142),
.C(n_146),
.Y(n_345)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_134),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_131),
.B(n_138),
.C(n_141),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_136),
.A2(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_148),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_137),
.B(n_148),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_143),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_147),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_324),
.B(n_330),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_314),
.B(n_323),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_213),
.B(n_297),
.C(n_313),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_193),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_153),
.B(n_193),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_172),
.C(n_183),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_154),
.A2(n_155),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_167),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_162),
.C(n_167),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B(n_171),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_172),
.A2(n_173),
.B1(n_183),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_183),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_190),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_192),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_202),
.B1(n_203),
.B2(n_212),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_194),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.CI(n_199),
.CON(n_194),
.SN(n_194)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_195),
.B(n_196),
.C(n_199),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_211),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_204),
.B(n_211),
.C(n_212),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_205),
.B(n_210),
.Y(n_311)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_290),
.B(n_296),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_245),
.B(n_289),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_237),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_237),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_236),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_219),
.B(n_225),
.C(n_229),
.Y(n_295)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.C(n_242),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_242),
.B1(n_243),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_283),
.B(n_288),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_273),
.B(n_282),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_261),
.B(n_272),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_268),
.B(n_271),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_281),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_281),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_287),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_295),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_312),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_312),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_302),
.C(n_304),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.C(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_340),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_338),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_340),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_350),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_353),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_348),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_354),
.B(n_357),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_356),
.Y(n_355)
);


endmodule