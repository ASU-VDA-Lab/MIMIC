module fake_jpeg_28178_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_45),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_39),
.Y(n_72)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_29),
.Y(n_88)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_59),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_35),
.B1(n_40),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_67),
.B1(n_54),
.B2(n_64),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_30),
.B1(n_22),
.B2(n_36),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_71),
.B1(n_24),
.B2(n_16),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_66),
.B(n_72),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_22),
.B1(n_41),
.B2(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_73),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_41),
.B1(n_28),
.B2(n_25),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_28),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_85),
.B1(n_87),
.B2(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_15),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_15),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_18),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_86),
.Y(n_95)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_17),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_44),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_91),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_37),
.C(n_19),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_62),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_23),
.B(n_27),
.C(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_14),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_113),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_45),
.B1(n_23),
.B2(n_27),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_108),
.B1(n_112),
.B2(n_74),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_16),
.B1(n_21),
.B2(n_37),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_59),
.B1(n_87),
.B2(n_63),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_37),
.C(n_29),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_69),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_65),
.A2(n_58),
.B1(n_32),
.B2(n_13),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_21),
.B1(n_16),
.B2(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_111),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_32),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_32),
.B1(n_12),
.B2(n_14),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_2),
.B(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_128),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_105),
.B1(n_109),
.B2(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_138),
.B1(n_106),
.B2(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_24),
.Y(n_132)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_115),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_68),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_159),
.B1(n_164),
.B2(n_167),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_95),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_175),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_92),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_126),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_101),
.C(n_95),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_155),
.C(n_126),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_99),
.B1(n_114),
.B2(n_118),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_171),
.B(n_122),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_117),
.A3(n_104),
.B1(n_89),
.B2(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_114),
.B1(n_100),
.B2(n_107),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_132),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_107),
.B1(n_85),
.B2(n_21),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_77),
.B1(n_29),
.B2(n_31),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_176),
.B1(n_144),
.B2(n_127),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_77),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_120),
.B1(n_130),
.B2(n_124),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_178),
.B1(n_127),
.B2(n_129),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_10),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_77),
.B1(n_31),
.B2(n_84),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_206),
.B1(n_148),
.B2(n_133),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_174),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_202),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_189),
.B(n_194),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_204),
.C(n_154),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_125),
.B(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_145),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_122),
.B(n_145),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_205),
.Y(n_228)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_207),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_203),
.Y(n_231)
);

XOR2x1_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_12),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_142),
.C(n_84),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_122),
.B(n_133),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_163),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_153),
.B1(n_159),
.B2(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_210),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_163),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_192),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_149),
.C(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_217),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_177),
.C(n_150),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_182),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_168),
.C(n_84),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_183),
.B1(n_199),
.B2(n_210),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_129),
.B1(n_84),
.B2(n_5),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_227),
.B1(n_205),
.B2(n_187),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_209),
.Y(n_250)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_237),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_252),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_253),
.B1(n_255),
.B2(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_184),
.B1(n_181),
.B2(n_202),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_257),
.B1(n_230),
.B2(n_236),
.Y(n_269)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_218),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_214),
.B(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_256),
.B(n_213),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_198),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_232),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_192),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_234),
.A2(n_184),
.B1(n_183),
.B2(n_195),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_190),
.B1(n_196),
.B2(n_193),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_197),
.B1(n_189),
.B2(n_191),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_185),
.B(n_212),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_211),
.B1(n_200),
.B2(n_5),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_223),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_261),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_252),
.B(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_257),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_218),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_248),
.C(n_216),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_290),
.C(n_288),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_286),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_250),
.B(n_249),
.C(n_213),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

A2O1A1O1Ixp25_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_255),
.B(n_245),
.C(n_246),
.D(n_243),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_287),
.B(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_242),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_253),
.B(n_220),
.C(n_241),
.D(n_217),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_221),
.C(n_222),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_262),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_294),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_277),
.A2(n_265),
.B1(n_261),
.B2(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_296),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_265),
.C(n_9),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_13),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_13),
.C(n_12),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_280),
.B1(n_289),
.B2(n_285),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_283),
.C(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_280),
.C(n_11),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_4),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_10),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_3),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_10),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_307),
.B(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_313),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_320),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_319),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_317),
.C(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.C(n_5),
.Y(n_326)
);

AOI221xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_6),
.B1(n_7),
.B2(n_225),
.C(n_185),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_6),
.Y(n_328)
);


endmodule