module fake_jpeg_27518_n_171 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_14),
.B(n_24),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_20),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_32),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_51),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_66),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_57),
.B1(n_15),
.B2(n_12),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_38),
.B1(n_30),
.B2(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_61),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_27),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_16),
.B(n_22),
.C(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_32),
.B(n_12),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_42),
.C(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_12),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_70),
.B(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_35),
.B1(n_60),
.B2(n_20),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_77),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_42),
.B(n_15),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_30),
.B1(n_37),
.B2(n_31),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_78),
.B1(n_59),
.B2(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_11),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_24),
.B1(n_14),
.B2(n_15),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_58),
.B1(n_50),
.B2(n_49),
.Y(n_78)
);

BUFx2_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_16),
.B1(n_14),
.B2(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_88),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_104),
.B1(n_68),
.B2(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_88),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_106),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_93),
.B1(n_91),
.B2(n_90),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_22),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_84),
.B1(n_86),
.B2(n_75),
.C(n_70),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_53),
.C(n_41),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_105),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_22),
.B1(n_19),
.B2(n_41),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_22),
.B(n_41),
.C(n_53),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_1),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_67),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_117),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_81),
.B1(n_75),
.B2(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_102),
.B(n_99),
.C(n_100),
.D(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_122),
.B(n_123),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_98),
.B1(n_102),
.B2(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_22),
.C(n_11),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_128),
.C(n_134),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_1),
.C(n_2),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_118),
.B(n_120),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_7),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_2),
.C(n_3),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_4),
.C(n_5),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_5),
.C(n_7),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_119),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_137),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_123),
.B1(n_117),
.B2(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_112),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_142),
.B(n_138),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.C(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_10),
.C(n_8),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_129),
.B(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_124),
.B(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_134),
.C(n_9),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_139),
.C(n_9),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_145),
.B1(n_147),
.B2(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_146),
.B1(n_8),
.B2(n_10),
.Y(n_160)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

NAND2x1p5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_157),
.B(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_162),
.B(n_153),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_167),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_169),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);


endmodule