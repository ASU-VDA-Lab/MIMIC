module fake_jpeg_16075_n_166 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_25),
.B1(n_24),
.B2(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_18),
.B1(n_29),
.B2(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_20),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_21),
.B1(n_15),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_16),
.B1(n_26),
.B2(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_21),
.B1(n_27),
.B2(n_15),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_59),
.B1(n_37),
.B2(n_19),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_33),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_70),
.B1(n_89),
.B2(n_42),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_40),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_84),
.C(n_92),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_85),
.B1(n_86),
.B2(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_57),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_40),
.B1(n_39),
.B2(n_16),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_40),
.B1(n_16),
.B2(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_18),
.B1(n_28),
.B2(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_28),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_42),
.B(n_46),
.C(n_18),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_113),
.B(n_63),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_18),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_28),
.B1(n_20),
.B2(n_30),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_6),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_79),
.B(n_70),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_121),
.B(n_95),
.C(n_30),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_73),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_1),
.C(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_119),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_73),
.CI(n_62),
.CON(n_118),
.SN(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_66),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_89),
.B(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_67),
.B1(n_87),
.B2(n_82),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_132),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_67),
.B1(n_82),
.B2(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_76),
.B1(n_64),
.B2(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_134),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_98),
.B1(n_104),
.B2(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_63),
.B1(n_8),
.B2(n_2),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_20),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_103),
.B1(n_109),
.B2(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_144),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_124),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_95),
.B(n_102),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_145),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_102),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_127),
.C(n_118),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_149),
.C(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_126),
.C(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_123),
.C(n_3),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_151),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_147),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_155),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_157),
.B(n_156),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_159),
.B(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_9),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_9),
.CI(n_11),
.CON(n_165),
.SN(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_12),
.Y(n_166)
);


endmodule