module real_jpeg_393_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g103 ( 
.A(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_48),
.Y(n_105)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_1),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_101),
.Y(n_220)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_2),
.B(n_26),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_2),
.B(n_60),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_4),
.B(n_38),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_4),
.B(n_31),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_4),
.B(n_48),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_4),
.B(n_60),
.Y(n_287)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_5),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_38),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_5),
.B(n_31),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_26),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_31),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_9),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_9),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_9),
.B(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_9),
.B(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_9),
.B(n_123),
.Y(n_197)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_11),
.B(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_11),
.B(n_48),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_11),
.B(n_101),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_79),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_11),
.B(n_123),
.Y(n_212)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_12),
.B(n_38),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_12),
.B(n_31),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_12),
.B(n_48),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_14),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_14),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_14),
.B(n_26),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI31xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.A3(n_161),
.B(n_321),
.Y(n_17)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_41),
.B(n_87),
.C(n_320),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_21),
.B(n_62),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_73),
.C(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_25),
.A2(n_40),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_26),
.Y(n_195)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_29),
.Y(n_321)
);

HAxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.CON(n_29),
.SN(n_29)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_43),
.C(n_46),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_30),
.B(n_191),
.C(n_198),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_30),
.A2(n_53),
.B1(n_198),
.B2(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_34),
.A2(n_35),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_35),
.B(n_100),
.C(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_37),
.B(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_43),
.A2(n_44),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_44),
.B(n_112),
.C(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_46),
.A2(n_47),
.B1(n_184),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.C(n_58),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_47),
.B(n_113),
.C(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g218 ( 
.A(n_48),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.C(n_55),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_58),
.A2(n_59),
.B1(n_77),
.B2(n_78),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_58),
.A2(n_59),
.B1(n_106),
.B2(n_146),
.Y(n_276)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_77),
.C(n_80),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_59),
.B(n_106),
.C(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_84),
.C(n_85),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_63),
.A2(n_64),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_76),
.C(n_81),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_65),
.A2(n_66),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_68),
.A2(n_69),
.B1(n_124),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_68),
.A2(n_69),
.B1(n_169),
.B2(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_120),
.C(n_124),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_69),
.B(n_163),
.C(n_169),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_73),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_73),
.B(n_164),
.C(n_166),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_73),
.A2(n_117),
.B1(n_164),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_76),
.B(n_81),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_78),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_77),
.B(n_95),
.C(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_77),
.A2(n_78),
.B1(n_255),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_78),
.B(n_255),
.C(n_256),
.Y(n_254)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_79),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_84),
.B(n_85),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_199),
.B(n_311),
.C(n_314),
.D(n_319),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_171),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_89),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_137),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_90),
.B(n_137),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_125),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_91),
.B(n_126),
.C(n_136),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_115),
.C(n_119),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_92),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.C(n_108),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_93),
.A2(n_94),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_100),
.B1(n_122),
.B2(n_152),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_104),
.B(n_108),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.C(n_107),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_107),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_111),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_112),
.A2(n_113),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_121),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_151),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_122),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_182)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_131),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_128),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_143),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_140),
.CI(n_143),
.CON(n_172),
.SN(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.C(n_162),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_158),
.CI(n_162),
.CON(n_174),
.SN(n_174)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_155),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_145),
.B(n_149),
.Y(n_236)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_152),
.B(n_153),
.C(n_154),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_150),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_150),
.A2(n_151),
.B1(n_252),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_154),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_155),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_168),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_172),
.B(n_173),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_172),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.C(n_178),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_174),
.B(n_175),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_174),
.Y(n_327)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_178),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.C(n_190),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_179),
.A2(n_180),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_185),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_181),
.B(n_183),
.CI(n_185),
.CON(n_265),
.SN(n_265)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_184),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_188),
.B(n_190),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_192),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_197),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_266),
.B(n_305),
.C(n_306),
.D(n_310),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_241),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_202),
.B(n_241),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_233),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_203),
.B(n_234),
.C(n_240),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_221),
.C(n_229),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_205),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_214),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_206),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_229),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_240),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_264),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_242),
.A2(n_264),
.B1(n_265),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.C(n_259),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_254),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_248),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_251),
.B1(n_254),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_257),
.A2(n_259),
.B1(n_260),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_265),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_299),
.B(n_304),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_291),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.C(n_281),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_269),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_274),
.CI(n_275),
.CON(n_269),
.SN(n_269)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_274),
.C(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.C(n_273),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.C(n_289),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_291),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.CI(n_296),
.CON(n_291),
.SN(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_303),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_308),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule