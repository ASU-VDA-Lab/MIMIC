module fake_netlist_6_1354_n_2086 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2086);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2086;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_52),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_113),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_108),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_26),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_75),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_123),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_157),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_73),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_31),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_195),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_197),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_173),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_168),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_158),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_26),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_54),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_72),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_160),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_24),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_88),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_207),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_109),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_79),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_182),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_5),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_4),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_59),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_172),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_183),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_218),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_94),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_10),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_19),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_105),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_103),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_79),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_147),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_46),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_144),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_161),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_18),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_151),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_116),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_82),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_180),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_152),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_134),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_46),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_227),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_201),
.Y(n_300)
);

INVxp33_ASAP7_75t_R g301 ( 
.A(n_70),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_32),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_80),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_229),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_29),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_119),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_154),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_27),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_10),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_184),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_65),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_83),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_143),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_66),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_202),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_159),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_57),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_93),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_193),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_86),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_104),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_57),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_127),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_84),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_92),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_122),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_135),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_78),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_138),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_18),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_62),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_64),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_64),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_81),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_107),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_83),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_74),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_23),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_100),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_176),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_118),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_89),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_42),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_11),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_129),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_169),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_128),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_222),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_120),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_209),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_215),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_115),
.Y(n_354)
);

INVxp33_ASAP7_75t_R g355 ( 
.A(n_13),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_102),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_140),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_136),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_73),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_75),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_53),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_117),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_44),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_178),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_192),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_12),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_60),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_15),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_24),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_22),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_165),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_204),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_69),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_175),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_6),
.Y(n_376)
);

BUFx8_ASAP7_75t_SL g377 ( 
.A(n_177),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_16),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_62),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_84),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_226),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_29),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_223),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_130),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_196),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_61),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_20),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_96),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_59),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_13),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_70),
.Y(n_391)
);

BUFx8_ASAP7_75t_SL g392 ( 
.A(n_213),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_87),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_41),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_58),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_208),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_211),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_200),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_131),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_230),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_8),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_3),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_112),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_142),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_114),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_155),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_9),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_148),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_101),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_98),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_188),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_42),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_174),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_164),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_36),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_179),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_47),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_91),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_225),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_81),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_181),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_39),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_216),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_54),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_3),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_28),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_121),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_77),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_191),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_166),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_206),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_162),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_214),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_219),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_30),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_16),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_67),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_56),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_203),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_14),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_99),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_149),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_47),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_106),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_60),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_19),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_186),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_63),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_217),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_7),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_39),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_167),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_30),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_224),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_163),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_126),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_11),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_12),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_137),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_292),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_314),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_271),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_277),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_334),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_292),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_274),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_292),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_280),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_292),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_292),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_284),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_286),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_292),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_292),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_289),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_292),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_297),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_339),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_243),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_245),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_339),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_293),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_234),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_245),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_234),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_279),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_383),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_234),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_279),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_234),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_234),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_319),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_388),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_319),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_319),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_319),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_319),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_249),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_406),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_401),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_303),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_305),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_249),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_283),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_411),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_239),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_306),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_401),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_240),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_257),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_239),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_283),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_281),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_298),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_310),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_290),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_246),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_332),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_309),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_313),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_333),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_256),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_335),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_336),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_338),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_345),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_316),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_324),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_346),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_369),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_370),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_374),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_256),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_270),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_326),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_320),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_379),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_330),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_340),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_264),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_239),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_386),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_391),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_261),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_360),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_422),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_261),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_270),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_361),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_435),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_363),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_320),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_261),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_367),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_453),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_290),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_368),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_413),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_341),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_371),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_302),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_246),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_390),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_320),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_390),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_382),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_302),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_425),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_431),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_425),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_302),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_377),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_359),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_389),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_394),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_417),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_237),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_395),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_565),
.B(n_328),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_461),
.B(n_480),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_487),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_490),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_490),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_494),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_507),
.B(n_259),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_582),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_543),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_461),
.B(n_237),
.Y(n_600)
);

NOR2x1_ASAP7_75t_L g601 ( 
.A(n_492),
.B(n_311),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_488),
.B(n_328),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_519),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_523),
.B(n_237),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_464),
.A2(n_273),
.B1(n_378),
.B2(n_312),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_493),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_493),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_491),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_496),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_543),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_465),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_462),
.B(n_407),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_497),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_568),
.B(n_342),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_486),
.B(n_343),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_466),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_467),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_500),
.B(n_244),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_560),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_498),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_498),
.B(n_311),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_587),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_499),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_499),
.Y(n_629)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_518),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_470),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_473),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_501),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_501),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_474),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_474),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_503),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_477),
.B(n_342),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_481),
.B(n_427),
.Y(n_640)
);

BUFx8_ASAP7_75t_L g641 ( 
.A(n_507),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_503),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_506),
.B(n_441),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_560),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_506),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_573),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_483),
.B(n_342),
.Y(n_647)
);

XNOR2x1_ASAP7_75t_L g648 ( 
.A(n_547),
.B(n_272),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_573),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_513),
.B(n_418),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_485),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_484),
.B(n_418),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_511),
.A2(n_449),
.B(n_441),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_463),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_514),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_524),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_524),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_466),
.B(n_272),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_478),
.B(n_418),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_571),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_572),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_572),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_574),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_478),
.B(n_247),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_529),
.B(n_248),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_580),
.B(n_380),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_577),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_489),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_579),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_580),
.B(n_275),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_516),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_520),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_522),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_525),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_588),
.B(n_449),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_528),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_531),
.B(n_236),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_637),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_651),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_623),
.B(n_515),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_604),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_651),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_667),
.B(n_468),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_637),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_603),
.B(n_468),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_630),
.B(n_548),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_630),
.B(n_619),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_598),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_636),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_636),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_636),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_636),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_651),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_659),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_632),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_604),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_612),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_638),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_638),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_654),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_638),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_632),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_627),
.B(n_570),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_603),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_633),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_681),
.B(n_588),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_633),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_671),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_610),
.B(n_471),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_612),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_598),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_612),
.B(n_471),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_612),
.B(n_472),
.Y(n_725)
);

BUFx6f_ASAP7_75t_SL g726 ( 
.A(n_627),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_609),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_609),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_682),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_682),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_598),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_599),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_659),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_682),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_599),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_599),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_590),
.B(n_475),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_602),
.B(n_475),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_662),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_674),
.B(n_540),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_609),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_662),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_644),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_658),
.B(n_482),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_644),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_600),
.B(n_482),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_662),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_662),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_662),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_663),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_665),
.A2(n_479),
.B1(n_540),
.B2(n_541),
.Y(n_754)
);

OAI22x1_ASAP7_75t_L g755 ( 
.A1(n_606),
.A2(n_551),
.B1(n_554),
.B2(n_510),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_663),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_591),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_665),
.A2(n_458),
.B1(n_428),
.B2(n_295),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_648),
.A2(n_376),
.B1(n_238),
.B2(n_258),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_613),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_663),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_663),
.Y(n_762)
);

NOR2x1p5_ASAP7_75t_L g763 ( 
.A(n_596),
.B(n_420),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_613),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_674),
.B(n_586),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_592),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_592),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_641),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_618),
.B(n_586),
.Y(n_769)
);

AO21x2_ASAP7_75t_L g770 ( 
.A1(n_653),
.A2(n_260),
.B(n_235),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_596),
.B(n_504),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_663),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_593),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_598),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_626),
.A2(n_643),
.B1(n_669),
.B2(n_618),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_613),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_647),
.B(n_555),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_663),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_639),
.B(n_504),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_650),
.A2(n_576),
.B1(n_512),
.B2(n_526),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_593),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_684),
.B(n_505),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_594),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_664),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_613),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_613),
.B(n_505),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_594),
.Y(n_787)
);

XOR2x2_ASAP7_75t_L g788 ( 
.A(n_606),
.B(n_301),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_664),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_644),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_684),
.B(n_512),
.Y(n_791)
);

AND3x1_ASAP7_75t_L g792 ( 
.A(n_669),
.B(n_355),
.C(n_532),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_647),
.B(n_533),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_652),
.B(n_527),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_605),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_605),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_607),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_607),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_620),
.B(n_527),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_664),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_652),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_608),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_641),
.B(n_534),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_641),
.B(n_534),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_664),
.Y(n_805)
);

BUFx6f_ASAP7_75t_SL g806 ( 
.A(n_626),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_644),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_608),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_589),
.B(n_535),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_611),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_664),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_641),
.B(n_542),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_653),
.A2(n_276),
.B(n_265),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_656),
.B(n_536),
.Y(n_814)
);

AND3x2_ASAP7_75t_L g815 ( 
.A(n_626),
.B(n_581),
.C(n_562),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_611),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_615),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_615),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_621),
.B(n_542),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_597),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_646),
.Y(n_821)
);

AND3x2_ASAP7_75t_L g822 ( 
.A(n_626),
.B(n_583),
.C(n_304),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_672),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_675),
.B(n_545),
.Y(n_824)
);

AND3x2_ASAP7_75t_L g825 ( 
.A(n_643),
.B(n_308),
.C(n_285),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_616),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_643),
.A2(n_538),
.B1(n_539),
.B2(n_537),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_648),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_L g829 ( 
.A(n_640),
.B(n_549),
.C(n_544),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_589),
.B(n_545),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_675),
.B(n_546),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_676),
.B(n_585),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_616),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_646),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_676),
.B(n_553),
.C(n_550),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_672),
.Y(n_836)
);

INVx5_ASAP7_75t_L g837 ( 
.A(n_621),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_677),
.B(n_546),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_648),
.Y(n_839)
);

NOR2x1_ASAP7_75t_L g840 ( 
.A(n_601),
.B(n_315),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_672),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_617),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_672),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_677),
.B(n_552),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_L g845 ( 
.A(n_689),
.B(n_320),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_706),
.B(n_721),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_745),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_706),
.B(n_721),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_691),
.B(n_556),
.C(n_552),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_814),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_621),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_742),
.B(n_556),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_714),
.B(n_621),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_771),
.B(n_688),
.C(n_799),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_693),
.B(n_559),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_705),
.A2(n_502),
.B1(n_509),
.B2(n_495),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_745),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_705),
.B(n_621),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_733),
.B(n_320),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_733),
.B(n_621),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_814),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_782),
.B(n_622),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_791),
.B(n_622),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_801),
.A2(n_679),
.B(n_680),
.C(n_678),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_738),
.B(n_559),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_801),
.B(n_622),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_759),
.A2(n_770),
.B1(n_813),
.B2(n_765),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_703),
.B(n_622),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_809),
.B(n_830),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_703),
.B(n_622),
.Y(n_870)
);

AND2x6_ASAP7_75t_L g871 ( 
.A(n_697),
.B(n_698),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_775),
.B(n_631),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_746),
.B(n_563),
.Y(n_873)
);

INVx4_ASAP7_75t_SL g874 ( 
.A(n_806),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_724),
.B(n_725),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_749),
.A2(n_578),
.B1(n_567),
.B2(n_362),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_765),
.A2(n_679),
.B(n_680),
.C(n_678),
.Y(n_877)
);

INVxp33_ASAP7_75t_L g878 ( 
.A(n_742),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_777),
.B(n_563),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_844),
.B(n_566),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_786),
.B(n_631),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_844),
.B(n_566),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_729),
.B(n_631),
.Y(n_883)
);

CKINVDCx16_ASAP7_75t_R g884 ( 
.A(n_820),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_819),
.B(n_320),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_769),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_834),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_831),
.B(n_569),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_839),
.B(n_569),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_757),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_766),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_766),
.B(n_643),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_838),
.B(n_720),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_697),
.A2(n_625),
.B(n_628),
.C(n_617),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_824),
.B(n_575),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_737),
.B(n_575),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_723),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_767),
.B(n_646),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_767),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_793),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_773),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_716),
.A2(n_585),
.B1(n_584),
.B2(n_385),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_773),
.B(n_646),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_781),
.B(n_649),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_L g905 ( 
.A(n_840),
.B(n_320),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_745),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_780),
.B(n_584),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_781),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_794),
.B(n_294),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_698),
.B(n_262),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_695),
.B(n_779),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_713),
.B(n_409),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_783),
.B(n_649),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_792),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_723),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_727),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_787),
.B(n_649),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_795),
.B(n_625),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_754),
.A2(n_421),
.B1(n_331),
.B2(n_348),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_729),
.B(n_262),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_795),
.B(n_628),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_796),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_796),
.B(n_629),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_797),
.B(n_629),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_797),
.B(n_634),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_792),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_839),
.B(n_614),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_730),
.B(n_262),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_282),
.B1(n_287),
.B2(n_278),
.Y(n_929)
);

BUFx6f_ASAP7_75t_SL g930 ( 
.A(n_820),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_798),
.B(n_802),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_798),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_763),
.A2(n_291),
.B1(n_296),
.B2(n_288),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_802),
.B(n_634),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_730),
.B(n_262),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_732),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_734),
.B(n_262),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_808),
.B(n_635),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_808),
.B(n_635),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_815),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_810),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_735),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_840),
.B(n_329),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_816),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_816),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_759),
.A2(n_357),
.B1(n_372),
.B2(n_405),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_817),
.B(n_645),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_832),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_817),
.B(n_645),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_747),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_806),
.A2(n_318),
.B1(n_299),
.B2(n_300),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_SL g952 ( 
.A(n_768),
.B(n_392),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_726),
.B(n_241),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_822),
.B(n_818),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_806),
.A2(n_381),
.B1(n_366),
.B2(n_364),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_818),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_826),
.B(n_666),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_726),
.B(n_241),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_735),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_826),
.B(n_666),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_833),
.B(n_666),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_833),
.B(n_666),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_709),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_758),
.B(n_412),
.C(n_402),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_734),
.B(n_357),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_825),
.Y(n_966)
);

NOR3xp33_ASAP7_75t_L g967 ( 
.A(n_828),
.B(n_558),
.C(n_557),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_842),
.A2(n_683),
.B(n_561),
.C(n_564),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_842),
.Y(n_969)
);

NAND3x1_ASAP7_75t_L g970 ( 
.A(n_788),
.B(n_614),
.C(n_354),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_739),
.B(n_357),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_739),
.B(n_357),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_768),
.B(n_242),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_709),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_726),
.A2(n_373),
.B1(n_307),
.B2(n_317),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_699),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_699),
.B(n_672),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_700),
.Y(n_978)
);

CKINVDCx16_ASAP7_75t_R g979 ( 
.A(n_820),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_700),
.B(n_242),
.Y(n_980)
);

OAI22xp33_ASAP7_75t_SL g981 ( 
.A1(n_828),
.A2(n_445),
.B1(n_426),
.B2(n_457),
.Y(n_981)
);

BUFx6f_ASAP7_75t_SL g982 ( 
.A(n_820),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_696),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_759),
.B(n_683),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_759),
.A2(n_357),
.B1(n_372),
.B2(n_358),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_755),
.A2(n_397),
.B1(n_321),
.B2(n_322),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_747),
.B(n_672),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_827),
.B(n_250),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_719),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_747),
.B(n_655),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_790),
.B(n_372),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_736),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_727),
.B(n_372),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_L g994 ( 
.A(n_829),
.B(n_655),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_790),
.B(n_642),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_790),
.B(n_642),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_807),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_869),
.A2(n_821),
.B1(n_807),
.B2(n_804),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_893),
.B(n_807),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_976),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_893),
.B(n_821),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_900),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_916),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_963),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_978),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_855),
.A2(n_803),
.B1(n_812),
.B2(n_755),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_855),
.A2(n_748),
.B1(n_785),
.B2(n_728),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_884),
.B(n_719),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_874),
.B(n_835),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_847),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_946),
.A2(n_829),
.B(n_835),
.C(n_403),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_875),
.A2(n_687),
.B(n_685),
.Y(n_1012)
);

AND2x6_ASAP7_75t_SL g1013 ( 
.A(n_896),
.B(n_788),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_974),
.Y(n_1014)
);

BUFx8_ASAP7_75t_L g1015 ( 
.A(n_930),
.Y(n_1015)
);

OAI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_850),
.A2(n_424),
.B1(n_426),
.B2(n_420),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_865),
.A2(n_748),
.B1(n_785),
.B2(n_728),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_875),
.B(n_727),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_890),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_888),
.B(n_687),
.Y(n_1020)
);

INVxp33_ASAP7_75t_SL g1021 ( 
.A(n_856),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_865),
.A2(n_748),
.B1(n_785),
.B2(n_728),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_878),
.B(n_694),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_891),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_888),
.B(n_692),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_900),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_847),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_SL g1028 ( 
.A(n_979),
.B(n_250),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_899),
.B(n_692),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_901),
.B(n_704),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_862),
.B(n_863),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_857),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_861),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_857),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_911),
.A2(n_880),
.B1(n_882),
.B2(n_854),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_908),
.B(n_704),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_916),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_922),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_932),
.B(n_710),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_852),
.B(n_879),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_954),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_989),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_886),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_911),
.A2(n_712),
.B1(n_715),
.B2(n_710),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_954),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_880),
.A2(n_715),
.B1(n_717),
.B2(n_712),
.Y(n_1046)
);

AND2x6_ASAP7_75t_SL g1047 ( 
.A(n_896),
.B(n_353),
.Y(n_1047)
);

OR2x2_ASAP7_75t_SL g1048 ( 
.A(n_964),
.B(n_927),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_872),
.A2(n_718),
.B(n_717),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_941),
.B(n_718),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_914),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_906),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_906),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_950),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_944),
.B(n_740),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_945),
.B(n_740),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_956),
.B(n_741),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_950),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_969),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_931),
.B(n_741),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_889),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_846),
.B(n_744),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_882),
.A2(n_750),
.B1(n_751),
.B2(n_744),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_867),
.B(n_760),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_997),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_848),
.B(n_750),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_909),
.B(n_359),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_984),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_966),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_L g1070 ( 
.A(n_940),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_874),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_871),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_871),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_948),
.B(n_415),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_946),
.A2(n_459),
.B(n_454),
.C(n_430),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_982),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_926),
.A2(n_843),
.B1(n_841),
.B2(n_836),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_851),
.B(n_853),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_912),
.A2(n_772),
.B1(n_823),
.B2(n_753),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_985),
.A2(n_444),
.B(n_452),
.C(n_433),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_874),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_881),
.A2(n_764),
.B(n_760),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_867),
.B(n_764),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_868),
.B(n_656),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_982),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_912),
.A2(n_751),
.B1(n_823),
.B2(n_752),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_868),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_970),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_873),
.B(n_424),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_870),
.B(n_661),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_876),
.Y(n_1091)
);

AND2x4_ASAP7_75t_SL g1092 ( 
.A(n_967),
.B(n_359),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_887),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_870),
.B(n_661),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_994),
.B(n_670),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_858),
.B(n_752),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_990),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_871),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_892),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_860),
.B(n_670),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_871),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_897),
.Y(n_1102)
);

AND2x2_ASAP7_75t_SL g1103 ( 
.A(n_985),
.B(n_753),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_980),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_871),
.Y(n_1105)
);

NOR2x1p5_ASAP7_75t_L g1106 ( 
.A(n_952),
.B(n_436),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_953),
.B(n_756),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_860),
.B(n_764),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_918),
.B(n_761),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_895),
.B(n_907),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_921),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_943),
.B(n_764),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_943),
.B(n_776),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_915),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_923),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_924),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_866),
.B(n_776),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_925),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_934),
.B(n_761),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_988),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_936),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_902),
.Y(n_1122)
);

AND2x2_ASAP7_75t_SL g1123 ( 
.A(n_905),
.B(n_762),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_919),
.A2(n_813),
.B1(n_770),
.B2(n_372),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_938),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_939),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_942),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_895),
.B(n_776),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_SL g1129 ( 
.A1(n_986),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_947),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_SL g1131 ( 
.A1(n_953),
.A2(n_437),
.B1(n_438),
.B2(n_440),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_959),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_949),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_992),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_845),
.A2(n_813),
.B1(n_770),
.B2(n_372),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_929),
.B(n_772),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_957),
.A2(n_778),
.B1(n_811),
.B2(n_805),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_973),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_849),
.B(n_440),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_955),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_958),
.B(n_445),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_960),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_933),
.A2(n_961),
.B1(n_962),
.B2(n_975),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_951),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_898),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_991),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_883),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_903),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_877),
.B(n_778),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_991),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_864),
.B(n_904),
.Y(n_1151)
);

AND2x4_ASAP7_75t_SL g1152 ( 
.A(n_958),
.B(n_776),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_894),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_913),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_977),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_859),
.A2(n_885),
.B1(n_917),
.B2(n_883),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_987),
.B(n_784),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_995),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_996),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_983),
.B(n_789),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_920),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_SL g1162 ( 
.A(n_968),
.B(n_252),
.C(n_251),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1110),
.A2(n_965),
.B(n_935),
.C(n_972),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1101),
.B(n_983),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1035),
.B(n_981),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1110),
.A2(n_935),
.B(n_972),
.C(n_971),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1091),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1042),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1078),
.A2(n_993),
.B(n_800),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_1061),
.B(n_928),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1040),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1012),
.A2(n_800),
.B(n_928),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1031),
.A2(n_965),
.B(n_937),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1089),
.B(n_1067),
.C(n_1074),
.Y(n_1174)
);

CKINVDCx6p67_ASAP7_75t_R g1175 ( 
.A(n_1014),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1025),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1113),
.A2(n_624),
.B(n_598),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1004),
.Y(n_1178)
);

AND2x2_ASAP7_75t_SL g1179 ( 
.A(n_1122),
.B(n_657),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1049),
.A2(n_624),
.B(n_702),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1114),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_SL g1182 ( 
.A1(n_1128),
.A2(n_910),
.B(n_601),
.C(n_372),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1115),
.B(n_707),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1025),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1021),
.A2(n_414),
.B1(n_323),
.B2(n_325),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1132),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1051),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1134),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1144),
.A2(n_1089),
.B1(n_1139),
.B2(n_1141),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1104),
.A2(n_711),
.B(n_708),
.C(n_707),
.Y(n_1190)
);

OA22x2_ASAP7_75t_L g1191 ( 
.A1(n_1006),
.A2(n_457),
.B1(n_451),
.B2(n_266),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1071),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1104),
.B(n_254),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1116),
.B(n_255),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1118),
.B(n_708),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1043),
.B(n_263),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1125),
.B(n_263),
.Y(n_1197)
);

AO32x1_ASAP7_75t_L g1198 ( 
.A1(n_998),
.A2(n_686),
.A3(n_701),
.B1(n_690),
.B2(n_711),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1134),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1069),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1002),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1020),
.A2(n_1130),
.B1(n_1133),
.B2(n_1126),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1074),
.A2(n_267),
.B(n_266),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1111),
.B(n_1099),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1064),
.A2(n_690),
.B(n_686),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1087),
.A2(n_267),
.B(n_268),
.C(n_269),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1041),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1111),
.B(n_701),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_999),
.A2(n_268),
.B1(n_269),
.B2(n_419),
.Y(n_1209)
);

AO22x1_ASAP7_75t_L g1210 ( 
.A1(n_1023),
.A2(n_419),
.B1(n_423),
.B2(n_429),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1043),
.B(n_423),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1099),
.B(n_657),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1026),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1001),
.A2(n_673),
.B(n_668),
.C(n_660),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1120),
.A2(n_429),
.B(n_434),
.C(n_439),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1082),
.A2(n_673),
.B(n_668),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1064),
.A2(n_910),
.B(n_837),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1101),
.A2(n_434),
.B1(n_439),
.B2(n_442),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1019),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1105),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1097),
.B(n_660),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1128),
.A2(n_668),
.B(n_673),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1068),
.B(n_660),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1011),
.A2(n_372),
.B(n_910),
.C(n_2),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_L g1225 ( 
.A1(n_1018),
.A2(n_910),
.B(n_722),
.C(n_774),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_R g1226 ( 
.A(n_1008),
.B(n_442),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1070),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1024),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1015),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1008),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_1083),
.A2(n_0),
.B(n_1),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_SL g1232 ( 
.A(n_1071),
.B(n_447),
.Y(n_1232)
);

OR2x6_ASAP7_75t_SL g1233 ( 
.A(n_1076),
.B(n_455),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1038),
.B(n_455),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1003),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1059),
.B(n_456),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1011),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1000),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1093),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1023),
.A2(n_398),
.B1(n_337),
.B2(n_344),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1101),
.A2(n_400),
.B1(n_347),
.B2(n_349),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1151),
.A2(n_837),
.B(n_743),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1140),
.B(n_327),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1146),
.A2(n_396),
.B(n_351),
.C(n_352),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1142),
.B(n_350),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1033),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1157),
.A2(n_837),
.B(n_212),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1155),
.B(n_356),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1003),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1138),
.B(n_365),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1155),
.B(n_375),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1083),
.A2(n_1123),
.B(n_1060),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_SL g1253 ( 
.A(n_1016),
.B(n_416),
.C(n_410),
.Y(n_1253)
);

AND2x2_ASAP7_75t_SL g1254 ( 
.A(n_1028),
.B(n_4),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1048),
.B(n_384),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1013),
.B(n_393),
.Y(n_1256)
);

BUFx4_ASAP7_75t_SL g1257 ( 
.A(n_1085),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1009),
.B(n_404),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1123),
.A2(n_774),
.B(n_731),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1145),
.B(n_408),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1148),
.B(n_595),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1009),
.B(n_595),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1095),
.B(n_595),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1005),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1062),
.A2(n_774),
.B(n_731),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1003),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1066),
.A2(n_774),
.B(n_731),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1112),
.A2(n_595),
.B(n_642),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1096),
.A2(n_731),
.B(n_722),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1154),
.B(n_595),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1084),
.B(n_595),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1084),
.B(n_642),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1030),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1150),
.A2(n_642),
.B(n_7),
.C(n_8),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1109),
.A2(n_696),
.B(n_232),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1129),
.A2(n_6),
.B1(n_9),
.B2(n_15),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1045),
.B(n_17),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1034),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1090),
.B(n_17),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1137),
.A2(n_145),
.B(n_231),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_R g1281 ( 
.A(n_1081),
.B(n_228),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1119),
.A2(n_696),
.B(n_221),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1075),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1283)
);

BUFx12f_ASAP7_75t_L g1284 ( 
.A(n_1015),
.Y(n_1284)
);

OAI21xp33_ASAP7_75t_L g1285 ( 
.A1(n_1092),
.A2(n_25),
.B(n_27),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1105),
.B(n_205),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1103),
.A2(n_198),
.B1(n_194),
.B2(n_185),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1070),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1088),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1136),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1092),
.B(n_33),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1095),
.B(n_33),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1105),
.B(n_171),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1094),
.B(n_34),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1105),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1158),
.B(n_34),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1136),
.A2(n_170),
.B1(n_156),
.B2(n_146),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1143),
.B(n_141),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1036),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1131),
.B(n_35),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1301)
);

INVx4_ASAP7_75t_L g1302 ( 
.A(n_1003),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1171),
.B(n_1207),
.Y(n_1303)
);

O2A1O1Ixp5_ASAP7_75t_L g1304 ( 
.A1(n_1298),
.A2(n_1143),
.B(n_1080),
.C(n_1075),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_1159),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1216),
.A2(n_1222),
.B(n_1172),
.Y(n_1306)
);

O2A1O1Ixp5_ASAP7_75t_L g1307 ( 
.A1(n_1174),
.A2(n_1080),
.B(n_1149),
.C(n_1153),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1243),
.A2(n_1106),
.B1(n_1107),
.B2(n_1016),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1299),
.B(n_1100),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1204),
.B(n_1100),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1255),
.A2(n_1156),
.B(n_1124),
.C(n_1152),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1247),
.A2(n_1117),
.B(n_1108),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1252),
.A2(n_1124),
.B(n_1135),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1202),
.B(n_1039),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1301),
.B(n_1050),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1293),
.B(n_1072),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1168),
.B(n_1102),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1252),
.A2(n_1135),
.B(n_1046),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1179),
.B(n_1152),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1183),
.B(n_1029),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1189),
.A2(n_1017),
.B1(n_1022),
.B2(n_1007),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1165),
.B(n_1219),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1300),
.A2(n_1162),
.B(n_1065),
.C(n_1055),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1228),
.B(n_1010),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1246),
.B(n_1027),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1169),
.A2(n_1180),
.B(n_1242),
.Y(n_1326)
);

BUFx2_ASAP7_75t_SL g1327 ( 
.A(n_1288),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1178),
.Y(n_1328)
);

NAND3x1_ASAP7_75t_L g1329 ( 
.A(n_1256),
.B(n_1291),
.C(n_1277),
.Y(n_1329)
);

AO21x1_ASAP7_75t_L g1330 ( 
.A1(n_1237),
.A2(n_1056),
.B(n_1057),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1238),
.B(n_1264),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1245),
.B(n_1032),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1203),
.A2(n_1166),
.B(n_1163),
.C(n_1253),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1187),
.B(n_1147),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1181),
.Y(n_1335)
);

NAND3xp33_ASAP7_75t_L g1336 ( 
.A(n_1290),
.B(n_1063),
.C(n_1044),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1193),
.B(n_1047),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1173),
.A2(n_1037),
.B(n_1160),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1257),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1250),
.A2(n_1162),
.B1(n_1073),
.B2(n_1072),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1258),
.A2(n_1098),
.B1(n_1052),
.B2(n_1053),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1239),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1192),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1254),
.B(n_1147),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1249),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1163),
.A2(n_1079),
.B(n_1086),
.C(n_1077),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1186),
.Y(n_1347)
);

BUFx2_ASAP7_75t_SL g1348 ( 
.A(n_1227),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1260),
.B(n_1054),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1175),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1188),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1212),
.B(n_1058),
.Y(n_1352)
);

AOI31xp67_ASAP7_75t_L g1353 ( 
.A1(n_1191),
.A2(n_1161),
.A3(n_1127),
.B(n_1147),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1276),
.A2(n_1147),
.B1(n_1121),
.B2(n_37),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1279),
.B(n_1121),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1199),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1280),
.A2(n_139),
.B(n_133),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1285),
.B(n_35),
.C(n_36),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1166),
.A2(n_125),
.B(n_124),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1194),
.A2(n_38),
.B(n_40),
.C(n_43),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1294),
.B(n_1196),
.Y(n_1361)
);

AO21x1_ASAP7_75t_L g1362 ( 
.A1(n_1237),
.A2(n_40),
.B(n_44),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_SL g1363 ( 
.A1(n_1274),
.A2(n_1244),
.B(n_1287),
.C(n_1206),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1164),
.A2(n_111),
.B(n_110),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1211),
.B(n_1234),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1276),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1201),
.Y(n_1367)
);

AOI22x1_ASAP7_75t_SL g1368 ( 
.A1(n_1230),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1275),
.A2(n_95),
.B(n_52),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1192),
.B(n_51),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1182),
.A2(n_53),
.B(n_55),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1197),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1275),
.A2(n_61),
.B(n_63),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1278),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1282),
.A2(n_66),
.B(n_67),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1231),
.A2(n_68),
.A3(n_71),
.B(n_74),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1176),
.B(n_68),
.C(n_71),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1289),
.B(n_76),
.Y(n_1378)
);

BUFx12f_ASAP7_75t_L g1379 ( 
.A(n_1229),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1282),
.A2(n_76),
.A3(n_77),
.B(n_78),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1213),
.B(n_80),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1292),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1200),
.B(n_1236),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1296),
.A2(n_82),
.A3(n_85),
.B(n_1198),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1265),
.A2(n_85),
.B(n_1267),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1214),
.A2(n_1190),
.B(n_1221),
.Y(n_1386)
);

NOR4xp25_ASAP7_75t_L g1387 ( 
.A(n_1283),
.B(n_1224),
.C(n_1184),
.D(n_1214),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1249),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1185),
.B(n_1232),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1195),
.B(n_1210),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1284),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1167),
.B(n_1191),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1208),
.B(n_1170),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1261),
.A2(n_1270),
.B(n_1265),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1209),
.B(n_1240),
.Y(n_1396)
);

BUFx2_ASAP7_75t_R g1397 ( 
.A(n_1233),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_SL g1398 ( 
.A(n_1293),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1223),
.B(n_1215),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1293),
.A2(n_1297),
.B1(n_1262),
.B2(n_1224),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1267),
.A2(n_1272),
.B(n_1269),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1190),
.A2(n_1225),
.B(n_1217),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1283),
.A2(n_1220),
.B1(n_1295),
.B2(n_1286),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1271),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1225),
.A2(n_1259),
.B(n_1269),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1220),
.B(n_1295),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1198),
.A2(n_1259),
.A3(n_1177),
.B(n_1218),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1198),
.A2(n_1263),
.B(n_1177),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1249),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1266),
.Y(n_1410)
);

AND3x4_ASAP7_75t_L g1411 ( 
.A(n_1226),
.B(n_1281),
.C(n_1286),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1241),
.B(n_1235),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1235),
.A2(n_1302),
.B(n_1205),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1266),
.A2(n_869),
.B1(n_893),
.B2(n_1035),
.Y(n_1414)
);

INVxp67_ASAP7_75t_SL g1415 ( 
.A(n_1266),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1302),
.B(n_1205),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1268),
.A2(n_1031),
.B(n_1180),
.Y(n_1417)
);

AO32x2_ASAP7_75t_L g1418 ( 
.A1(n_1202),
.A2(n_919),
.A3(n_1287),
.B1(n_1068),
.B2(n_998),
.Y(n_1418)
);

AOI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1174),
.A2(n_1110),
.B(n_869),
.Y(n_1419)
);

AOI221x1_ASAP7_75t_L g1420 ( 
.A1(n_1174),
.A2(n_1110),
.B1(n_893),
.B2(n_869),
.C(n_1252),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1252),
.A2(n_1049),
.B(n_1173),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_SL g1422 ( 
.A1(n_1298),
.A2(n_1011),
.B(n_1080),
.C(n_1075),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1216),
.A2(n_1222),
.B(n_1172),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1293),
.B(n_1071),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1168),
.B(n_927),
.Y(n_1425)
);

OAI22x1_ASAP7_75t_L g1426 ( 
.A1(n_1174),
.A2(n_1006),
.B1(n_1035),
.B2(n_1091),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1178),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1216),
.A2(n_1222),
.B(n_1172),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1174),
.A2(n_869),
.B1(n_893),
.B2(n_1035),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1252),
.A2(n_1049),
.B(n_1173),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1239),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1273),
.B(n_893),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1192),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1257),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1168),
.B(n_927),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1273),
.B(n_893),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1174),
.B(n_869),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1174),
.B(n_974),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1178),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1192),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1273),
.B(n_893),
.Y(n_1441)
);

INVx3_ASAP7_75t_SL g1442 ( 
.A(n_1339),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1434),
.Y(n_1443)
);

OAI211xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1419),
.A2(n_1308),
.B(n_1365),
.C(n_1361),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1425),
.B(n_1435),
.Y(n_1445)
);

OAI211xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1419),
.A2(n_1441),
.B(n_1432),
.C(n_1436),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1429),
.B(n_1437),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1316),
.Y(n_1448)
);

INVx4_ASAP7_75t_SL g1449 ( 
.A(n_1398),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1429),
.A2(n_1424),
.B1(n_1396),
.B2(n_1316),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1328),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1390),
.A2(n_1333),
.B(n_1311),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1401),
.A2(n_1405),
.B(n_1338),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1316),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1439),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1431),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1417),
.A2(n_1312),
.B(n_1395),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1317),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1358),
.A2(n_1377),
.B1(n_1366),
.B2(n_1426),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1367),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_SL g1462 ( 
.A(n_1337),
.B(n_1373),
.C(n_1389),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1402),
.A2(n_1385),
.B(n_1408),
.Y(n_1463)
);

AO32x2_ASAP7_75t_L g1464 ( 
.A1(n_1366),
.A2(n_1354),
.A3(n_1414),
.B1(n_1321),
.B2(n_1400),
.Y(n_1464)
);

NAND2x1_ASAP7_75t_L g1465 ( 
.A(n_1424),
.B(n_1440),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1373),
.A2(n_1371),
.B(n_1362),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1335),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1358),
.B(n_1420),
.C(n_1377),
.Y(n_1468)
);

CKINVDCx6p67_ASAP7_75t_R g1469 ( 
.A(n_1379),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1411),
.A2(n_1398),
.B1(n_1414),
.B2(n_1400),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1383),
.A2(n_1329),
.B1(n_1438),
.B2(n_1344),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1354),
.A2(n_1336),
.B1(n_1321),
.B2(n_1393),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1392),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1322),
.A2(n_1427),
.B1(n_1319),
.B2(n_1309),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1330),
.A2(n_1346),
.A3(n_1403),
.B(n_1416),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1409),
.Y(n_1476)
);

AO221x2_ASAP7_75t_L g1477 ( 
.A1(n_1359),
.A2(n_1371),
.B1(n_1313),
.B2(n_1318),
.C(n_1336),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1304),
.A2(n_1314),
.B(n_1323),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1413),
.A2(n_1386),
.B(n_1307),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1318),
.A2(n_1314),
.B(n_1360),
.C(n_1372),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1327),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_SL g1482 ( 
.A(n_1350),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1305),
.B(n_1310),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1427),
.A2(n_1391),
.B1(n_1367),
.B2(n_1340),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1386),
.A2(n_1369),
.B(n_1413),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1397),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1403),
.Y(n_1487)
);

BUFx2_ASAP7_75t_R g1488 ( 
.A(n_1348),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1315),
.A2(n_1320),
.B(n_1422),
.Y(n_1489)
);

CKINVDCx8_ASAP7_75t_R g1490 ( 
.A(n_1303),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1345),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1399),
.A2(n_1320),
.B(n_1315),
.Y(n_1492)
);

BUFx2_ASAP7_75t_SL g1493 ( 
.A(n_1345),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1364),
.B(n_1353),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1387),
.A2(n_1363),
.B(n_1412),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1332),
.B(n_1349),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1355),
.B(n_1394),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1341),
.A2(n_1404),
.B1(n_1324),
.B2(n_1325),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1345),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1378),
.A2(n_1381),
.B1(n_1375),
.B2(n_1347),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1357),
.A2(n_1421),
.B(n_1430),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1351),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1421),
.A2(n_1352),
.B(n_1375),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1325),
.B(n_1356),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1374),
.B(n_1370),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1388),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_SL g1507 ( 
.A(n_1370),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1410),
.A2(n_1387),
.B1(n_1368),
.B2(n_1406),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1415),
.B(n_1388),
.Y(n_1509)
);

CKINVDCx6p67_ASAP7_75t_R g1510 ( 
.A(n_1388),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1343),
.B(n_1433),
.Y(n_1511)
);

INVx4_ASAP7_75t_L g1512 ( 
.A(n_1343),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1407),
.A2(n_1418),
.B(n_1384),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1407),
.A2(n_1418),
.B(n_1384),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1380),
.A2(n_1376),
.B(n_1433),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1316),
.B(n_1424),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1345),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1425),
.B(n_869),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1331),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1316),
.B(n_1424),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1328),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1342),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1367),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1432),
.A2(n_869),
.B1(n_893),
.B2(n_1091),
.Y(n_1524)
);

NAND2x1p5_ASAP7_75t_L g1525 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1525)
);

CKINVDCx16_ASAP7_75t_R g1526 ( 
.A(n_1379),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1527)
);

NOR2xp67_ASAP7_75t_L g1528 ( 
.A(n_1317),
.B(n_974),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1425),
.B(n_869),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1328),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1339),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1392),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1432),
.A2(n_869),
.B1(n_893),
.B2(n_1091),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1429),
.A2(n_869),
.B(n_893),
.C(n_888),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1316),
.B(n_1424),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1342),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1437),
.A2(n_869),
.B(n_893),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1437),
.B(n_869),
.C(n_893),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1425),
.Y(n_1539)
);

OAI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1366),
.A2(n_1035),
.B1(n_869),
.B2(n_1358),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1331),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1398),
.A2(n_1091),
.B1(n_1021),
.B2(n_1174),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1429),
.A2(n_1437),
.B1(n_1110),
.B2(n_1358),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1313),
.A2(n_893),
.B(n_1110),
.C(n_1437),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1429),
.A2(n_1437),
.B1(n_1110),
.B2(n_1358),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1326),
.A2(n_1402),
.B(n_1401),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1326),
.A2(n_1402),
.B(n_1401),
.Y(n_1547)
);

NAND2x1_ASAP7_75t_L g1548 ( 
.A(n_1316),
.B(n_1424),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1328),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1326),
.A2(n_1402),
.B(n_1401),
.Y(n_1550)
);

CKINVDCx11_ASAP7_75t_R g1551 ( 
.A(n_1392),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1367),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1425),
.B(n_869),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1328),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1328),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1437),
.A2(n_869),
.B(n_893),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1342),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_SL g1559 ( 
.A(n_1358),
.B(n_884),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1366),
.A2(n_1035),
.B1(n_869),
.B2(n_1358),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1437),
.A2(n_869),
.B(n_893),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1427),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1328),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1328),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_SL g1565 ( 
.A1(n_1333),
.A2(n_1298),
.B(n_1311),
.C(n_1359),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1331),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1342),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1317),
.B(n_974),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1306),
.A2(n_1428),
.B(n_1423),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1342),
.Y(n_1570)
);

A2O1A1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1313),
.A2(n_893),
.B(n_1110),
.C(n_1437),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1427),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1429),
.A2(n_1437),
.B1(n_1110),
.B2(n_1358),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1337),
.A2(n_1091),
.B1(n_1021),
.B2(n_893),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1331),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1306),
.A2(n_1428),
.B(n_1423),
.Y(n_1576)
);

BUFx8_ASAP7_75t_L g1577 ( 
.A(n_1398),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1337),
.A2(n_1091),
.B1(n_1021),
.B2(n_893),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1314),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1366),
.A2(n_1035),
.B1(n_869),
.B2(n_1358),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1316),
.B(n_1424),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1306),
.A2(n_1428),
.B(n_1423),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1432),
.B(n_1436),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1425),
.B(n_869),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1313),
.A2(n_893),
.B(n_1110),
.C(n_1437),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1432),
.B(n_1436),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1328),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1306),
.A2(n_1428),
.B(n_1423),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1425),
.B(n_869),
.Y(n_1589)
);

BUFx8_ASAP7_75t_L g1590 ( 
.A(n_1398),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1382),
.B(n_1425),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1548),
.B(n_1478),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1574),
.B(n_1578),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1544),
.A2(n_1585),
.B(n_1571),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1544),
.A2(n_1585),
.B(n_1571),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1472),
.A2(n_1543),
.B1(n_1573),
.B2(n_1545),
.Y(n_1596)
);

O2A1O1Ixp5_ASAP7_75t_L g1597 ( 
.A1(n_1447),
.A2(n_1540),
.B(n_1560),
.C(n_1580),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1579),
.B(n_1447),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1445),
.Y(n_1599)
);

BUFx4f_ASAP7_75t_L g1600 ( 
.A(n_1442),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1492),
.B(n_1545),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1481),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1456),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1486),
.A2(n_1460),
.B1(n_1573),
.B2(n_1470),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1591),
.B(n_1539),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1534),
.A2(n_1462),
.B(n_1560),
.C(n_1580),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1445),
.B(n_1459),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1497),
.B(n_1505),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1497),
.B(n_1496),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1537),
.B(n_1557),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1565),
.A2(n_1477),
.B(n_1561),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1458),
.A2(n_1515),
.B(n_1453),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1472),
.A2(n_1538),
.B1(n_1540),
.B2(n_1524),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1533),
.A2(n_1508),
.B1(n_1554),
.B2(n_1529),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1461),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1513),
.A2(n_1514),
.B(n_1503),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1508),
.A2(n_1589),
.B1(n_1529),
.B2(n_1584),
.Y(n_1617)
);

AOI221x1_ASAP7_75t_SL g1618 ( 
.A1(n_1468),
.A2(n_1554),
.B1(n_1589),
.B2(n_1518),
.C(n_1584),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1492),
.B(n_1483),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1477),
.A2(n_1480),
.B(n_1452),
.Y(n_1620)
);

CKINVDCx8_ASAP7_75t_R g1621 ( 
.A(n_1443),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1480),
.A2(n_1444),
.B(n_1446),
.C(n_1466),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1461),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1492),
.B(n_1519),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1502),
.Y(n_1625)
);

AOI21x1_ASAP7_75t_SL g1626 ( 
.A1(n_1583),
.A2(n_1586),
.B(n_1467),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1541),
.B(n_1566),
.Y(n_1627)
);

BUFx4f_ASAP7_75t_L g1628 ( 
.A(n_1442),
.Y(n_1628)
);

CKINVDCx8_ASAP7_75t_R g1629 ( 
.A(n_1443),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1523),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1518),
.B(n_1575),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1559),
.A2(n_1471),
.B(n_1500),
.C(n_1568),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1553),
.B(n_1484),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1549),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1474),
.B(n_1562),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1500),
.A2(n_1487),
.B1(n_1488),
.B2(n_1464),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1572),
.B(n_1450),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1487),
.A2(n_1464),
.B1(n_1507),
.B2(n_1490),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1457),
.B(n_1522),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1464),
.A2(n_1507),
.B1(n_1581),
.B2(n_1535),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1551),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1495),
.B(n_1475),
.Y(n_1643)
);

O2A1O1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1498),
.A2(n_1495),
.B(n_1465),
.C(n_1528),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1530),
.B(n_1555),
.Y(n_1645)
);

OAI31xp33_ASAP7_75t_L g1646 ( 
.A1(n_1455),
.A2(n_1527),
.A3(n_1525),
.B(n_1552),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1509),
.Y(n_1647)
);

OA22x2_ASAP7_75t_L g1648 ( 
.A1(n_1448),
.A2(n_1454),
.B1(n_1451),
.B2(n_1521),
.Y(n_1648)
);

AOI221x1_ASAP7_75t_SL g1649 ( 
.A1(n_1464),
.A2(n_1570),
.B1(n_1567),
.B2(n_1536),
.C(n_1558),
.Y(n_1649)
);

AOI21x1_ASAP7_75t_SL g1650 ( 
.A1(n_1511),
.A2(n_1449),
.B(n_1590),
.Y(n_1650)
);

CKINVDCx16_ASAP7_75t_R g1651 ( 
.A(n_1532),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1485),
.A2(n_1564),
.B1(n_1587),
.B2(n_1549),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1455),
.A2(n_1552),
.B(n_1494),
.C(n_1485),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1485),
.A2(n_1556),
.B1(n_1587),
.B2(n_1563),
.Y(n_1655)
);

AOI21x1_ASAP7_75t_SL g1656 ( 
.A1(n_1449),
.A2(n_1590),
.B(n_1577),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1449),
.B(n_1563),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1476),
.B(n_1491),
.Y(n_1658)
);

O2A1O1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1494),
.A2(n_1476),
.B(n_1463),
.C(n_1547),
.Y(n_1659)
);

AOI21x1_ASAP7_75t_SL g1660 ( 
.A1(n_1577),
.A2(n_1590),
.B(n_1482),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1494),
.A2(n_1547),
.B(n_1546),
.C(n_1550),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1482),
.A2(n_1510),
.B1(n_1512),
.B2(n_1526),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1577),
.B(n_1499),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1473),
.A2(n_1531),
.B1(n_1506),
.B2(n_1517),
.C(n_1493),
.Y(n_1664)
);

AND2x2_ASAP7_75t_SL g1665 ( 
.A(n_1546),
.B(n_1550),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1469),
.A2(n_1517),
.B1(n_1531),
.B2(n_1551),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1517),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1569),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1576),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1582),
.B(n_1588),
.Y(n_1670)
);

O2A1O1Ixp5_ASAP7_75t_L g1671 ( 
.A1(n_1478),
.A2(n_1373),
.B(n_1447),
.C(n_1540),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1579),
.B(n_1447),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1544),
.A2(n_1398),
.B(n_1571),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1574),
.A2(n_1578),
.B1(n_1542),
.B2(n_1189),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1481),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1516),
.B(n_1520),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1501),
.A2(n_1478),
.B(n_1479),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1445),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1472),
.A2(n_1366),
.B1(n_1545),
.B2(n_1543),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1461),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1501),
.A2(n_1478),
.B(n_1479),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1544),
.A2(n_1398),
.B(n_1571),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1579),
.B(n_1447),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1445),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_SL g1685 ( 
.A1(n_1574),
.A2(n_1578),
.B1(n_1542),
.B2(n_1189),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1591),
.B(n_1539),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1472),
.A2(n_1366),
.B1(n_1545),
.B2(n_1543),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1461),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1579),
.B(n_1447),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1472),
.A2(n_1366),
.B1(n_1545),
.B2(n_1543),
.Y(n_1690)
);

OR2x6_ASAP7_75t_L g1691 ( 
.A(n_1548),
.B(n_1424),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1579),
.A2(n_1489),
.B(n_1565),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1445),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1472),
.A2(n_1366),
.B1(n_1545),
.B2(n_1543),
.Y(n_1694)
);

O2A1O1Ixp5_ASAP7_75t_L g1695 ( 
.A1(n_1478),
.A2(n_1373),
.B(n_1447),
.C(n_1540),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1544),
.A2(n_1398),
.B(n_1571),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1472),
.A2(n_1366),
.B1(n_1545),
.B2(n_1543),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1591),
.B(n_1539),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1579),
.A2(n_1489),
.B(n_1565),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1461),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1544),
.A2(n_1398),
.B(n_1571),
.Y(n_1701)
);

AO21x1_ASAP7_75t_SL g1702 ( 
.A1(n_1643),
.A2(n_1653),
.B(n_1598),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1624),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1608),
.B(n_1609),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1616),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1619),
.B(n_1624),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_R g1707 ( 
.A(n_1642),
.B(n_1621),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1669),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1592),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1619),
.B(n_1601),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1601),
.B(n_1653),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1598),
.B(n_1672),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1692),
.A2(n_1699),
.B(n_1620),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1592),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1672),
.B(n_1683),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1674),
.A2(n_1685),
.B1(n_1694),
.B2(n_1687),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1615),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1599),
.B(n_1678),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1689),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1623),
.Y(n_1720)
);

AO21x2_ASAP7_75t_L g1721 ( 
.A1(n_1670),
.A2(n_1661),
.B(n_1611),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1671),
.A2(n_1695),
.B(n_1597),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1659),
.B(n_1654),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1677),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1606),
.A2(n_1613),
.B1(n_1614),
.B2(n_1617),
.C(n_1618),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1633),
.B(n_1688),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1680),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1677),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1681),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1684),
.B(n_1693),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1625),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1647),
.B(n_1610),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1612),
.Y(n_1735)
);

AOI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1655),
.A2(n_1652),
.B(n_1668),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1700),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1592),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1648),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1648),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1665),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1691),
.Y(n_1742)
);

OR2x2_ASAP7_75t_SL g1743 ( 
.A(n_1651),
.B(n_1637),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1593),
.A2(n_1622),
.B1(n_1632),
.B2(n_1682),
.C(n_1673),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1649),
.Y(n_1745)
);

AO21x1_ASAP7_75t_SL g1746 ( 
.A1(n_1635),
.A2(n_1627),
.B(n_1631),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1649),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1676),
.B(n_1691),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1630),
.Y(n_1749)
);

INVx4_ASAP7_75t_L g1750 ( 
.A(n_1691),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1644),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1676),
.B(n_1638),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1607),
.B(n_1605),
.Y(n_1753)
);

AO21x2_ASAP7_75t_L g1754 ( 
.A1(n_1655),
.A2(n_1652),
.B(n_1596),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1686),
.B(n_1698),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1638),
.B(n_1641),
.Y(n_1756)
);

NOR3xp33_ASAP7_75t_L g1757 ( 
.A(n_1604),
.B(n_1687),
.C(n_1679),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1639),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1645),
.Y(n_1759)
);

AO21x2_ASAP7_75t_L g1760 ( 
.A1(n_1690),
.A2(n_1697),
.B(n_1694),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1636),
.B(n_1603),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1696),
.B(n_1701),
.Y(n_1762)
);

AO21x2_ASAP7_75t_L g1763 ( 
.A1(n_1690),
.A2(n_1697),
.B(n_1636),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1627),
.B(n_1640),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1618),
.B(n_1634),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1708),
.Y(n_1767)
);

INVxp67_ASAP7_75t_SL g1768 ( 
.A(n_1705),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1710),
.B(n_1667),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1710),
.B(n_1706),
.Y(n_1770)
);

OAI222xp33_ASAP7_75t_L g1771 ( 
.A1(n_1716),
.A2(n_1722),
.B1(n_1744),
.B2(n_1713),
.C1(n_1756),
.C2(n_1761),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1741),
.B(n_1711),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1703),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_SL g1774 ( 
.A(n_1746),
.B(n_1666),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1703),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1717),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1711),
.B(n_1657),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1705),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1716),
.B(n_1646),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_SL g1780 ( 
.A(n_1746),
.B(n_1666),
.Y(n_1780)
);

INVx6_ASAP7_75t_L g1781 ( 
.A(n_1750),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1735),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1757),
.A2(n_1664),
.B1(n_1628),
.B2(n_1600),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1750),
.B(n_1658),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1702),
.B(n_1675),
.Y(n_1785)
);

OAI21xp33_ASAP7_75t_L g1786 ( 
.A1(n_1726),
.A2(n_1662),
.B(n_1663),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1735),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1709),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1722),
.B(n_1662),
.C(n_1602),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1720),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1733),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1719),
.B(n_1626),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1719),
.B(n_1629),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1712),
.B(n_1715),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1709),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1722),
.A2(n_1656),
.B1(n_1660),
.B2(n_1650),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1709),
.B(n_1724),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1728),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1715),
.B(n_1727),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1737),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1764),
.B(n_1734),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1750),
.B(n_1748),
.Y(n_1802)
);

AOI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1760),
.A2(n_1763),
.B1(n_1751),
.B2(n_1765),
.C(n_1732),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1758),
.B(n_1754),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1779),
.A2(n_1722),
.B(n_1760),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1803),
.B(n_1722),
.C(n_1723),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1790),
.Y(n_1807)
);

OAI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1803),
.A2(n_1723),
.B1(n_1762),
.B2(n_1724),
.C(n_1739),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1772),
.B(n_1714),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1771),
.A2(n_1760),
.B1(n_1763),
.B2(n_1718),
.C(n_1749),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1767),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1795),
.Y(n_1812)
);

NOR2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1789),
.B(n_1756),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1786),
.A2(n_1763),
.B1(n_1723),
.B2(n_1762),
.Y(n_1814)
);

NAND2xp33_ASAP7_75t_R g1815 ( 
.A(n_1766),
.B(n_1707),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1789),
.A2(n_1743),
.B1(n_1762),
.B2(n_1761),
.Y(n_1816)
);

OAI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1786),
.A2(n_1723),
.B1(n_1762),
.B2(n_1724),
.C(n_1739),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1790),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1801),
.B(n_1759),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1798),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1772),
.B(n_1714),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1777),
.B(n_1738),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1777),
.B(n_1738),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1792),
.A2(n_1740),
.B(n_1736),
.C(n_1747),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1783),
.A2(n_1762),
.B1(n_1724),
.B2(n_1740),
.C(n_1755),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1783),
.Y(n_1826)
);

CKINVDCx16_ASAP7_75t_R g1827 ( 
.A(n_1784),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1797),
.A2(n_1743),
.B1(n_1709),
.B2(n_1724),
.Y(n_1828)
);

OA21x2_ASAP7_75t_L g1829 ( 
.A1(n_1768),
.A2(n_1725),
.B(n_1731),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1782),
.Y(n_1830)
);

NAND2x1_ASAP7_75t_L g1831 ( 
.A(n_1781),
.B(n_1709),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1804),
.B(n_1754),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1778),
.A2(n_1729),
.B(n_1725),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1794),
.B(n_1755),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1798),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1804),
.B(n_1754),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1800),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1800),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1788),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1773),
.Y(n_1840)
);

OAI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1792),
.A2(n_1736),
.B(n_1745),
.C(n_1747),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1793),
.A2(n_1752),
.B1(n_1748),
.B2(n_1704),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1769),
.B(n_1758),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1797),
.A2(n_1748),
.B1(n_1752),
.B2(n_1758),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1801),
.B(n_1753),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1776),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1791),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1769),
.B(n_1721),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1799),
.B(n_1721),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_1812),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1812),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1827),
.Y(n_1852)
);

OA21x2_ASAP7_75t_L g1853 ( 
.A1(n_1806),
.A2(n_1730),
.B(n_1729),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1847),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1847),
.Y(n_1855)
);

INVx3_ASAP7_75t_L g1856 ( 
.A(n_1829),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1840),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1832),
.B(n_1836),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1812),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1848),
.B(n_1770),
.Y(n_1860)
);

BUFx8_ASAP7_75t_L g1861 ( 
.A(n_1824),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1848),
.B(n_1807),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1833),
.Y(n_1863)
);

OR2x6_ASAP7_75t_L g1864 ( 
.A(n_1805),
.B(n_1797),
.Y(n_1864)
);

OR2x6_ASAP7_75t_L g1865 ( 
.A(n_1831),
.B(n_1797),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1837),
.B(n_1773),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1810),
.B(n_1797),
.C(n_1796),
.Y(n_1867)
);

NOR2x1_ASAP7_75t_L g1868 ( 
.A(n_1813),
.B(n_1787),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1812),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1838),
.B(n_1775),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1811),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1818),
.B(n_1775),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1808),
.A2(n_1771),
.B(n_1796),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1839),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1831),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1818),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1839),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1852),
.B(n_1827),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1852),
.B(n_1826),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1875),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1854),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1868),
.B(n_1813),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1862),
.B(n_1849),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1868),
.B(n_1830),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1865),
.B(n_1822),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1857),
.B(n_1841),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1854),
.Y(n_1887)
);

INVx4_ASAP7_75t_L g1888 ( 
.A(n_1875),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1855),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1855),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1865),
.B(n_1802),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1865),
.B(n_1864),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1856),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1875),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1864),
.B(n_1823),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1860),
.B(n_1820),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1875),
.B(n_1802),
.Y(n_1897)
);

NAND2x1p5_ASAP7_75t_L g1898 ( 
.A(n_1875),
.B(n_1795),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1856),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1864),
.B(n_1809),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1864),
.B(n_1809),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1864),
.B(n_1821),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1864),
.B(n_1821),
.Y(n_1903)
);

NAND2xp33_ASAP7_75t_SL g1904 ( 
.A(n_1875),
.B(n_1826),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1858),
.B(n_1774),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1860),
.B(n_1820),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1858),
.B(n_1774),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1867),
.B(n_1846),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1858),
.B(n_1780),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1875),
.B(n_1780),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1871),
.Y(n_1911)
);

AND2x4_ASAP7_75t_SL g1912 ( 
.A(n_1857),
.B(n_1785),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1866),
.B(n_1835),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1856),
.Y(n_1914)
);

NOR2x1_ASAP7_75t_R g1915 ( 
.A(n_1861),
.B(n_1846),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1850),
.B(n_1843),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1886),
.B(n_1866),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1882),
.B(n_1850),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1882),
.B(n_1853),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1879),
.B(n_1874),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1893),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1881),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1893),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1881),
.Y(n_1924)
);

NOR2xp67_ASAP7_75t_SL g1925 ( 
.A(n_1888),
.B(n_1867),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1878),
.B(n_1850),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1879),
.B(n_1874),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1886),
.B(n_1870),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1908),
.B(n_1834),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1878),
.B(n_1869),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1915),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1888),
.B(n_1851),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1908),
.B(n_1825),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1910),
.B(n_1869),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1887),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1887),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1888),
.B(n_1869),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1904),
.Y(n_1938)
);

NAND2xp67_ASAP7_75t_L g1939 ( 
.A(n_1910),
.B(n_1793),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1896),
.B(n_1870),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1905),
.B(n_1851),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1889),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1889),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1890),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1915),
.B(n_1845),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1905),
.B(n_1851),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1893),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1916),
.B(n_1819),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1899),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1907),
.B(n_1859),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1913),
.A2(n_1873),
.B1(n_1817),
.B2(n_1814),
.C(n_1816),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1896),
.B(n_1872),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1890),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1916),
.Y(n_1954)
);

OR2x6_ASAP7_75t_L g1955 ( 
.A(n_1888),
.B(n_1873),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1907),
.B(n_1859),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1912),
.Y(n_1957)
);

NAND2x1_ASAP7_75t_SL g1958 ( 
.A(n_1880),
.B(n_1853),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1884),
.Y(n_1959)
);

OAI32xp33_ASAP7_75t_L g1960 ( 
.A1(n_1898),
.A2(n_1877),
.A3(n_1876),
.B1(n_1815),
.B2(n_1828),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1933),
.A2(n_1861),
.B1(n_1892),
.B2(n_1891),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1922),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1924),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1937),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1926),
.B(n_1909),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1918),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1954),
.B(n_1913),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1919),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1926),
.B(n_1909),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1932),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1935),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1929),
.B(n_1877),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1930),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1931),
.B(n_1885),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1936),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1930),
.B(n_1897),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1942),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1951),
.A2(n_1912),
.B1(n_1844),
.B2(n_1842),
.Y(n_1978)
);

INVx3_ASAP7_75t_SL g1979 ( 
.A(n_1955),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1943),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1948),
.B(n_1906),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1945),
.B(n_1939),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1944),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1917),
.B(n_1906),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1934),
.B(n_1897),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1917),
.B(n_1883),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1934),
.B(n_1897),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1941),
.B(n_1897),
.Y(n_1988)
);

CKINVDCx16_ASAP7_75t_R g1989 ( 
.A(n_1931),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1941),
.B(n_1885),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1973),
.B(n_1989),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1962),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1989),
.B(n_1938),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1979),
.A2(n_1955),
.B1(n_1920),
.B2(n_1927),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1984),
.B(n_1928),
.Y(n_1995)
);

OAI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1974),
.A2(n_1925),
.B(n_1939),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1976),
.B(n_1955),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1970),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1976),
.B(n_1955),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1972),
.A2(n_1925),
.B1(n_1861),
.B2(n_1928),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1970),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1962),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1964),
.B(n_1957),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1984),
.B(n_1940),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1986),
.B(n_1940),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1963),
.Y(n_2006)
);

AOI222xp33_ASAP7_75t_L g2007 ( 
.A1(n_1978),
.A2(n_1960),
.B1(n_1861),
.B2(n_1918),
.C1(n_1892),
.C2(n_1957),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1961),
.A2(n_1919),
.B(n_1946),
.Y(n_2008)
);

NOR2x1_ASAP7_75t_L g2009 ( 
.A(n_1964),
.B(n_1880),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1963),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1968),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1982),
.A2(n_1919),
.B(n_1932),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1971),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1985),
.B(n_1946),
.Y(n_2014)
);

AOI322xp5_ASAP7_75t_L g2015 ( 
.A1(n_1966),
.A2(n_1863),
.A3(n_1900),
.B1(n_1903),
.B2(n_1901),
.C1(n_1902),
.C2(n_1895),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1993),
.A2(n_1979),
.B1(n_1981),
.B2(n_1966),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2001),
.B(n_1985),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1995),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_2014),
.B(n_1987),
.Y(n_2019)
);

NAND2xp33_ASAP7_75t_L g2020 ( 
.A(n_2000),
.B(n_1979),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2001),
.B(n_1987),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1998),
.Y(n_2022)
);

INVx1_ASAP7_75t_SL g2023 ( 
.A(n_1991),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_2005),
.B(n_1967),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_2004),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_2000),
.B(n_1968),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_2003),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1993),
.A2(n_1988),
.B1(n_1990),
.B2(n_1861),
.Y(n_2028)
);

NOR2x1_ASAP7_75t_L g2029 ( 
.A(n_2011),
.B(n_1971),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_2016),
.A2(n_2008),
.B1(n_1994),
.B2(n_1996),
.Y(n_2030)
);

OAI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_2016),
.A2(n_2007),
.B1(n_2012),
.B2(n_2015),
.C(n_1999),
.Y(n_2031)
);

AOI221xp5_ASAP7_75t_L g2032 ( 
.A1(n_2026),
.A2(n_1994),
.B1(n_1998),
.B2(n_2003),
.C(n_1992),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2027),
.B(n_2003),
.Y(n_2033)
);

OR2x6_ASAP7_75t_L g2034 ( 
.A(n_2017),
.B(n_1997),
.Y(n_2034)
);

OAI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_2023),
.A2(n_1988),
.B(n_1990),
.Y(n_2035)
);

NOR3x1_ASAP7_75t_L g2036 ( 
.A(n_2021),
.B(n_2006),
.C(n_2002),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_2026),
.A2(n_2009),
.B(n_2011),
.Y(n_2037)
);

OAI211xp5_ASAP7_75t_L g2038 ( 
.A1(n_2029),
.A2(n_2013),
.B(n_2010),
.C(n_1975),
.Y(n_2038)
);

O2A1O1Ixp5_ASAP7_75t_L g2039 ( 
.A1(n_2022),
.A2(n_1959),
.B(n_1880),
.C(n_1894),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_2020),
.A2(n_1965),
.B1(n_1969),
.B2(n_1932),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2025),
.A2(n_1975),
.B1(n_1983),
.B2(n_1980),
.C(n_1977),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2030),
.A2(n_2019),
.B1(n_2028),
.B2(n_2018),
.Y(n_2042)
);

XOR2x2_ASAP7_75t_L g2043 ( 
.A(n_2031),
.B(n_2024),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2033),
.Y(n_2044)
);

INVxp67_ASAP7_75t_L g2045 ( 
.A(n_2034),
.Y(n_2045)
);

NOR2x1_ASAP7_75t_L g2046 ( 
.A(n_2038),
.B(n_1977),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2032),
.A2(n_1969),
.B1(n_1965),
.B2(n_1894),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2040),
.A2(n_1986),
.B1(n_1952),
.B2(n_1898),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2046),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_2043),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2044),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_2045),
.B(n_2037),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2047),
.B(n_2036),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2042),
.B(n_2035),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2048),
.B(n_2041),
.Y(n_2055)
);

OAI32xp33_ASAP7_75t_L g2056 ( 
.A1(n_2045),
.A2(n_1983),
.A3(n_1980),
.B1(n_1959),
.B2(n_1880),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2052),
.B(n_1950),
.Y(n_2057)
);

XOR2x2_ASAP7_75t_L g2058 ( 
.A(n_2054),
.B(n_1898),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2050),
.B(n_1950),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2050),
.A2(n_2039),
.B(n_1953),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2049),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_2050),
.B(n_1894),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_R g2063 ( 
.A(n_2051),
.B(n_2053),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_L g2064 ( 
.A(n_2062),
.B(n_2052),
.C(n_2053),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_SL g2065 ( 
.A(n_2059),
.B(n_2056),
.C(n_2055),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2057),
.B(n_1956),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_2058),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_R g2068 ( 
.A(n_2061),
.B(n_1894),
.Y(n_2068)
);

NOR3xp33_ASAP7_75t_L g2069 ( 
.A(n_2064),
.B(n_2063),
.C(n_2060),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2066),
.B(n_1959),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2067),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_2070),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2069),
.B(n_2065),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2072),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2073),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2072),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_2074),
.B(n_2071),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2076),
.A2(n_2068),
.B(n_1923),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2075),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_SL g2080 ( 
.A1(n_2077),
.A2(n_1952),
.B1(n_1921),
.B2(n_1947),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_SL g2081 ( 
.A1(n_2080),
.A2(n_2079),
.B1(n_2078),
.B2(n_1921),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_2081),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_2082),
.A2(n_1923),
.B1(n_1947),
.B2(n_1949),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2083),
.A2(n_1949),
.B(n_1958),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_2084),
.A2(n_1899),
.B1(n_1914),
.B2(n_1956),
.Y(n_2085)
);

AOI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2085),
.A2(n_1899),
.B(n_1914),
.C(n_1911),
.Y(n_2086)
);


endmodule