module fake_jpeg_20439_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_1),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_3),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_68),
.B1(n_40),
.B2(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_3),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_73),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_41),
.B1(n_42),
.B2(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_48),
.B1(n_45),
.B2(n_52),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_51),
.B1(n_62),
.B2(n_54),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_78),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_79),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_75),
.B1(n_56),
.B2(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_53),
.C(n_44),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_102),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_56),
.B1(n_59),
.B2(n_5),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_92),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_96),
.B1(n_93),
.B2(n_97),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_6),
.B(n_7),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_105),
.C(n_108),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_113),
.B(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_114),
.B1(n_16),
.B2(n_17),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_15),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_114),
.C(n_34),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_37),
.Y(n_124)
);


endmodule