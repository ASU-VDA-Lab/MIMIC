module fake_jpeg_31108_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_46),
.B1(n_37),
.B2(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_63),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_21),
.B1(n_32),
.B2(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_41),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_45),
.B(n_48),
.Y(n_68)
);

OR2x4_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_78),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_19),
.B1(n_36),
.B2(n_33),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_3),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_18),
.B1(n_30),
.B2(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_89),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_62),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_87),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_14),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_5),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_70),
.B1(n_71),
.B2(n_7),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_82),
.A3(n_6),
.B1(n_13),
.B2(n_17),
.C(n_25),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_95),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_22),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_83),
.C(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_99),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_94),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_101),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_91),
.C(n_100),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_94),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_10),
.C(n_27),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_28),
.Y(n_106)
);


endmodule