module fake_jpeg_27592_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_44),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_74),
.B1(n_49),
.B2(n_36),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_27),
.B1(n_35),
.B2(n_16),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_25),
.B1(n_16),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_67),
.Y(n_83)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_61),
.Y(n_105)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_20),
.B1(n_22),
.B2(n_19),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_22),
.B1(n_20),
.B2(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_85),
.Y(n_135)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_82),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_49),
.B1(n_36),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_44),
.B1(n_53),
.B2(n_40),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_28),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_93),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_22),
.B1(n_21),
.B2(n_34),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_120)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_19),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_106),
.Y(n_122)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_114),
.Y(n_134)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_59),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_37),
.Y(n_145)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_33),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_10),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_125),
.B1(n_144),
.B2(n_105),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_44),
.B1(n_28),
.B2(n_21),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_119),
.A2(n_113),
.B1(n_86),
.B2(n_91),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_143),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_39),
.B1(n_38),
.B2(n_42),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_110),
.B(n_25),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_39),
.C(n_38),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_82),
.C(n_96),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_39),
.B1(n_26),
.B2(n_34),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_122),
.B1(n_134),
.B2(n_135),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_78),
.B(n_101),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_29),
.B(n_77),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_154),
.B(n_155),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_41),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_150),
.B(n_157),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_158),
.B1(n_166),
.B2(n_168),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_142),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_105),
.B(n_41),
.C(n_42),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_25),
.B(n_1),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_162),
.B(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_120),
.B1(n_124),
.B2(n_125),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_41),
.C(n_89),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_136),
.B(n_123),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_0),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_169),
.B1(n_167),
.B2(n_178),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_2),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_167),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_91),
.B(n_89),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_3),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_37),
.B1(n_109),
.B2(n_12),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_9),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_9),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_15),
.C(n_14),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_14),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_178),
.B(n_4),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_4),
.B(n_5),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_127),
.B1(n_136),
.B2(n_130),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_187),
.B(n_190),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_142),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_139),
.B1(n_133),
.B2(n_130),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_200),
.B1(n_202),
.B2(n_205),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_12),
.C(n_13),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_139),
.B1(n_133),
.B2(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_177),
.B(n_159),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_136),
.B1(n_140),
.B2(n_123),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_155),
.C(n_146),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_12),
.B1(n_13),
.B2(n_8),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_5),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_156),
.Y(n_213)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_214),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_154),
.C(n_162),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_227),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_154),
.C(n_163),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_154),
.C(n_163),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_180),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_154),
.B1(n_176),
.B2(n_169),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_238),
.B(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_239),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_203),
.B1(n_199),
.B2(n_184),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_183),
.B1(n_189),
.B2(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_252),
.B1(n_257),
.B2(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_237),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_254),
.B(n_210),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_219),
.B1(n_235),
.B2(n_227),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_192),
.B(n_206),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_262),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_183),
.B1(n_195),
.B2(n_204),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_212),
.A2(n_148),
.B1(n_182),
.B2(n_192),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_181),
.B1(n_182),
.B2(n_179),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_236),
.B1(n_232),
.B2(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_179),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_215),
.C(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_267),
.C(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_271),
.B1(n_279),
.B2(n_245),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_215),
.C(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_241),
.B(n_237),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_243),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_240),
.B1(n_241),
.B2(n_248),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_213),
.C(n_218),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_252),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_247),
.A2(n_214),
.B1(n_226),
.B2(n_208),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_249),
.B(n_256),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_201),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_287),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_271),
.Y(n_302)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_245),
.B(n_250),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_292),
.A2(n_293),
.B(n_284),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_251),
.C(n_257),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_211),
.C(n_7),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_277),
.C(n_279),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_5),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_272),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_264),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_306),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_302),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_284),
.B1(n_286),
.B2(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_282),
.C(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_268),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_273),
.B1(n_290),
.B2(n_269),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_319),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_306),
.C(n_307),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_266),
.C(n_274),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_290),
.B1(n_269),
.B2(n_270),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_303),
.B1(n_300),
.B2(n_308),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_309),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_325),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_274),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_317),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_320),
.B1(n_314),
.B2(n_319),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_328),
.B(n_324),
.Y(n_334)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.A3(n_318),
.B1(n_325),
.B2(n_331),
.C(n_326),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_268),
.B(n_7),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_7),
.B(n_8),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_7),
.C(n_8),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);


endmodule