module fake_jpeg_23486_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_18),
.B(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.C(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_20),
.B1(n_25),
.B2(n_23),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_15),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_57),
.B1(n_17),
.B2(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_56),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_59),
.B(n_49),
.C(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_21),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_48),
.B1(n_42),
.B2(n_44),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_71),
.Y(n_94)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_45),
.B1(n_41),
.B2(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_31),
.B1(n_48),
.B2(n_34),
.Y(n_91)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_73),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_42),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_58),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_R g92 ( 
.A(n_78),
.B(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_70),
.C(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_84),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_85),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_29),
.B1(n_34),
.B2(n_24),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_96),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_96),
.B1(n_89),
.B2(n_85),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_95),
.Y(n_101)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_2),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_73),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_104),
.B1(n_90),
.B2(n_87),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_69),
.B1(n_77),
.B2(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_R g133 ( 
.A(n_116),
.B(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_126),
.B1(n_130),
.B2(n_118),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_134),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_84),
.B1(n_67),
.B2(n_95),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_95),
.B1(n_72),
.B2(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_74),
.C(n_117),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_101),
.B1(n_112),
.B2(n_114),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_141),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_101),
.A3(n_108),
.B1(n_112),
.B2(n_116),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_130),
.Y(n_155)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_133),
.B1(n_122),
.B2(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_120),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_125),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_37),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_135),
.C(n_121),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_39),
.Y(n_174)
);

AOI321xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_116),
.A3(n_127),
.B1(n_65),
.B2(n_114),
.C(n_86),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_143),
.B(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

AOI321xp33_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_176),
.A3(n_161),
.B1(n_160),
.B2(n_162),
.C(n_37),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_161),
.A2(n_147),
.B1(n_150),
.B2(n_141),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_51),
.B1(n_37),
.B2(n_33),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_155),
.C(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_129),
.B1(n_51),
.B2(n_30),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_51),
.B1(n_33),
.B2(n_5),
.Y(n_181)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_181),
.C(n_33),
.Y(n_190)
);

AOI31xp67_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_183),
.A3(n_4),
.B(n_6),
.Y(n_189)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_167),
.B(n_168),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_184),
.B(n_176),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_3),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_171),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_191),
.C(n_7),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_189),
.B1(n_14),
.B2(n_7),
.Y(n_194)
);

NAND4xp25_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_170),
.C(n_171),
.D(n_10),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_190),
.B(n_7),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_9),
.C(n_13),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_183),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_193),
.B(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_14),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_8),
.B(n_185),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_192),
.B(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_198),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_8),
.Y(n_204)
);


endmodule