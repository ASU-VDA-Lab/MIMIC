module real_jpeg_27650_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_244;
wire n_295;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_0),
.B(n_51),
.Y(n_82)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_0),
.B(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_0),
.B(n_228),
.Y(n_233)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_4),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_30),
.B1(n_43),
.B2(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_30),
.B1(n_49),
.B2(n_51),
.Y(n_120)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_4),
.A2(n_6),
.B1(n_29),
.B2(n_65),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_5),
.B1(n_29),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_5),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_134),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_5),
.A2(n_43),
.B1(n_47),
.B2(n_134),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_5),
.A2(n_49),
.B1(n_51),
.B2(n_134),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_43),
.B1(n_47),
.B2(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_49),
.B1(n_51),
.B2(n_65),
.Y(n_149)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_7),
.A2(n_10),
.B(n_49),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_9),
.A2(n_10),
.B(n_43),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_29),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_43),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_49),
.B1(n_51),
.B2(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_21),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_10),
.B(n_60),
.Y(n_223)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_109),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_108),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_90),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_16),
.B(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_69),
.C(n_77),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_17),
.B(n_69),
.CI(n_77),
.CON(n_140),
.SN(n_140)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_37),
.B2(n_38),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_18),
.A2(n_19),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_56),
.C(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_20),
.B(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_21),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_23),
.B(n_29),
.C(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_22),
.A2(n_33),
.B(n_35),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_22),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_24),
.B(n_26),
.Y(n_170)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_25),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_25),
.B(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_55),
.B(n_61),
.C(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_28),
.B(n_33),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_32),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_34),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_35),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_36),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_56),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_39),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_39),
.A2(n_107),
.B1(n_156),
.B2(n_157),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_52),
.B(n_53),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_41),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_41),
.B(n_54),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_41),
.B(n_201),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_43),
.A2(n_45),
.B(n_55),
.C(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_48),
.B(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_51),
.B(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_52),
.A2(n_75),
.B(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_52),
.B(n_55),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_55),
.B(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B(n_66),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_57),
.B(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_57),
.B(n_159),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_57),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_60),
.B(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_67),
.B(n_167),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_69),
.A2(n_70),
.B(n_73),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_71),
.A2(n_102),
.B(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_72),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_74),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_75),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_89),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_78),
.A2(n_79),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_81),
.B1(n_89),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_80),
.A2(n_81),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_81),
.B(n_193),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_82),
.B(n_85),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_82),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_85),
.Y(n_116)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx5_ASAP7_75t_SL g244 ( 
.A(n_83),
.Y(n_244)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_86),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_88),
.B(n_210),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_89),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_106),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_105),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_97),
.B(n_155),
.Y(n_272)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_101),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_154),
.C(n_156),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_141),
.B(n_298),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_140),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_111),
.B(n_140),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_135),
.C(n_136),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_112),
.A2(n_113),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_123),
.C(n_126),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_114),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_115),
.B(n_122),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_116),
.B(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_117),
.A2(n_149),
.B(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_118),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_123),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_125),
.B(n_158),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_135),
.B(n_136),
.Y(n_296)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_140),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_292),
.B(n_297),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_279),
.B(n_291),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_187),
.B(n_262),
.C(n_278),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_175),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_145),
.B(n_175),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_160),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_147),
.B(n_153),
.C(n_160),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_148),
.B(n_151),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_150),
.B(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_152),
.B(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_162),
.B(n_165),
.C(n_168),
.Y(n_276)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_176),
.A2(n_177),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.C(n_185),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_185),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_233),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_261),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_254),
.B(n_260),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_212),
.B(n_253),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_202),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_191),
.B(n_202),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.C(n_198),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_192),
.B(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_209),
.C(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_248),
.B(n_252),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_229),
.B(n_247),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_220),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_236),
.B(n_246),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_240),
.B(n_245),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_276),
.B2(n_277),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_268),
.C(n_277),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_287),
.B2(n_288),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_288),
.C(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);


endmodule