module fake_ariane_1206_n_1808 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1808);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1808;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_73),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_9),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_0),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_60),
.Y(n_182)
);

BUFx8_ASAP7_75t_SL g183 ( 
.A(n_20),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_78),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_32),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_35),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_75),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_36),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_54),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_98),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_57),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_48),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_139),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_80),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_71),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_42),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_11),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_109),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_165),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_135),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_13),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_74),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_105),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_43),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_20),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_56),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_52),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_83),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_62),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_81),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_11),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_65),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_24),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_140),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_29),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_70),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_16),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_50),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_35),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_119),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_91),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_51),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_52),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_112),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_25),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_15),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_101),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_133),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_28),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_126),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_29),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_47),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_158),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_55),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_31),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_94),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_8),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_124),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_160),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_53),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_168),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_100),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_14),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_14),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_36),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_79),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_68),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_162),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_12),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_87),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_143),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_147),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_44),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_113),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_103),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_61),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_39),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_39),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_41),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_82),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_131),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_167),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_46),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_108),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_93),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_23),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_21),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_59),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_156),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_115),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_17),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_49),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_7),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_2),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_10),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_26),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_63),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_159),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_85),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_3),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_95),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_148),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_30),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_22),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_50),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_187),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_203),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_214),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_175),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_314),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_183),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_268),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_268),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_300),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_264),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_268),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_181),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_181),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_243),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_263),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_263),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_308),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_224),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_307),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_218),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_218),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_276),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_184),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_180),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_249),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_270),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_216),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_217),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_257),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_180),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_264),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_302),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_184),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_275),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_175),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_319),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_289),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_284),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_180),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_270),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_284),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_284),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_176),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_171),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_312),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_335),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_331),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_189),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_192),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_196),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_190),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_204),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_205),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_171),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_209),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_272),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_173),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_213),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_229),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_178),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_232),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_272),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_272),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_260),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_347),
.B(n_309),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_415),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_283),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_409),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_341),
.A2(n_252),
.B1(n_245),
.B2(n_316),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_372),
.B(n_173),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_343),
.A2(n_348),
.B(n_366),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_362),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_173),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

OAI22x1_ASAP7_75t_SL g445 ( 
.A1(n_346),
.A2(n_324),
.B1(n_317),
.B2(n_225),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_365),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_283),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_373),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_195),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_398),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_239),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_398),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_399),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_399),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_353),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_390),
.B(n_242),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_405),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_402),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_380),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_408),
.A2(n_255),
.B(n_244),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_355),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_408),
.B(n_178),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_355),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_357),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_182),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_384),
.Y(n_483)
);

INVx6_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_416),
.B(n_262),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_357),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_419),
.B(n_265),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_358),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_356),
.B(n_182),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_406),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_358),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_393),
.B(n_359),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_351),
.Y(n_495)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_364),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_388),
.B(n_271),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_337),
.A2(n_286),
.B(n_277),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_338),
.B(n_303),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_439),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

NAND2x1p5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_475),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_SL g507 ( 
.A1(n_429),
.A2(n_379),
.B(n_350),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

NOR2x1p5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_346),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_433),
.B(n_397),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_496),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_467),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_497),
.A2(n_361),
.B1(n_354),
.B2(n_432),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_467),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_467),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_438),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_482),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_460),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_460),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_484),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_467),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_496),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_441),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_460),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_460),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_494),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_460),
.Y(n_533)
);

AND2x2_ASAP7_75t_SL g534 ( 
.A(n_433),
.B(n_173),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_433),
.B(n_397),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_460),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_491),
.B(n_412),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_432),
.B(n_345),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_465),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_467),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_467),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_427),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_470),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_477),
.B(n_412),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_482),
.B(n_418),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_436),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_458),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_470),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_470),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_496),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_471),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_482),
.B(n_378),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_458),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_464),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_480),
.B(n_367),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_480),
.B(n_367),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_480),
.B(n_371),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_426),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_496),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_497),
.A2(n_383),
.B1(n_400),
.B2(n_342),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_426),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_496),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_434),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_471),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_480),
.B(n_371),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_492),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_427),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_494),
.B(n_418),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_427),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_474),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_427),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_496),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_497),
.A2(n_354),
.B1(n_361),
.B2(n_223),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_480),
.B(n_381),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_434),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_494),
.B(n_381),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_434),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_461),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_494),
.B(n_387),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_429),
.B(n_173),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_434),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_431),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_490),
.B(n_387),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_434),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_431),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_429),
.B(n_392),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_497),
.B(n_339),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_476),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_449),
.B(n_392),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_474),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_490),
.B(n_395),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_431),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_481),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_484),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_431),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_489),
.B(n_327),
.C(n_320),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_497),
.B(n_340),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_489),
.Y(n_618)
);

AO21x2_ASAP7_75t_L g619 ( 
.A1(n_498),
.A2(n_376),
.B(n_375),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_449),
.B(n_395),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_442),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_442),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_461),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_443),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_497),
.A2(n_174),
.B1(n_322),
.B2(n_305),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_443),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_490),
.A2(n_322),
.B1(n_179),
.B2(n_305),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_423),
.B(n_349),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_444),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_444),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_478),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_447),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_499),
.A2(n_389),
.B1(n_377),
.B2(n_385),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_431),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_447),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_484),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_448),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_478),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_449),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_499),
.B(n_382),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_499),
.A2(n_394),
.B1(n_391),
.B2(n_386),
.Y(n_642)
);

AO22x2_ASAP7_75t_L g643 ( 
.A1(n_499),
.A2(n_414),
.B1(n_212),
.B2(n_363),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_478),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_463),
.B(n_420),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_422),
.B(n_421),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_463),
.B(n_185),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_484),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_484),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_423),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_595),
.B(n_623),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_508),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_596),
.B(n_422),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_532),
.B(n_495),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_463),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_579),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_520),
.A2(n_452),
.B1(n_495),
.B2(n_463),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_508),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_512),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_604),
.A2(n_313),
.B1(n_323),
.B2(n_325),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_640),
.B(n_532),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_532),
.B(n_580),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_580),
.B(n_463),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_535),
.B(n_452),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_507),
.A2(n_485),
.B(n_487),
.C(n_450),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_580),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_554),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_646),
.B(n_455),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_580),
.B(n_462),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_629),
.B(n_462),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_625),
.A2(n_485),
.B1(n_487),
.B2(n_450),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_534),
.B(n_466),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_595),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_534),
.A2(n_469),
.B1(n_472),
.B2(n_453),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_534),
.B(n_466),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_526),
.B(n_558),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_560),
.B(n_446),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_526),
.B(n_466),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_558),
.B(n_466),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_554),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_625),
.B(n_475),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_566),
.B(n_475),
.Y(n_684)
);

OR2x2_ASAP7_75t_SL g685 ( 
.A(n_514),
.B(n_445),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_560),
.B(n_451),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_572),
.B(n_469),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_572),
.B(n_472),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_516),
.Y(n_689)
);

AND2x6_ASAP7_75t_SL g690 ( 
.A(n_604),
.B(n_445),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_575),
.B(n_455),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_522),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_539),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_522),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_516),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_575),
.B(n_448),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_603),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_607),
.B(n_453),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_437),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_589),
.B(n_454),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_604),
.A2(n_179),
.B1(n_188),
.B2(n_194),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_573),
.B(n_468),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_539),
.A2(n_430),
.B1(n_483),
.B2(n_313),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_589),
.B(n_581),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_511),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_620),
.B(n_454),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_593),
.B(n_456),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_569),
.B(n_437),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_527),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_600),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_584),
.B(n_456),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_628),
.B(n_493),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_590),
.B(n_186),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_628),
.B(n_493),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_537),
.B(n_457),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_527),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_581),
.B(n_457),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_552),
.B(n_459),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_616),
.B(n_459),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_479),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_583),
.B(n_479),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_586),
.B(n_479),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_528),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_586),
.B(n_486),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_486),
.Y(n_725)
);

BUFx6f_ASAP7_75t_SL g726 ( 
.A(n_604),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_604),
.A2(n_191),
.B1(n_193),
.B2(n_304),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_617),
.A2(n_188),
.B1(n_194),
.B2(n_323),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_501),
.B(n_486),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_617),
.A2(n_191),
.B1(n_193),
.B2(n_304),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_609),
.B(n_553),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_L g732 ( 
.A(n_507),
.B(n_326),
.C(n_325),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_528),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_517),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_608),
.B(n_488),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_608),
.B(n_488),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_517),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_578),
.B(n_198),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_612),
.B(n_488),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_647),
.B(n_326),
.C(n_334),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_591),
.B(n_360),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_645),
.B(n_641),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_643),
.A2(n_498),
.B1(n_437),
.B2(n_363),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_515),
.B(n_310),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_613),
.B(n_310),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_519),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_613),
.B(n_315),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_618),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_618),
.B(n_315),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_621),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_641),
.B(n_329),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_515),
.B(n_329),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_621),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_641),
.B(n_330),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_509),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_641),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_622),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_503),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_515),
.B(n_330),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_641),
.B(n_230),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_509),
.B(n_360),
.Y(n_761)
);

INVx8_ASAP7_75t_L g762 ( 
.A(n_617),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_617),
.B(n_231),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_503),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_332),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_515),
.B(n_332),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_617),
.A2(n_206),
.B1(n_208),
.B2(n_299),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_504),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_511),
.B(n_234),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_624),
.Y(n_770)
);

BUFx6f_ASAP7_75t_SL g771 ( 
.A(n_597),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_624),
.B(n_236),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_627),
.B(n_240),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_515),
.B(n_172),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_511),
.A2(n_597),
.B1(n_631),
.B2(n_627),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_634),
.B(n_335),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_505),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_511),
.B(n_246),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_525),
.B(n_172),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_630),
.B(n_248),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_505),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_253),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_633),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_633),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_636),
.B(n_254),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_636),
.B(n_258),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_638),
.B(n_259),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_638),
.B(n_266),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_642),
.B(n_267),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_597),
.B(n_269),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_597),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_549),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_597),
.B(n_274),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_551),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_524),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_550),
.B(n_278),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_648),
.B(n_279),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_524),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_597),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_555),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_524),
.B(n_606),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_606),
.A2(n_290),
.B1(n_280),
.B2(n_282),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_597),
.B(n_288),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_643),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_556),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_555),
.A2(n_295),
.B1(n_296),
.B2(n_220),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_550),
.B(n_1),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_525),
.B(n_172),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_756),
.B(n_648),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_652),
.Y(n_810)
);

INVx5_ASAP7_75t_L g811 ( 
.A(n_762),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_762),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_SL g813 ( 
.A1(n_685),
.A2(n_506),
.B1(n_643),
.B2(n_256),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_659),
.B(n_606),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_658),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_670),
.B(n_562),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_656),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_689),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_743),
.B(n_643),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_659),
.B(n_648),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_695),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_673),
.A2(n_649),
.B1(n_614),
.B2(n_637),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_756),
.B(n_649),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_675),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_659),
.B(n_614),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_659),
.B(n_614),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_668),
.B(n_637),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_660),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_734),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_665),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_762),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_670),
.B(n_562),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_737),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_672),
.B(n_563),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_755),
.B(n_649),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_668),
.B(n_637),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_653),
.B(n_563),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_650),
.B(n_564),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_650),
.B(n_564),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_698),
.B(n_568),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_673),
.B(n_525),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_651),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_684),
.A2(n_807),
.B(n_683),
.C(n_752),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_686),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_705),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_726),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_697),
.B(n_550),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_710),
.B(n_561),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_761),
.B(n_561),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_698),
.B(n_568),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_727),
.B(n_730),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_714),
.A2(n_644),
.B1(n_639),
.B2(n_605),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_662),
.B(n_525),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_758),
.Y(n_856)
);

NOR2x2_ASAP7_75t_L g857 ( 
.A(n_702),
.B(n_576),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_706),
.B(n_605),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_795),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_743),
.A2(n_644),
.B1(n_639),
.B2(n_611),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_682),
.Y(n_861)
);

INVx5_ASAP7_75t_L g862 ( 
.A(n_729),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_692),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_694),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_763),
.B(n_525),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_709),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_SL g867 ( 
.A(n_732),
.B(n_506),
.C(n_200),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_716),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_706),
.B(n_611),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_723),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_733),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_763),
.B(n_543),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_726),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_764),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_748),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_750),
.B(n_626),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_669),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_753),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_742),
.A2(n_547),
.B1(n_542),
.B2(n_531),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_705),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_795),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_757),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_798),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_663),
.B(n_543),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_768),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_770),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_783),
.B(n_626),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_784),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_666),
.B(n_632),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_664),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_666),
.B(n_632),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_703),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_729),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_690),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_671),
.B(n_543),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_760),
.A2(n_506),
.B1(n_235),
.B2(n_238),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_742),
.B(n_635),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_777),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_781),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_667),
.B(n_557),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_729),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_SL g903 ( 
.A(n_654),
.B(n_561),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_767),
.B(n_543),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_792),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_797),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_674),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_729),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_794),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_729),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_800),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_676),
.B(n_559),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_676),
.B(n_559),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_760),
.A2(n_654),
.B1(n_731),
.B2(n_738),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_805),
.B(n_570),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_711),
.B(n_570),
.Y(n_916)
);

BUFx8_ASAP7_75t_SL g917 ( 
.A(n_797),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_717),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_712),
.B(n_635),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_657),
.B(n_543),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_776),
.A2(n_577),
.B1(n_619),
.B2(n_541),
.Y(n_921)
);

BUFx8_ASAP7_75t_L g922 ( 
.A(n_771),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_720),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_798),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_684),
.A2(n_500),
.B(n_502),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_799),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_711),
.B(n_577),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_661),
.B(n_582),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_721),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_707),
.B(n_582),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_655),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_707),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_701),
.B(n_582),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_775),
.B(n_547),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_791),
.B(n_521),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_722),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_751),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_715),
.B(n_585),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_724),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_715),
.A2(n_533),
.B(n_538),
.C(n_540),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_SL g941 ( 
.A1(n_728),
.A2(n_221),
.B1(n_197),
.B2(n_201),
.Y(n_941)
);

NAND2x1_ASAP7_75t_L g942 ( 
.A(n_735),
.B(n_547),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_718),
.B(n_585),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_718),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_691),
.B(n_585),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_736),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_738),
.A2(n_530),
.B1(n_531),
.B2(n_533),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_754),
.B(n_588),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_739),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_687),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_688),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_683),
.A2(n_804),
.B1(n_713),
.B2(n_677),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_771),
.Y(n_953)
);

AO22x1_ASAP7_75t_L g954 ( 
.A1(n_740),
.A2(n_565),
.B1(n_437),
.B2(n_226),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_696),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_700),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_791),
.B(n_588),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_780),
.B(n_588),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_780),
.B(n_599),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_787),
.B(n_599),
.Y(n_960)
);

BUFx8_ASAP7_75t_L g961 ( 
.A(n_806),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_787),
.B(n_599),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_788),
.B(n_602),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_719),
.B(n_565),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_788),
.A2(n_619),
.B1(n_541),
.B2(n_529),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_680),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_678),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_704),
.B(n_789),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_681),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_725),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_772),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_807),
.A2(n_542),
.B(n_530),
.C(n_538),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_801),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_774),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_774),
.Y(n_975)
);

NOR2x2_ASAP7_75t_L g976 ( 
.A(n_806),
.B(n_592),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_769),
.A2(n_546),
.B1(n_540),
.B2(n_513),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_773),
.B(n_602),
.Y(n_978)
);

BUFx12f_ASAP7_75t_SL g979 ( 
.A(n_778),
.Y(n_979)
);

INVx5_ASAP7_75t_L g980 ( 
.A(n_699),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_782),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_778),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_745),
.B(n_610),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_785),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_786),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_779),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_747),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_790),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_749),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_842),
.A2(n_708),
.B(n_741),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_944),
.B(n_765),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_812),
.B(n_793),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_842),
.A2(n_752),
.B(n_744),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_844),
.B(n_802),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_932),
.B(n_796),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_R g996 ( 
.A(n_817),
.B(n_803),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_SL g997 ( 
.A(n_961),
.B(n_565),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_820),
.B(n_501),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_811),
.B(n_812),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_852),
.A2(n_869),
.B(n_858),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_852),
.A2(n_766),
.B(n_759),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_811),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_818),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_861),
.Y(n_1004)
);

HAxp5_ASAP7_75t_L g1005 ( 
.A(n_819),
.B(n_846),
.CON(n_1005),
.SN(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_858),
.A2(n_759),
.B(n_808),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_810),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_853),
.A2(n_971),
.B(n_989),
.C(n_987),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_825),
.B(n_610),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_811),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_869),
.A2(n_808),
.B(n_500),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_981),
.A2(n_635),
.B(n_610),
.C(n_615),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_873),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_811),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_L g1015 ( 
.A(n_897),
.B(n_867),
.C(n_941),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_816),
.A2(n_502),
.B(n_546),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_822),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_898),
.A2(n_594),
.B(n_598),
.C(n_601),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_926),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_819),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_984),
.A2(n_615),
.B(n_594),
.C(n_601),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_918),
.A2(n_615),
.B1(n_598),
.B2(n_529),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_815),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_820),
.A2(n_548),
.B1(n_523),
.B2(n_536),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_829),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_813),
.A2(n_548),
.B1(n_523),
.B2(n_536),
.Y(n_1026)
);

AOI22x1_ASAP7_75t_L g1027 ( 
.A1(n_958),
.A2(n_521),
.B1(n_545),
.B2(n_513),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_877),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_816),
.A2(n_513),
.B(n_544),
.Y(n_1029)
);

XNOR2xp5_ASAP7_75t_L g1030 ( 
.A(n_892),
.B(n_619),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_832),
.B(n_518),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_919),
.B(n_518),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_867),
.B(n_518),
.C(n_544),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_919),
.A2(n_961),
.B1(n_898),
.B2(n_906),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_893),
.A2(n_544),
.B1(n_545),
.B2(n_437),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_979),
.B(n_922),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_830),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_833),
.A2(n_587),
.B1(n_574),
.B2(n_571),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_835),
.A2(n_587),
.B1(n_574),
.B2(n_571),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_985),
.A2(n_424),
.B(n_425),
.C(n_571),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_834),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_936),
.B(n_571),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_937),
.B(n_571),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_851),
.B(n_5),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_962),
.A2(n_424),
.B(n_425),
.C(n_8),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_851),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_895),
.B(n_5),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_841),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_832),
.B(n_565),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_809),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_831),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_939),
.B(n_574),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_946),
.B(n_574),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_959),
.A2(n_7),
.B(n_9),
.C(n_12),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_873),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_SL g1056 ( 
.A1(n_896),
.A2(n_437),
.B(n_172),
.C(n_215),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_848),
.B(n_565),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_924),
.B(n_587),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_587),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_835),
.A2(n_587),
.B(n_250),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_838),
.A2(n_297),
.B1(n_207),
.B2(n_210),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_849),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_924),
.B(n_247),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_809),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_924),
.B(n_241),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_922),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_959),
.A2(n_960),
.B(n_963),
.C(n_956),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_849),
.A2(n_251),
.B1(n_219),
.B2(n_202),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_856),
.Y(n_1069)
);

CKINVDCx8_ASAP7_75t_R g1070 ( 
.A(n_836),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_923),
.B(n_437),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_894),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_929),
.B(n_437),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_SL g1074 ( 
.A(n_953),
.B(n_565),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_838),
.A2(n_273),
.B(n_298),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_960),
.A2(n_237),
.B(n_293),
.C(n_292),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_894),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_963),
.A2(n_228),
.B(n_287),
.C(n_281),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_901),
.A2(n_925),
.B(n_896),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_889),
.B(n_172),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_955),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_845),
.A2(n_211),
.B(n_222),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_931),
.B(n_850),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_894),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_824),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_917),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_901),
.A2(n_261),
.B(n_233),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_889),
.B(n_172),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_953),
.B(n_426),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_940),
.A2(n_23),
.B(n_26),
.C(n_27),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_847),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_928),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_R g1093 ( 
.A(n_903),
.B(n_106),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_857),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_925),
.A2(n_426),
.B(n_110),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_924),
.B(n_426),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_957),
.B(n_426),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_891),
.B(n_215),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_863),
.A2(n_868),
.B1(n_882),
.B2(n_870),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_902),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_864),
.B(n_34),
.C(n_37),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_916),
.A2(n_927),
.B(n_891),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_SL g1103 ( 
.A(n_866),
.B(n_37),
.C(n_40),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_874),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_871),
.Y(n_1105)
);

BUFx2_ASAP7_75t_SL g1106 ( 
.A(n_862),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_875),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_878),
.B(n_45),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_SL g1109 ( 
.A1(n_978),
.A2(n_48),
.B(n_215),
.C(n_172),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_902),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_886),
.B(n_172),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_902),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_908),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_SL g1114 ( 
.A(n_862),
.B(n_58),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_L g1115 ( 
.A1(n_845),
.A2(n_215),
.B(n_67),
.C(n_69),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_839),
.B(n_215),
.Y(n_1116)
);

AOI22x1_ASAP7_75t_L g1117 ( 
.A1(n_973),
.A2(n_215),
.B1(n_77),
.B2(n_84),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_950),
.B(n_66),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_938),
.A2(n_215),
.B(n_88),
.C(n_90),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_839),
.B(n_215),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_824),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_888),
.B(n_169),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_916),
.A2(n_86),
.B(n_96),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_909),
.B(n_117),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_933),
.A2(n_120),
.B(n_121),
.C(n_122),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_957),
.B(n_123),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_951),
.B(n_125),
.Y(n_1127)
);

INVx3_ASAP7_75t_SL g1128 ( 
.A(n_976),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_983),
.A2(n_128),
.B(n_129),
.C(n_132),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_840),
.B(n_150),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_938),
.A2(n_153),
.B(n_163),
.C(n_843),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_935),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_935),
.B(n_862),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_890),
.B(n_862),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_965),
.A2(n_972),
.B(n_930),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_908),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1128),
.B(n_890),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1083),
.B(n_967),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_1091),
.B(n_908),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1135),
.A2(n_965),
.B(n_840),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1121),
.B(n_910),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1000),
.A2(n_943),
.B(n_927),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1102),
.A2(n_945),
.B(n_915),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1007),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1015),
.B(n_1008),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1038),
.A2(n_945),
.B(n_915),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1044),
.B(n_907),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_998),
.B(n_907),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1038),
.A2(n_865),
.B(n_872),
.Y(n_1149)
);

NAND3x1_ASAP7_75t_L g1150 ( 
.A(n_1034),
.B(n_970),
.C(n_947),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1090),
.B(n_968),
.C(n_879),
.Y(n_1151)
);

AOI221x1_ASAP7_75t_L g1152 ( 
.A1(n_1082),
.A2(n_988),
.B1(n_912),
.B2(n_913),
.C(n_966),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1023),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1030),
.A2(n_968),
.B1(n_920),
.B2(n_912),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_SL g1155 ( 
.A(n_1081),
.B(n_952),
.C(n_921),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1050),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1118),
.A2(n_1127),
.B(n_1067),
.C(n_1082),
.Y(n_1157)
);

NOR4xp25_ASAP7_75t_L g1158 ( 
.A(n_1107),
.B(n_952),
.C(n_921),
.D(n_948),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1014),
.B(n_967),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_1094),
.B(n_968),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1064),
.B(n_854),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1079),
.A2(n_942),
.B(n_934),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1025),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1135),
.A2(n_823),
.B(n_977),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1039),
.A2(n_980),
.B(n_876),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1039),
.A2(n_855),
.B(n_884),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1095),
.A2(n_934),
.B(n_876),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_997),
.B(n_910),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1085),
.B(n_854),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1051),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_1107),
.A2(n_988),
.B1(n_913),
.B2(n_967),
.C(n_975),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1105),
.B(n_969),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1016),
.A2(n_887),
.B(n_860),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1014),
.B(n_910),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_1036),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1131),
.A2(n_904),
.B(n_973),
.C(n_974),
.Y(n_1176)
);

AND2x6_ASAP7_75t_L g1177 ( 
.A(n_1133),
.B(n_986),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1009),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1046),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_995),
.B(n_860),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1027),
.A2(n_821),
.B(n_814),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1011),
.A2(n_821),
.B(n_826),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_993),
.A2(n_1001),
.B(n_1006),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1092),
.A2(n_986),
.B(n_974),
.C(n_883),
.Y(n_1184)
);

AO21x1_ASAP7_75t_L g1185 ( 
.A1(n_1130),
.A2(n_827),
.B(n_828),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1066),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_990),
.A2(n_900),
.A3(n_911),
.B(n_905),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1130),
.A2(n_980),
.B(n_837),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_SL g1189 ( 
.A(n_1086),
.B(n_859),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1029),
.A2(n_1056),
.B(n_1115),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1042),
.A2(n_881),
.B(n_954),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1014),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1004),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1133),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_994),
.B(n_885),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1099),
.B(n_899),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1099),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1126),
.A2(n_964),
.B(n_880),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_999),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1052),
.A2(n_964),
.B(n_1053),
.Y(n_1200)
);

AND2x6_ASAP7_75t_L g1201 ( 
.A(n_999),
.B(n_1084),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_991),
.B(n_1070),
.Y(n_1202)
);

AOI221x1_ASAP7_75t_L g1203 ( 
.A1(n_1119),
.A2(n_1033),
.B1(n_1123),
.B2(n_1022),
.C(n_1087),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1003),
.B(n_1017),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1045),
.A2(n_1054),
.B(n_1021),
.C(n_1125),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1037),
.B(n_1041),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1048),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1022),
.A2(n_1065),
.B(n_1063),
.C(n_1058),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1080),
.A2(n_1098),
.B(n_1088),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1018),
.A2(n_1040),
.B(n_1053),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1122),
.A2(n_1124),
.B(n_1059),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1069),
.Y(n_1212)
);

AOI221x1_ASAP7_75t_L g1213 ( 
.A1(n_1061),
.A2(n_1060),
.B1(n_1098),
.B2(n_1080),
.C(n_1088),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1116),
.A2(n_1120),
.B(n_1117),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1104),
.Y(n_1215)
);

O2A1O1Ixp5_ASAP7_75t_L g1216 ( 
.A1(n_1096),
.A2(n_1097),
.B(n_1061),
.C(n_1109),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1028),
.B(n_1020),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1116),
.A2(n_1120),
.B(n_1059),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1134),
.A2(n_1129),
.B(n_1089),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1108),
.B(n_1132),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1071),
.A2(n_1073),
.A3(n_1076),
.B(n_1078),
.Y(n_1221)
);

AO21x1_ASAP7_75t_L g1222 ( 
.A1(n_1043),
.A2(n_1012),
.B(n_1075),
.Y(n_1222)
);

NAND3xp33_ASAP7_75t_L g1223 ( 
.A(n_1101),
.B(n_1103),
.C(n_1062),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1032),
.A2(n_1073),
.B(n_1071),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1089),
.A2(n_1110),
.B(n_1113),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1110),
.A2(n_1113),
.B(n_1002),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1002),
.A2(n_1111),
.B(n_1024),
.Y(n_1227)
);

AOI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1114),
.A2(n_992),
.B(n_1031),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_992),
.A2(n_1031),
.B(n_1049),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_996),
.B(n_1068),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1047),
.B(n_1005),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1026),
.A2(n_1035),
.B(n_1106),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1057),
.B(n_1136),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_992),
.A2(n_1074),
.B(n_1112),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1057),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_SL g1236 ( 
.A(n_1013),
.B(n_1055),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1084),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1074),
.A2(n_1136),
.B(n_1112),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1093),
.A2(n_1077),
.B(n_1072),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1072),
.A2(n_1077),
.B(n_1010),
.Y(n_1240)
);

NAND3x1_ASAP7_75t_L g1241 ( 
.A(n_1019),
.B(n_997),
.C(n_1010),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1019),
.B(n_1100),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1100),
.A2(n_845),
.B(n_1135),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1019),
.A2(n_1000),
.B(n_1102),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1000),
.A2(n_1102),
.B(n_1038),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1000),
.A2(n_1102),
.B(n_1038),
.Y(n_1246)
);

AO21x1_ASAP7_75t_L g1247 ( 
.A1(n_1067),
.A2(n_1082),
.B(n_1015),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1067),
.A2(n_833),
.B(n_816),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1083),
.B(n_982),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1094),
.B(n_844),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1008),
.A2(n_914),
.B(n_932),
.C(n_672),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1008),
.A2(n_914),
.B(n_932),
.C(n_672),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1135),
.A2(n_1079),
.B(n_845),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_SL g1254 ( 
.A1(n_1067),
.A2(n_1102),
.B(n_1135),
.Y(n_1254)
);

AOI31xp67_ASAP7_75t_L g1255 ( 
.A1(n_1080),
.A2(n_896),
.A3(n_1098),
.B(n_1088),
.Y(n_1255)
);

BUFx8_ASAP7_75t_L g1256 ( 
.A(n_1086),
.Y(n_1256)
);

OAI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1015),
.A2(n_672),
.B(n_383),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1102),
.B(n_918),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1135),
.A2(n_845),
.B(n_1082),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1008),
.A2(n_914),
.B(n_932),
.C(n_672),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1007),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1083),
.B(n_982),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1079),
.A2(n_1095),
.B(n_925),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1128),
.B(n_560),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1004),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1014),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1009),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_991),
.A2(n_853),
.B(n_672),
.C(n_573),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1000),
.A2(n_1102),
.B(n_1038),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1083),
.B(n_932),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1094),
.A2(n_539),
.B1(n_432),
.B2(n_813),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1083),
.B(n_932),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1007),
.Y(n_1273)
);

AOI221x1_ASAP7_75t_L g1274 ( 
.A1(n_1015),
.A2(n_813),
.B1(n_1082),
.B2(n_897),
.C(n_867),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1000),
.A2(n_1102),
.B(n_1038),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1036),
.Y(n_1276)
);

O2A1O1Ixp5_ASAP7_75t_L g1277 ( 
.A1(n_1082),
.A2(n_853),
.B(n_1135),
.C(n_995),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1083),
.B(n_932),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1008),
.A2(n_914),
.B(n_932),
.C(n_672),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1083),
.B(n_932),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1000),
.A2(n_1102),
.B(n_1038),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1007),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1079),
.A2(n_1095),
.B(n_925),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1000),
.A2(n_1102),
.B(n_1038),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1246),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1257),
.A2(n_1186),
.B(n_1230),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1284),
.A2(n_1269),
.B(n_1245),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1275),
.A2(n_1281),
.B(n_1183),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1183),
.A2(n_1214),
.B(n_1190),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1192),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1140),
.A2(n_1259),
.B(n_1157),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1175),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1228),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1153),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1209),
.A2(n_1218),
.B(n_1167),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1277),
.A2(n_1252),
.B(n_1251),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1259),
.A2(n_1213),
.B(n_1152),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1278),
.B(n_1280),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1211),
.B(n_1234),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1244),
.A2(n_1162),
.B(n_1143),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1140),
.A2(n_1171),
.B(n_1243),
.Y(n_1302)
);

INVxp67_ASAP7_75t_SL g1303 ( 
.A(n_1196),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1173),
.A2(n_1142),
.B(n_1165),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1271),
.A2(n_1155),
.B1(n_1247),
.B2(n_1145),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1193),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1164),
.A2(n_1154),
.B1(n_1151),
.B2(n_1264),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1163),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1248),
.A2(n_1146),
.B(n_1258),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1265),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1249),
.B(n_1262),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1187),
.Y(n_1312)
);

NAND2x1_ASAP7_75t_L g1313 ( 
.A(n_1254),
.B(n_1198),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1201),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1170),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1182),
.A2(n_1200),
.B(n_1243),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1260),
.A2(n_1279),
.B(n_1268),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1258),
.A2(n_1164),
.B(n_1158),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1274),
.A2(n_1208),
.B(n_1216),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1139),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1188),
.A2(n_1149),
.B(n_1166),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1178),
.B(n_1179),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1256),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1256),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1210),
.A2(n_1224),
.B(n_1181),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1223),
.A2(n_1151),
.B1(n_1197),
.B2(n_1267),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1210),
.A2(n_1219),
.B(n_1191),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1194),
.B(n_1199),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1266),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1253),
.A2(n_1185),
.B(n_1227),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1199),
.B(n_1266),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1168),
.A2(n_1203),
.B(n_1253),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1148),
.B(n_1220),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1223),
.A2(n_1180),
.B1(n_1205),
.B2(n_1150),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1261),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1179),
.B(n_1172),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1239),
.B(n_1159),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1242),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1276),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1201),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1226),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1250),
.B(n_1138),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1158),
.A2(n_1176),
.B(n_1184),
.Y(n_1343)
);

BUFx8_ASAP7_75t_L g1344 ( 
.A(n_1137),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1161),
.A2(n_1169),
.B1(n_1195),
.B2(n_1231),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1148),
.A2(n_1222),
.B(n_1232),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1225),
.A2(n_1229),
.B(n_1238),
.Y(n_1347)
);

NAND2x1p5_ASAP7_75t_L g1348 ( 
.A(n_1189),
.B(n_1235),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1240),
.A2(n_1241),
.B(n_1174),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1202),
.B(n_1233),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1174),
.A2(n_1282),
.B(n_1273),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1160),
.B(n_1217),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1201),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1237),
.A2(n_1255),
.B(n_1206),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1141),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1177),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1204),
.A2(n_1206),
.B(n_1215),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1207),
.A2(n_1212),
.B1(n_1204),
.B2(n_1177),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1177),
.B(n_1141),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1236),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1177),
.B(n_1221),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_SL g1362 ( 
.A1(n_1221),
.A2(n_1157),
.B(n_1279),
.C(n_1252),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1193),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1175),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1193),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1144),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1144),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1271),
.A2(n_813),
.B1(n_820),
.B2(n_432),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1194),
.B(n_1014),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1271),
.A2(n_813),
.B1(n_820),
.B2(n_432),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1183),
.A2(n_1246),
.B(n_1245),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1187),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1144),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1175),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1147),
.B(n_1178),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1274),
.A2(n_702),
.B1(n_590),
.B2(n_914),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1156),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1187),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1192),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1213),
.A2(n_1157),
.A3(n_1152),
.B(n_1171),
.Y(n_1385)
);

BUFx8_ASAP7_75t_SL g1386 ( 
.A(n_1175),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1144),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1157),
.A2(n_1277),
.B(n_1252),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1144),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1156),
.Y(n_1391)
);

AO31x2_ASAP7_75t_L g1392 ( 
.A1(n_1213),
.A2(n_1157),
.A3(n_1152),
.B(n_1171),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1144),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1271),
.A2(n_813),
.B1(n_820),
.B2(n_432),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1193),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1147),
.B(n_1178),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1144),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1213),
.A2(n_1157),
.A3(n_1152),
.B(n_1171),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1183),
.A2(n_1246),
.B(n_1245),
.Y(n_1401)
);

NAND2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1189),
.B(n_1093),
.Y(n_1402)
);

AND2x6_ASAP7_75t_L g1403 ( 
.A(n_1197),
.B(n_1133),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1257),
.A2(n_702),
.B1(n_590),
.B2(n_1157),
.C(n_573),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1144),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1144),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1157),
.A2(n_1277),
.B(n_1252),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1263),
.A2(n_1283),
.B(n_1281),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1156),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1306),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1404),
.A2(n_1305),
.B1(n_1307),
.B2(n_1381),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_SL g1414 ( 
.A1(n_1292),
.A2(n_1366),
.B(n_1299),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1317),
.A2(n_1334),
.B(n_1314),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1344),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1354),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1309),
.A2(n_1362),
.B(n_1389),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1354),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1380),
.B(n_1398),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1362),
.A2(n_1408),
.B(n_1297),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1344),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1330),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1305),
.A2(n_1307),
.B1(n_1372),
.B2(n_1370),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1370),
.A2(n_1396),
.B1(n_1372),
.B2(n_1286),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1352),
.B(n_1350),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1287),
.A2(n_1363),
.B(n_1285),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1333),
.B(n_1336),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1322),
.B(n_1382),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1396),
.A2(n_1360),
.B1(n_1326),
.B2(n_1311),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1338),
.B(n_1391),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1411),
.B(n_1295),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1386),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1308),
.B(n_1315),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1330),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1314),
.A2(n_1340),
.B(n_1319),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_SL g1437 ( 
.A(n_1300),
.B(n_1340),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1335),
.B(n_1368),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1369),
.B(n_1376),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1344),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1388),
.B(n_1390),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1394),
.B(n_1399),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1406),
.B(n_1407),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1342),
.B(n_1303),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1287),
.A2(n_1410),
.B(n_1285),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1332),
.A2(n_1402),
.B(n_1313),
.C(n_1327),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1348),
.A2(n_1345),
.B1(n_1358),
.B2(n_1331),
.Y(n_1447)
);

AOI31xp33_ASAP7_75t_L g1448 ( 
.A1(n_1324),
.A2(n_1320),
.A3(n_1402),
.B(n_1328),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1327),
.A2(n_1358),
.B(n_1351),
.C(n_1288),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1363),
.A2(n_1410),
.B(n_1375),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1357),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1357),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1357),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1348),
.A2(n_1331),
.B1(n_1367),
.B2(n_1323),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1373),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1397),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1325),
.A2(n_1353),
.B(n_1356),
.C(n_1294),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1318),
.B(n_1291),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1324),
.A2(n_1323),
.B(n_1386),
.Y(n_1459)
);

BUFx4f_ASAP7_75t_L g1460 ( 
.A(n_1356),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1310),
.B(n_1364),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1290),
.B(n_1384),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1401),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1403),
.B(n_1300),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1403),
.B(n_1349),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1293),
.A2(n_1365),
.B1(n_1378),
.B2(n_1339),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1375),
.A2(n_1409),
.B(n_1405),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1346),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1301),
.A2(n_1298),
.B(n_1304),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1328),
.A2(n_1329),
.B1(n_1293),
.B2(n_1365),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1329),
.A2(n_1378),
.B1(n_1339),
.B2(n_1302),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1349),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1302),
.A2(n_1298),
.B1(n_1355),
.B2(n_1337),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_SL g1474 ( 
.A1(n_1302),
.A2(n_1361),
.B1(n_1359),
.B2(n_1337),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1355),
.B(n_1343),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1346),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1385),
.B(n_1392),
.Y(n_1477)
);

AOI21x1_ASAP7_75t_SL g1478 ( 
.A1(n_1289),
.A2(n_1400),
.B(n_1392),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1385),
.B(n_1392),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1294),
.A2(n_1341),
.B(n_1371),
.C(n_1383),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1377),
.A2(n_1409),
.B(n_1405),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1371),
.A2(n_1341),
.B1(n_1400),
.B2(n_1312),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1316),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1316),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1347),
.B(n_1321),
.Y(n_1485)
);

BUFx10_ASAP7_75t_L g1486 ( 
.A(n_1400),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1347),
.B(n_1289),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1304),
.A2(n_1379),
.B(n_1393),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1374),
.A2(n_1321),
.B1(n_1296),
.B2(n_1377),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_SL g1490 ( 
.A1(n_1296),
.A2(n_1379),
.B(n_1387),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1395),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1395),
.B(n_1380),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1317),
.B(n_1157),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1380),
.B(n_1398),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1432),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1434),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1492),
.B(n_1486),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1429),
.B(n_1444),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1490),
.A2(n_1469),
.B(n_1488),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1451),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1486),
.B(n_1494),
.Y(n_1501)
);

AOI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1493),
.A2(n_1424),
.B1(n_1425),
.B2(n_1430),
.C(n_1413),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1438),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1431),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1418),
.A2(n_1458),
.B(n_1449),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1477),
.B(n_1479),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1491),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1452),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1439),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1420),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1441),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1426),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1442),
.Y(n_1513)
);

BUFx2_ASAP7_75t_SL g1514 ( 
.A(n_1412),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1443),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1428),
.B(n_1493),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1485),
.A2(n_1449),
.B(n_1453),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1468),
.A2(n_1476),
.B(n_1489),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1468),
.A2(n_1476),
.B(n_1446),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1412),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1421),
.B(n_1456),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1473),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1475),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1455),
.B(n_1463),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1455),
.B(n_1463),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1482),
.B(n_1423),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1423),
.B(n_1435),
.Y(n_1527)
);

INVx5_ASAP7_75t_SL g1528 ( 
.A(n_1464),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1465),
.B(n_1472),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1471),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1435),
.B(n_1491),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1483),
.B(n_1484),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1478),
.A2(n_1472),
.B(n_1480),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1433),
.B(n_1466),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1483),
.B(n_1484),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1462),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1415),
.A2(n_1447),
.B1(n_1454),
.B2(n_1448),
.C(n_1461),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1416),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1417),
.B(n_1419),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1474),
.B(n_1436),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1417),
.B(n_1487),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1498),
.B(n_1457),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1496),
.B(n_1457),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1500),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1524),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1541),
.B(n_1524),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1525),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1541),
.B(n_1525),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1498),
.B(n_1445),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1497),
.B(n_1427),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1514),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1527),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1529),
.B(n_1437),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1497),
.B(n_1481),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1505),
.B(n_1481),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1540),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1505),
.B(n_1481),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1505),
.B(n_1450),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1539),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1533),
.B(n_1460),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1505),
.B(n_1517),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1506),
.B(n_1450),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1517),
.B(n_1467),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1562),
.A2(n_1565),
.B(n_1559),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1562),
.A2(n_1502),
.B(n_1534),
.C(n_1470),
.Y(n_1567)
);

AOI33xp33_ASAP7_75t_L g1568 ( 
.A1(n_1562),
.A2(n_1515),
.A3(n_1509),
.B1(n_1503),
.B2(n_1513),
.B3(n_1511),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1544),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1563),
.Y(n_1570)
);

AO21x2_ASAP7_75t_L g1571 ( 
.A1(n_1565),
.A2(n_1518),
.B(n_1517),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1547),
.B(n_1495),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1544),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1547),
.B(n_1563),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1543),
.A2(n_1565),
.B1(n_1522),
.B2(n_1530),
.C(n_1558),
.Y(n_1575)
);

OAI322xp33_ASAP7_75t_L g1576 ( 
.A1(n_1564),
.A2(n_1516),
.A3(n_1526),
.B1(n_1512),
.B2(n_1521),
.C1(n_1513),
.C2(n_1515),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1551),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1578)
);

OAI31xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1545),
.A2(n_1537),
.A3(n_1531),
.B(n_1535),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1552),
.B(n_1511),
.Y(n_1580)
);

OA332x1_ASAP7_75t_L g1581 ( 
.A1(n_1545),
.A2(n_1433),
.A3(n_1459),
.B1(n_1414),
.B2(n_1538),
.B3(n_1504),
.C1(n_1499),
.C2(n_1532),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1542),
.A2(n_1523),
.B1(n_1540),
.B2(n_1501),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1542),
.A2(n_1523),
.B1(n_1540),
.B2(n_1501),
.Y(n_1583)
);

AND2x6_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1528),
.Y(n_1584)
);

OAI31xp33_ASAP7_75t_L g1585 ( 
.A1(n_1542),
.A2(n_1526),
.A3(n_1507),
.B(n_1531),
.Y(n_1585)
);

NAND4xp25_ASAP7_75t_L g1586 ( 
.A(n_1556),
.B(n_1538),
.C(n_1532),
.D(n_1535),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1561),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.B(n_1536),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1556),
.A2(n_1518),
.B(n_1519),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1560),
.B(n_1510),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1554),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1546),
.B(n_1507),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1529),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1548),
.B(n_1520),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1551),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1569),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1566),
.B(n_1555),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1569),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1566),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1566),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1577),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1596),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1589),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1584),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1587),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1538),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1589),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1570),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1591),
.Y(n_1614)
);

AO21x2_ASAP7_75t_L g1615 ( 
.A1(n_1571),
.A2(n_1556),
.B(n_1558),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1559),
.C(n_1558),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1584),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1578),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1574),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1574),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1575),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1567),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1594),
.B(n_1555),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1580),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1571),
.Y(n_1627)
);

INVx6_ASAP7_75t_L g1628 ( 
.A(n_1616),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1624),
.A2(n_1583),
.B1(n_1582),
.B2(n_1557),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1621),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1615),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1579),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1614),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_L g1634 ( 
.A(n_1618),
.B(n_1586),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1613),
.B(n_1590),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1614),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1605),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1597),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1608),
.B(n_1616),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1616),
.B(n_1571),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1605),
.Y(n_1641)
);

OAI33xp33_ASAP7_75t_L g1642 ( 
.A1(n_1624),
.A2(n_1618),
.A3(n_1613),
.B1(n_1620),
.B2(n_1617),
.B3(n_1626),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1615),
.Y(n_1643)
);

AO21x2_ASAP7_75t_L g1644 ( 
.A1(n_1607),
.A2(n_1611),
.B(n_1627),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1623),
.B(n_1579),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1606),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1626),
.B(n_1590),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1597),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1617),
.B(n_1620),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1608),
.B(n_1594),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1592),
.Y(n_1651)
);

NAND4xp25_ASAP7_75t_L g1652 ( 
.A(n_1610),
.B(n_1586),
.C(n_1585),
.D(n_1581),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1599),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1585),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1622),
.B(n_1610),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1599),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1616),
.B(n_1592),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1619),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1619),
.B(n_1595),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1602),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1602),
.B(n_1571),
.Y(n_1664)
);

AOI322xp5_ASAP7_75t_L g1665 ( 
.A1(n_1598),
.A2(n_1559),
.A3(n_1555),
.B1(n_1550),
.B2(n_1576),
.C1(n_1593),
.C2(n_1587),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1615),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1602),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1631),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1628),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1635),
.B(n_1612),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1632),
.A2(n_1615),
.B(n_1602),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1639),
.B(n_1625),
.Y(n_1674)
);

INVxp33_ASAP7_75t_L g1675 ( 
.A(n_1639),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1641),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1634),
.B(n_1625),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1601),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1638),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1645),
.A2(n_1602),
.B(n_1604),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1637),
.B(n_1646),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1634),
.B(n_1598),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1648),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1658),
.B(n_1598),
.Y(n_1685)
);

NAND2x1_ASAP7_75t_SL g1686 ( 
.A(n_1630),
.B(n_1600),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1642),
.A2(n_1604),
.B1(n_1600),
.B2(n_1611),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1628),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1653),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1653),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1631),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1658),
.B(n_1609),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1631),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1628),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1651),
.B(n_1609),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1606),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1601),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1659),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1647),
.B(n_1603),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1643),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1657),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1643),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1686),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1673),
.A2(n_1683),
.B1(n_1652),
.B2(n_1697),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1672),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1672),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1686),
.Y(n_1709)
);

AOI22x1_ASAP7_75t_L g1710 ( 
.A1(n_1676),
.A2(n_1659),
.B1(n_1663),
.B2(n_1668),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1683),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1655),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1671),
.B(n_1649),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1700),
.B(n_1656),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1670),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1682),
.B(n_1688),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1673),
.A2(n_1600),
.B1(n_1604),
.B2(n_1654),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1675),
.B(n_1662),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1670),
.B(n_1650),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1674),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1674),
.B(n_1660),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1697),
.B(n_1688),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1679),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1679),
.Y(n_1724)
);

CKINVDCx16_ASAP7_75t_R g1725 ( 
.A(n_1694),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1694),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1677),
.B(n_1660),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1671),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1692),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

NAND2x1_ASAP7_75t_SL g1731 ( 
.A(n_1722),
.B(n_1719),
.Y(n_1731)
);

NOR4xp25_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1687),
.C(n_1677),
.D(n_1690),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1707),
.Y(n_1733)
);

OAI21xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1722),
.A2(n_1665),
.B(n_1685),
.Y(n_1734)
);

NAND2xp67_ASAP7_75t_SL g1735 ( 
.A(n_1727),
.B(n_1692),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1707),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1705),
.A2(n_1681),
.B1(n_1640),
.B2(n_1667),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1708),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1712),
.A2(n_1664),
.B1(n_1667),
.B2(n_1654),
.C(n_1640),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1710),
.A2(n_1665),
.B(n_1698),
.C(n_1663),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1728),
.B(n_1680),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1719),
.Y(n_1742)
);

OAI21xp33_ASAP7_75t_L g1743 ( 
.A1(n_1718),
.A2(n_1696),
.B(n_1678),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1725),
.B(n_1696),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1661),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1725),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1716),
.B(n_1685),
.C(n_1684),
.D(n_1703),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1729),
.B(n_1699),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1719),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1709),
.A2(n_1640),
.B1(n_1654),
.B2(n_1667),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1731),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1746),
.B(n_1726),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1746),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1742),
.B(n_1715),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1748),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1744),
.B(n_1715),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1733),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1734),
.B(n_1719),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1749),
.B(n_1720),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1738),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1743),
.B(n_1720),
.Y(n_1762)
);

AOI211xp5_ASAP7_75t_L g1763 ( 
.A1(n_1758),
.A2(n_1732),
.B(n_1740),
.C(n_1709),
.Y(n_1763)
);

OAI21xp33_ASAP7_75t_L g1764 ( 
.A1(n_1753),
.A2(n_1727),
.B(n_1714),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1751),
.A2(n_1745),
.B(n_1741),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1754),
.B(n_1721),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1751),
.A2(n_1737),
.B1(n_1711),
.B2(n_1710),
.Y(n_1767)
);

AOI221xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1752),
.A2(n_1747),
.B1(n_1741),
.B2(n_1711),
.C(n_1735),
.Y(n_1768)
);

NAND4xp75_ASAP7_75t_L g1769 ( 
.A(n_1756),
.B(n_1739),
.C(n_1721),
.D(n_1750),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1759),
.A2(n_1717),
.B1(n_1713),
.B2(n_1678),
.C(n_1724),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_SL g1771 ( 
.A(n_1755),
.B(n_1708),
.Y(n_1771)
);

OAI31xp33_ASAP7_75t_L g1772 ( 
.A1(n_1761),
.A2(n_1640),
.A3(n_1664),
.B(n_1713),
.Y(n_1772)
);

OAI21xp33_ASAP7_75t_L g1773 ( 
.A1(n_1762),
.A2(n_1689),
.B(n_1684),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1763),
.A2(n_1754),
.B1(n_1699),
.B2(n_1701),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1767),
.A2(n_1760),
.B(n_1757),
.Y(n_1775)
);

AOI222xp33_ASAP7_75t_L g1776 ( 
.A1(n_1770),
.A2(n_1730),
.B1(n_1724),
.B2(n_1723),
.C1(n_1664),
.C2(n_1607),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1766),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1769),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1765),
.A2(n_1695),
.B1(n_1669),
.B2(n_1704),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1774),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

NAND3xp33_ASAP7_75t_L g1782 ( 
.A(n_1778),
.B(n_1768),
.C(n_1764),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1775),
.B(n_1771),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1776),
.B(n_1651),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1779),
.Y(n_1785)
);

XNOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1778),
.B(n_1723),
.Y(n_1786)
);

AOI311xp33_ASAP7_75t_L g1787 ( 
.A1(n_1783),
.A2(n_1730),
.A3(n_1773),
.B(n_1772),
.C(n_1703),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1782),
.A2(n_1689),
.B1(n_1690),
.B2(n_1701),
.C(n_1695),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1786),
.B(n_1633),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1781),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1782),
.A2(n_1633),
.B(n_1636),
.Y(n_1791)
);

A2O1A1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1785),
.B(n_1784),
.C(n_1780),
.Y(n_1792)
);

AO22x1_ASAP7_75t_L g1793 ( 
.A1(n_1790),
.A2(n_1636),
.B1(n_1661),
.B2(n_1662),
.Y(n_1793)
);

NOR3xp33_ASAP7_75t_L g1794 ( 
.A(n_1789),
.B(n_1704),
.C(n_1702),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1793),
.B(n_1788),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1795),
.A2(n_1792),
.B1(n_1787),
.B2(n_1794),
.C(n_1704),
.Y(n_1796)
);

NAND4xp25_ASAP7_75t_L g1797 ( 
.A(n_1796),
.B(n_1664),
.C(n_1422),
.D(n_1440),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_1702),
.B1(n_1695),
.B2(n_1693),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1798),
.B(n_1702),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1797),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1799),
.Y(n_1801)
);

XOR2xp5_ASAP7_75t_L g1802 ( 
.A(n_1800),
.B(n_1629),
.Y(n_1802)
);

AOI222xp33_ASAP7_75t_SL g1803 ( 
.A1(n_1801),
.A2(n_1693),
.B1(n_1691),
.B2(n_1669),
.C1(n_1657),
.C2(n_1607),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1803),
.B(n_1802),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1804),
.B(n_1669),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1693),
.B1(n_1691),
.B2(n_1644),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1691),
.B1(n_1644),
.B2(n_1611),
.C(n_1607),
.Y(n_1807)
);

AOI211xp5_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1666),
.B(n_1611),
.C(n_1627),
.Y(n_1808)
);


endmodule