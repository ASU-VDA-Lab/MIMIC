module real_jpeg_25359_n_3 (n_0, n_21, n_1, n_2, n_20, n_3);

input n_0;
input n_21;
input n_1;
input n_2;
input n_20;

output n_3;

wire n_17;
wire n_8;
wire n_10;
wire n_9;
wire n_12;
wire n_6;
wire n_11;
wire n_14;
wire n_7;
wire n_18;
wire n_5;
wire n_4;
wire n_16;
wire n_15;
wire n_13;

INVx6_ASAP7_75t_SL g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g3 ( 
.A(n_4),
.B(n_11),
.Y(n_3)
);

NOR2xp33_ASAP7_75t_SL g4 ( 
.A(n_5),
.B(n_10),
.Y(n_4)
);

INVx1_ASAP7_75t_L g5 ( 
.A(n_6),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_9),
.Y(n_6)
);

INVx6_ASAP7_75t_SL g7 ( 
.A(n_8),
.Y(n_7)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_17),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_14),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_20),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_21),
.Y(n_16)
);


endmodule