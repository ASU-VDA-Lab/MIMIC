module fake_aes_11378_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NOR2x1p5_ASAP7_75t_L g3 ( .A(n_1), .B(n_2), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_1), .B(n_0), .Y(n_4) );
NAND2xp33_ASAP7_75t_SL g5 ( .A(n_0), .B(n_2), .Y(n_5) );
INVx2_ASAP7_75t_SL g6 ( .A(n_3), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_4), .B(n_5), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_6), .B(n_7), .Y(n_9) );
NOR3xp33_ASAP7_75t_L g10 ( .A(n_9), .B(n_7), .C(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
endmodule