module real_aes_16042_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_855, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_855;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g118 ( .A(n_0), .B(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_1), .A2(n_3), .B1(n_156), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_2), .A2(n_43), .B1(n_163), .B2(n_269), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_4), .A2(n_24), .B1(n_234), .B2(n_269), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_5), .A2(n_16), .B1(n_153), .B2(n_202), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_6), .A2(n_60), .B1(n_181), .B2(n_236), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_7), .A2(n_18), .B1(n_163), .B2(n_185), .Y(n_568) );
INVx1_ASAP7_75t_L g119 ( .A(n_8), .Y(n_119) );
INVx1_ASAP7_75t_L g496 ( .A(n_9), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_10), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_11), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_12), .A2(n_19), .B1(n_180), .B2(n_183), .Y(n_179) );
BUFx2_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
OR2x2_ASAP7_75t_L g135 ( .A(n_13), .B(n_39), .Y(n_135) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_15), .Y(n_207) );
INVx1_ASAP7_75t_L g497 ( .A(n_17), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_20), .A2(n_101), .B1(n_153), .B2(n_156), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_21), .A2(n_40), .B1(n_197), .B2(n_199), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_22), .B(n_154), .Y(n_247) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_23), .A2(n_56), .B(n_172), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_25), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_26), .Y(n_663) );
INVx4_ASAP7_75t_R g580 ( .A(n_27), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_28), .B(n_160), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_29), .A2(n_47), .B1(n_213), .B2(n_215), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_30), .A2(n_67), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_30), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_31), .A2(n_53), .B1(n_153), .B2(n_215), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_32), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_33), .B(n_197), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_34), .Y(n_260) );
INVx1_ASAP7_75t_L g593 ( .A(n_35), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_36), .B(n_269), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_SL g529 ( .A1(n_37), .A2(n_159), .B(n_163), .C(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_38), .A2(n_54), .B1(n_163), .B2(n_215), .Y(n_661) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_41), .A2(n_87), .B1(n_163), .B2(n_233), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_42), .A2(n_46), .B1(n_163), .B2(n_185), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_44), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_45), .A2(n_58), .B1(n_153), .B2(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g615 ( .A(n_48), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_49), .B(n_163), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_50), .Y(n_555) );
INVx2_ASAP7_75t_L g126 ( .A(n_51), .Y(n_126) );
INVx1_ASAP7_75t_L g113 ( .A(n_52), .Y(n_113) );
BUFx3_ASAP7_75t_L g839 ( .A(n_52), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_55), .A2(n_89), .B1(n_163), .B2(n_215), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_57), .Y(n_581) );
XNOR2xp5_ASAP7_75t_SL g507 ( .A(n_59), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_61), .A2(n_75), .B1(n_162), .B2(n_213), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_62), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_63), .A2(n_77), .B1(n_163), .B2(n_185), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_64), .A2(n_100), .B1(n_153), .B2(n_183), .Y(n_257) );
AND2x4_ASAP7_75t_L g149 ( .A(n_65), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g172 ( .A(n_66), .Y(n_172) );
INVx1_ASAP7_75t_L g509 ( .A(n_67), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_68), .A2(n_92), .B1(n_213), .B2(n_215), .Y(n_589) );
AO22x1_ASAP7_75t_L g546 ( .A1(n_69), .A2(n_76), .B1(n_199), .B2(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g150 ( .A(n_70), .Y(n_150) );
AND2x2_ASAP7_75t_L g533 ( .A(n_71), .B(n_253), .Y(n_533) );
INVx1_ASAP7_75t_L g490 ( .A(n_72), .Y(n_490) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_72), .B(n_494), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_73), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_74), .B(n_236), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_78), .B(n_269), .Y(n_556) );
INVx2_ASAP7_75t_L g160 ( .A(n_79), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_80), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_81), .B(n_253), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_82), .A2(n_99), .B1(n_215), .B2(n_236), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_83), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_84), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_85), .B(n_170), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_86), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_88), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_90), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_91), .B(n_253), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_93), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_94), .B(n_253), .Y(n_552) );
INVx1_ASAP7_75t_L g117 ( .A(n_95), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_95), .B(n_133), .Y(n_132) );
NAND2xp33_ASAP7_75t_L g250 ( .A(n_96), .B(n_154), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_97), .A2(n_187), .B(n_236), .C(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g582 ( .A(n_98), .B(n_583), .Y(n_582) );
NAND2xp33_ASAP7_75t_L g560 ( .A(n_102), .B(n_198), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_120), .B(n_848), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_111), .Y(n_105) );
OR2x6_ASAP7_75t_L g853 ( .A(n_106), .B(n_111), .Y(n_853) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2x1p5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_116), .Y(n_513) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g832 ( .A(n_117), .Y(n_832) );
OR2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_501), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_504), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g836 ( .A(n_126), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_126), .B(n_845), .Y(n_844) );
AOI31xp67_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_136), .A3(n_498), .B(n_501), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
CKINVDCx8_ASAP7_75t_R g503 ( .A(n_131), .Y(n_503) );
AND2x6_ASAP7_75t_SL g131 ( .A(n_132), .B(n_134), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_134), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2x1_ASAP7_75t_L g847 ( .A(n_135), .B(n_839), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_491), .Y(n_136) );
NAND2xp33_ASAP7_75t_SL g137 ( .A(n_138), .B(n_490), .Y(n_137) );
INVx2_ASAP7_75t_L g494 ( .A(n_138), .Y(n_494) );
OAI22x1_ASAP7_75t_L g511 ( .A1(n_138), .A2(n_512), .B1(n_514), .B2(n_831), .Y(n_511) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_399), .Y(n_138) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_139), .A2(n_399), .B(n_493), .Y(n_500) );
NOR2x1_ASAP7_75t_L g139 ( .A(n_140), .B(n_338), .Y(n_139) );
NAND4xp25_ASAP7_75t_L g140 ( .A(n_141), .B(n_289), .C(n_308), .D(n_319), .Y(n_140) );
O2A1O1Ixp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_220), .B(n_227), .C(n_261), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_192), .Y(n_142) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_143), .B(n_354), .C(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_L g435 ( .A(n_143), .B(n_317), .Y(n_435) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_176), .Y(n_143) );
AND2x2_ASAP7_75t_L g279 ( .A(n_144), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g297 ( .A(n_144), .B(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g314 ( .A(n_144), .Y(n_314) );
AND2x2_ASAP7_75t_L g359 ( .A(n_144), .B(n_194), .Y(n_359) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g224 ( .A(n_145), .Y(n_224) );
AND2x4_ASAP7_75t_L g307 ( .A(n_145), .B(n_298), .Y(n_307) );
AO31x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_151), .A3(n_167), .B(n_173), .Y(n_145) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_146), .A2(n_188), .A3(n_256), .B(n_259), .Y(n_255) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_147), .A2(n_575), .B(n_578), .Y(n_574) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AO31x2_ASAP7_75t_L g177 ( .A1(n_148), .A2(n_178), .A3(n_188), .B(n_190), .Y(n_177) );
AO31x2_ASAP7_75t_L g194 ( .A1(n_148), .A2(n_195), .A3(n_204), .B(n_206), .Y(n_194) );
AO31x2_ASAP7_75t_L g266 ( .A1(n_148), .A2(n_267), .A3(n_271), .B(n_272), .Y(n_266) );
AO31x2_ASAP7_75t_L g566 ( .A1(n_148), .A2(n_175), .A3(n_567), .B(n_570), .Y(n_566) );
BUFx10_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
INVx1_ASAP7_75t_L g532 ( .A(n_149), .Y(n_532) );
BUFx10_ASAP7_75t_L g564 ( .A(n_149), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_158), .B1(n_161), .B2(n_164), .Y(n_151) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_154), .Y(n_547) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g157 ( .A(n_155), .Y(n_157) );
INVx3_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
INVx1_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
INVx2_ASAP7_75t_L g234 ( .A(n_155), .Y(n_234) );
INVx1_ASAP7_75t_L g236 ( .A(n_155), .Y(n_236) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_155), .Y(n_269) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_157), .B(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_158), .A2(n_179), .B1(n_184), .B2(n_186), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_158), .A2(n_164), .B1(n_196), .B2(n_201), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_164), .B1(n_212), .B2(n_214), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_158), .A2(n_232), .B1(n_235), .B2(n_237), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_158), .A2(n_249), .B(n_250), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_158), .A2(n_186), .B1(n_257), .B2(n_258), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_158), .A2(n_164), .B1(n_268), .B2(n_270), .Y(n_267) );
OAI22x1_ASAP7_75t_L g567 ( .A1(n_158), .A2(n_237), .B1(n_568), .B2(n_569), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_158), .A2(n_237), .B1(n_589), .B2(n_590), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_158), .A2(n_542), .B1(n_660), .B2(n_661), .Y(n_659) );
INVx6_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g245 ( .A1(n_159), .A2(n_185), .B(n_246), .C(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_159), .B(n_546), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_159), .A2(n_560), .B(n_561), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_159), .A2(n_541), .B(n_546), .C(n_549), .Y(n_601) );
BUFx8_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
INVx1_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
INVx1_ASAP7_75t_L g528 ( .A(n_160), .Y(n_528) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g183 ( .A(n_163), .Y(n_183) );
INVx4_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g542 ( .A(n_165), .Y(n_542) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g558 ( .A(n_166), .Y(n_558) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_167), .A2(n_211), .A3(n_216), .B(n_218), .Y(n_210) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_167), .A2(n_574), .B(n_582), .Y(n_573) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g190 ( .A(n_169), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_169), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g175 ( .A(n_170), .Y(n_175) );
INVx2_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_170), .A2(n_532), .B(n_544), .Y(n_549) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_175), .B(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g225 ( .A(n_176), .B(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g282 ( .A(n_176), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_176), .Y(n_305) );
INVx1_ASAP7_75t_L g316 ( .A(n_176), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_176), .B(n_208), .Y(n_325) );
INVx2_ASAP7_75t_L g332 ( .A(n_176), .Y(n_332) );
INVx4_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g277 ( .A(n_177), .B(n_194), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_177), .B(n_284), .Y(n_350) );
AND2x2_ASAP7_75t_L g358 ( .A(n_177), .B(n_210), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_177), .B(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g411 ( .A(n_177), .Y(n_411) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_182), .B(n_577), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_185), .A2(n_555), .B(n_556), .C(n_557), .Y(n_554) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
AOI21x1_ASAP7_75t_L g520 ( .A1(n_188), .A2(n_521), .B(n_533), .Y(n_520) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_188), .A2(n_216), .A3(n_588), .B(n_592), .Y(n_587) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_189), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g583 ( .A(n_189), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_189), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_189), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g427 ( .A(n_193), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_208), .Y(n_193) );
INVx1_ASAP7_75t_L g226 ( .A(n_194), .Y(n_226) );
INVx1_ASAP7_75t_L g284 ( .A(n_194), .Y(n_284) );
INVx2_ASAP7_75t_L g318 ( .A(n_194), .Y(n_318) );
OR2x2_ASAP7_75t_L g322 ( .A(n_194), .B(n_210), .Y(n_322) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_194), .Y(n_371) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g213 ( .A(n_198), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_198), .A2(n_203), .B1(n_580), .B2(n_581), .Y(n_579) );
OAI21xp33_ASAP7_75t_SL g611 ( .A1(n_199), .A2(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AO31x2_ASAP7_75t_L g230 ( .A1(n_204), .A2(n_216), .A3(n_231), .B(n_238), .Y(n_230) );
BUFx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_205), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_SL g243 ( .A(n_205), .Y(n_243) );
INVx4_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_205), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_205), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g619 ( .A(n_205), .B(n_564), .Y(n_619) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g344 ( .A(n_209), .B(n_224), .Y(n_344) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_210), .Y(n_280) );
INVx2_ASAP7_75t_L g298 ( .A(n_210), .Y(n_298) );
AND2x4_ASAP7_75t_L g317 ( .A(n_210), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g405 ( .A(n_210), .Y(n_405) );
INVx2_ASAP7_75t_L g591 ( .A(n_215), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_215), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_SL g251 ( .A(n_217), .Y(n_251) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_225), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_223), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g386 ( .A(n_224), .Y(n_386) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2x1_ASAP7_75t_L g228 ( .A(n_229), .B(n_240), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_229), .B(n_241), .Y(n_336) );
INVx1_ASAP7_75t_L g434 ( .A(n_229), .Y(n_434) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g274 ( .A(n_230), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g288 ( .A(n_230), .B(n_266), .Y(n_288) );
AND2x4_ASAP7_75t_L g311 ( .A(n_230), .B(n_254), .Y(n_311) );
INVx2_ASAP7_75t_L g328 ( .A(n_230), .Y(n_328) );
AND2x2_ASAP7_75t_L g354 ( .A(n_230), .B(n_255), .Y(n_354) );
INVx1_ASAP7_75t_L g419 ( .A(n_230), .Y(n_419) );
INVx2_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_234), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_237), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g379 ( .A(n_240), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_254), .Y(n_240) );
AND2x2_ASAP7_75t_L g345 ( .A(n_241), .B(n_302), .Y(n_345) );
AND2x4_ASAP7_75t_L g361 ( .A(n_241), .B(n_328), .Y(n_361) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g355 ( .A(n_242), .Y(n_355) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_242) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_276) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_248), .B(n_251), .Y(n_244) );
INVx2_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_253), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g287 ( .A(n_254), .Y(n_287) );
INVx3_ASAP7_75t_L g293 ( .A(n_254), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_254), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_254), .B(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g327 ( .A(n_255), .B(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g451 ( .A(n_255), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_277), .A3(n_278), .B1(n_279), .B2(n_281), .B3(n_285), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NOR2x1_ASAP7_75t_L g263 ( .A(n_264), .B(n_274), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g385 ( .A(n_265), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_276), .Y(n_294) );
INVx2_ASAP7_75t_L g302 ( .A(n_266), .Y(n_302) );
INVx1_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_269), .B(n_524), .Y(n_523) );
AO31x2_ASAP7_75t_L g658 ( .A1(n_271), .A2(n_564), .A3(n_659), .B(n_662), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_274), .A2(n_330), .B1(n_333), .B2(n_337), .Y(n_329) );
OR2x2_ASAP7_75t_L g469 ( .A(n_274), .B(n_287), .Y(n_469) );
AND2x4_ASAP7_75t_L g373 ( .A(n_275), .B(n_335), .Y(n_373) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_276), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_277), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g337 ( .A(n_277), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_277), .B(n_313), .Y(n_415) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g388 ( .A(n_279), .Y(n_388) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g446 ( .A(n_282), .B(n_314), .Y(n_446) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_282), .B(n_313), .Y(n_464) );
AND2x2_ASAP7_75t_L g488 ( .A(n_282), .B(n_307), .Y(n_488) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g478 ( .A(n_286), .B(n_355), .Y(n_478) );
NOR2x1p5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g412 ( .A(n_287), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g380 ( .A(n_288), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .B1(n_299), .B2(n_303), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
AND2x2_ASAP7_75t_L g387 ( .A(n_292), .B(n_355), .Y(n_387) );
AND2x2_ASAP7_75t_L g424 ( .A(n_292), .B(n_373), .Y(n_424) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g299 ( .A(n_293), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_293), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g465 ( .A(n_293), .B(n_294), .Y(n_465) );
AND2x2_ASAP7_75t_L g326 ( .A(n_294), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g445 ( .A(n_294), .B(n_311), .Y(n_445) );
AND2x2_ASAP7_75t_L g489 ( .A(n_294), .B(n_354), .Y(n_489) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_299), .A2(n_424), .B1(n_425), .B2(n_428), .C1(n_430), .C2(n_431), .Y(n_423) );
AND2x2_ASAP7_75t_L g346 ( .A(n_300), .B(n_314), .Y(n_346) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g377 ( .A(n_301), .Y(n_377) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_301), .Y(n_422) );
INVx2_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g392 ( .A(n_305), .Y(n_392) );
INVx2_ASAP7_75t_L g398 ( .A(n_306), .Y(n_398) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g382 ( .A(n_307), .B(n_371), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x4_ASAP7_75t_L g413 ( .A(n_310), .B(n_361), .Y(n_413) );
INVx2_ASAP7_75t_L g460 ( .A(n_310), .Y(n_460) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g403 ( .A(n_314), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g437 ( .A(n_314), .B(n_322), .Y(n_437) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_317), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g449 ( .A(n_317), .B(n_365), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_324), .B(n_326), .C(n_329), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
OR2x2_ASAP7_75t_L g330 ( .A(n_322), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g366 ( .A(n_322), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_323), .B(n_358), .Y(n_462) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g438 ( .A(n_325), .B(n_407), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_327), .B(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_327), .A2(n_343), .B1(n_385), .B2(n_387), .Y(n_384) );
AND2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_355), .Y(n_390) );
AND2x2_ASAP7_75t_L g459 ( .A(n_327), .B(n_460), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_330), .A2(n_432), .B(n_453), .C(n_456), .Y(n_452) );
INVx2_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g443 ( .A(n_335), .Y(n_443) );
INVx1_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_337), .A2(n_384), .B1(n_388), .B2(n_389), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_351), .C(n_374), .Y(n_338) );
AO22x1_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B1(n_346), .B2(n_347), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_344), .Y(n_477) );
OR2x2_ASAP7_75t_L g484 ( .A(n_344), .B(n_365), .Y(n_484) );
AND2x2_ASAP7_75t_L g396 ( .A(n_345), .B(n_354), .Y(n_396) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g472 ( .A(n_350), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .C(n_362), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
AND2x4_ASAP7_75t_SL g430 ( .A(n_354), .B(n_373), .Y(n_430) );
INVx1_ASAP7_75t_SL g441 ( .A(n_354), .Y(n_441) );
OR2x2_ASAP7_75t_L g393 ( .A(n_355), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x4_ASAP7_75t_L g370 ( .A(n_358), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g428 ( .A(n_359), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g450 ( .A(n_361), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g475 ( .A(n_361), .B(n_455), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_369), .B2(n_372), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x4_ASAP7_75t_L g410 ( .A(n_366), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g432 ( .A(n_366), .Y(n_432) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g487 ( .A(n_370), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_383), .C(n_391), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_381), .Y(n_375) );
INVx1_ASAP7_75t_L g456 ( .A(n_377), .Y(n_456) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_382), .A2(n_480), .B1(n_483), .B2(n_485), .C1(n_487), .C2(n_489), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_385), .B(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g408 ( .A(n_386), .Y(n_408) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_395), .C(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_457), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_423), .C(n_433), .D(n_444), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_412), .B1(n_414), .B2(n_416), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .C(n_409), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_403), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_407), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g454 ( .A(n_419), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_421), .Y(n_486) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_436), .C(n_442), .Y(n_433) );
AOI21xp33_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_438), .B(n_439), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_437), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_447), .B2(n_450), .C(n_452), .Y(n_444) );
INVx1_ASAP7_75t_L g482 ( .A(n_445), .Y(n_482) );
AOI31xp33_ASAP7_75t_L g466 ( .A1(n_448), .A2(n_467), .A3(n_468), .B(n_469), .Y(n_466) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g455 ( .A(n_451), .Y(n_455) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_470), .C(n_479), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B1(n_463), .B2(n_465), .C(n_466), .Y(n_458) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g467 ( .A(n_465), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B1(n_476), .B2(n_478), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g493 ( .A(n_490), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_494), .B(n_495), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_495), .A2(n_499), .B(n_500), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
NOR2xp67_ASAP7_75t_SL g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_833), .B(n_840), .Y(n_504) );
XNOR2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_731), .Y(n_515) );
NAND3xp33_ASAP7_75t_SL g516 ( .A(n_517), .B(n_634), .C(n_693), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_534), .B1(n_621), .B2(n_627), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g690 ( .A(n_519), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_519), .B(n_608), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_519), .B(n_654), .Y(n_801) );
AND2x2_ASAP7_75t_L g807 ( .A(n_519), .B(n_633), .Y(n_807) );
INVxp67_ASAP7_75t_L g812 ( .A(n_519), .Y(n_812) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g625 ( .A(n_520), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_529), .B(n_532), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_525), .B(n_527), .Y(n_522) );
BUFx4f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_528), .B(n_615), .Y(n_614) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_584), .B(n_594), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_565), .Y(n_536) );
INVx1_ASAP7_75t_L g728 ( .A(n_537), .Y(n_728) );
AND2x2_ASAP7_75t_L g757 ( .A(n_537), .B(n_719), .Y(n_757) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_550), .Y(n_537) );
AND2x2_ASAP7_75t_L g651 ( .A(n_538), .B(n_573), .Y(n_651) );
INVx1_ASAP7_75t_L g706 ( .A(n_538), .Y(n_706) );
AND2x2_ASAP7_75t_L g756 ( .A(n_538), .B(n_572), .Y(n_756) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g631 ( .A(n_539), .B(n_572), .Y(n_631) );
AND2x4_ASAP7_75t_L g775 ( .A(n_539), .B(n_573), .Y(n_775) );
AOI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_545), .B(n_548), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_542), .A2(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g700 ( .A(n_550), .Y(n_700) );
AND2x2_ASAP7_75t_L g769 ( .A(n_550), .B(n_573), .Y(n_769) );
AND2x2_ASAP7_75t_L g776 ( .A(n_550), .B(n_602), .Y(n_776) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g598 ( .A(n_551), .Y(n_598) );
BUFx3_ASAP7_75t_L g633 ( .A(n_551), .Y(n_633) );
AND2x2_ASAP7_75t_L g644 ( .A(n_551), .B(n_630), .Y(n_644) );
AND2x2_ASAP7_75t_L g707 ( .A(n_551), .B(n_566), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_551), .B(n_573), .Y(n_712) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_559), .B(n_562), .Y(n_553) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_565), .B(n_718), .Y(n_820) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_572), .Y(n_565) );
INVx2_ASAP7_75t_L g602 ( .A(n_566), .Y(n_602) );
OR2x2_ASAP7_75t_L g605 ( .A(n_566), .B(n_573), .Y(n_605) );
INVx2_ASAP7_75t_L g630 ( .A(n_566), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_566), .B(n_600), .Y(n_646) );
AND2x2_ASAP7_75t_L g719 ( .A(n_566), .B(n_573), .Y(n_719) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g647 ( .A(n_573), .Y(n_647) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_585), .B(n_682), .Y(n_828) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
AND2x2_ASAP7_75t_L g626 ( .A(n_587), .B(n_608), .Y(n_626) );
INVx1_ASAP7_75t_L g674 ( .A(n_587), .Y(n_674) );
OR2x2_ASAP7_75t_L g679 ( .A(n_587), .B(n_658), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_587), .B(n_658), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_587), .B(n_657), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_587), .B(n_625), .Y(n_764) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_603), .B(n_606), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
OR2x2_ASAP7_75t_L g604 ( .A(n_597), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g755 ( .A(n_597), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g785 ( .A(n_597), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_598), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g753 ( .A(n_598), .Y(n_753) );
OR2x2_ASAP7_75t_L g666 ( .A(n_599), .B(n_667), .Y(n_666) );
INVxp33_ASAP7_75t_L g784 ( .A(n_599), .Y(n_784) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx2_ASAP7_75t_L g688 ( .A(n_600), .Y(n_688) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g750 ( .A1(n_604), .A2(n_675), .B1(n_680), .B2(n_751), .C(n_754), .Y(n_750) );
OR2x2_ASAP7_75t_L g737 ( .A(n_605), .B(n_688), .Y(n_737) );
INVx2_ASAP7_75t_L g786 ( .A(n_605), .Y(n_786) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g686 ( .A(n_607), .Y(n_686) );
OR2x2_ASAP7_75t_L g689 ( .A(n_607), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_607), .Y(n_730) );
OR2x2_ASAP7_75t_L g743 ( .A(n_607), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_620), .Y(n_607) );
NAND2x1p5_ASAP7_75t_SL g639 ( .A(n_608), .B(n_624), .Y(n_639) );
INVx3_ASAP7_75t_L g654 ( .A(n_608), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_608), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g677 ( .A(n_608), .Y(n_677) );
AND2x2_ASAP7_75t_L g758 ( .A(n_608), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g765 ( .A(n_608), .B(n_672), .Y(n_765) );
AND2x4_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_616), .B(n_619), .Y(n_610) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
AND2x2_ASAP7_75t_L g817 ( .A(n_622), .B(n_676), .Y(n_817) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g721 ( .A(n_624), .B(n_691), .Y(n_721) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g656 ( .A(n_625), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g682 ( .A(n_625), .B(n_658), .Y(n_682) );
AND2x4_ASAP7_75t_L g779 ( .A(n_626), .B(n_749), .Y(n_779) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_632), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g698 ( .A(n_631), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_632), .B(n_719), .Y(n_803) );
AND2x2_ASAP7_75t_L g810 ( .A(n_632), .B(n_770), .Y(n_810) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g735 ( .A(n_633), .Y(n_735) );
AOI321xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_648), .A3(n_664), .B1(n_665), .B2(n_668), .C(n_683), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_645), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_641), .B(n_643), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g648 ( .A1(n_638), .A2(n_649), .B(n_652), .Y(n_648) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g747 ( .A(n_639), .B(n_679), .Y(n_747) );
INVx1_ASAP7_75t_L g739 ( .A(n_640), .Y(n_739) );
INVx2_ASAP7_75t_L g724 ( .A(n_641), .Y(n_724) );
OAI32xp33_ASAP7_75t_L g827 ( .A1(n_641), .A2(n_789), .A3(n_800), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g742 ( .A(n_642), .Y(n_742) );
INVx1_ASAP7_75t_L g692 ( .A(n_643), .Y(n_692) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_SL g780 ( .A(n_644), .B(n_687), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_645), .B(n_649), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_645), .A2(n_721), .B1(n_782), .B2(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g770 ( .A(n_646), .Y(n_770) );
INVx1_ASAP7_75t_L g667 ( .A(n_647), .Y(n_667) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g752 ( .A(n_651), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_652), .B(n_669), .C(n_675), .D(n_680), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVxp67_ASAP7_75t_L g694 ( .A(n_653), .Y(n_694) );
AND2x2_ASAP7_75t_L g773 ( .A(n_653), .B(n_682), .Y(n_773) );
OR2x2_ASAP7_75t_L g782 ( .A(n_653), .B(n_656), .Y(n_782) );
AND2x2_ASAP7_75t_L g806 ( .A(n_653), .B(n_678), .Y(n_806) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g720 ( .A(n_654), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g727 ( .A(n_654), .B(n_674), .Y(n_727) );
INVx1_ASAP7_75t_L g791 ( .A(n_655), .Y(n_791) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g699 ( .A(n_656), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g749 ( .A(n_656), .Y(n_749) );
INVx1_ASAP7_75t_L g691 ( .A(n_657), .Y(n_691) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g672 ( .A(n_658), .Y(n_672) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
AND2x4_ASAP7_75t_L g685 ( .A(n_671), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g726 ( .A(n_671), .Y(n_726) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_673), .Y(n_790) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x2_ASAP7_75t_L g681 ( .A(n_677), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g767 ( .A(n_679), .Y(n_767) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g744 ( .A(n_682), .Y(n_744) );
AND2x2_ASAP7_75t_L g787 ( .A(n_682), .B(n_727), .Y(n_787) );
O2A1O1Ixp33_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_687), .B(n_689), .C(n_692), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g798 ( .A(n_687), .B(n_776), .Y(n_798) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g702 ( .A(n_690), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_708), .C(n_722), .Y(n_693) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .B(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_697), .A2(n_805), .B(n_808), .Y(n_804) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g718 ( .A(n_700), .Y(n_718) );
AND2x2_ASAP7_75t_L g778 ( .A(n_700), .B(n_775), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g797 ( .A(n_705), .Y(n_797) );
AND2x2_ASAP7_75t_L g823 ( .A(n_705), .B(n_786), .Y(n_823) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g711 ( .A(n_706), .Y(n_711) );
INVx2_ASAP7_75t_L g762 ( .A(n_707), .Y(n_762) );
NAND2x1_ASAP7_75t_L g796 ( .A(n_707), .B(n_797), .Y(n_796) );
AOI33xp33_ASAP7_75t_L g814 ( .A1(n_707), .A2(n_727), .A3(n_765), .B1(n_775), .B2(n_807), .B3(n_855), .Y(n_814) );
OAI22xp33_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_713), .B1(n_716), .B2(n_720), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g741 ( .A(n_712), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_713), .B(n_800), .Y(n_799) );
OR2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
OR2x2_ASAP7_75t_L g826 ( .A(n_715), .B(n_760), .Y(n_826) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
OAI22xp33_ASAP7_75t_SL g722 ( .A1(n_723), .A2(n_725), .B1(n_728), .B2(n_729), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_726), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_726), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g748 ( .A(n_727), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g813 ( .A(n_727), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_792), .Y(n_731) );
NOR4xp25_ASAP7_75t_L g732 ( .A(n_733), .B(n_750), .C(n_771), .D(n_788), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_738), .B1(n_740), .B2(n_743), .C(n_745), .Y(n_733) );
O2A1O1Ixp33_ASAP7_75t_SL g788 ( .A1(n_734), .A2(n_789), .B(n_790), .C(n_791), .Y(n_788) );
NAND2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g821 ( .A(n_737), .Y(n_821) );
INVx2_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_741), .A2(n_746), .B(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OR2x6_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_757), .B(n_758), .C(n_761), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g800 ( .A(n_760), .B(n_801), .Y(n_800) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_760), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_766), .B2(n_768), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B(n_777), .C(n_783), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_775), .A2(n_823), .B1(n_824), .B2(n_825), .C(n_827), .Y(n_822) );
INVx3_ASAP7_75t_L g830 ( .A(n_775), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_777) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI21xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B(n_787), .Y(n_783) );
INVx1_ASAP7_75t_L g789 ( .A(n_786), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_815), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_804), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_798), .B(n_799), .C(n_802), .Y(n_794) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_798), .B(n_819), .C(n_821), .Y(n_818) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_811), .B(n_814), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OR2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_818), .B(n_822), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
AND2x2_ASAP7_75t_L g846 ( .A(n_832), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx5_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AND2x6_ASAP7_75t_SL g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
INVx6_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
BUFx10_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx5_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
endmodule