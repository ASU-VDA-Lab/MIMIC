module fake_ariane_1156_n_1720 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1720);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1720;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_42),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_11),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_47),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_14),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_63),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_0),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_55),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_35),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_13),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_23),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_53),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_112),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_54),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_94),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_23),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_109),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_31),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_33),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_88),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_126),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_99),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_83),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_27),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_106),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_33),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_41),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_9),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_67),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_2),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_79),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_46),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_21),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_104),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_115),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_129),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_61),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_19),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_15),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_59),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_11),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_40),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_39),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_66),
.Y(n_217)
);

INVx4_ASAP7_75t_R g218 ( 
.A(n_122),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_76),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_114),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_120),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_7),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_90),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g228 ( 
.A(n_118),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_10),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_8),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_43),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_8),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_93),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_37),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_26),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_27),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_75),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_34),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_18),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_111),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_69),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_16),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_124),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_102),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_0),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_16),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_135),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_6),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_65),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_84),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_70),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_132),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_96),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_39),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_22),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_100),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_34),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_131),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_128),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_143),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_42),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_82),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_64),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_45),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_38),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_68),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_3),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_101),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_108),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_71),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_72),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_37),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_12),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_77),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_56),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_146),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_29),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_73),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_152),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_170),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_169),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_197),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_200),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_202),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_163),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_206),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_242),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_276),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_175),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_201),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_193),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_194),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_201),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_201),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_190),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_157),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_225),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_237),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_148),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_178),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_180),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_187),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_195),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_208),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_243),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_154),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_275),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_149),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_279),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_154),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_155),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_155),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_182),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_182),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_149),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_151),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_196),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_196),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_151),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_252),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_289),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_214),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_219),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_158),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_158),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_239),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_160),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_203),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_160),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_241),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_248),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_307),
.B(n_252),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_277),
.B1(n_162),
.B2(n_284),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_228),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_296),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_309),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_159),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_297),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_321),
.B(n_162),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_189),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_326),
.B(n_251),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_306),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_298),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_298),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_304),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_299),
.A2(n_198),
.B(n_191),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_359),
.A2(n_166),
.B1(n_164),
.B2(n_211),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_303),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_303),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_307),
.B(n_278),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_210),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_343),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

AND3x2_ASAP7_75t_L g409 ( 
.A(n_312),
.B(n_185),
.C(n_292),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_317),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_305),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_308),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_320),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_334),
.B(n_153),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_322),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_342),
.B(n_227),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_316),
.B(n_167),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_310),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_326),
.B(n_245),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_363),
.A2(n_290),
.B1(n_277),
.B2(n_281),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_351),
.A2(n_294),
.B1(n_300),
.B2(n_335),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_347),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_347),
.A2(n_256),
.B(n_246),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_318),
.B(n_265),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_319),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_348),
.B(n_163),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_430),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_371),
.A2(n_281),
.B1(n_284),
.B2(n_286),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_370),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_356),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_398),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_381),
.B(n_333),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_398),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_400),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

XOR2x2_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_330),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_398),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_327),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_357),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_395),
.B(n_362),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_420),
.B(n_153),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

AO22x2_ASAP7_75t_L g470 ( 
.A1(n_368),
.A2(n_422),
.B1(n_385),
.B2(n_366),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_404),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_368),
.A2(n_286),
.B1(n_287),
.B2(n_255),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_416),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_367),
.B(n_349),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_369),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_372),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_372),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_432),
.B(n_406),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_425),
.B(n_156),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_375),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_425),
.B(n_156),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_417),
.B(n_353),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_375),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_376),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_376),
.A2(n_282),
.B(n_270),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_410),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_429),
.A2(n_355),
.B1(n_352),
.B2(n_354),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_388),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_407),
.Y(n_502)
);

OR2x6_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_360),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_423),
.A2(n_287),
.B1(n_204),
.B2(n_205),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_389),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_422),
.B(n_360),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_383),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_390),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_370),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_427),
.B(n_364),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

OAI22xp33_ASAP7_75t_L g522 ( 
.A1(n_423),
.A2(n_271),
.B1(n_212),
.B2(n_215),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_374),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_378),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_394),
.A2(n_261),
.B1(n_253),
.B2(n_224),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_427),
.B(n_350),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_427),
.B(n_350),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_427),
.B(n_364),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_422),
.B(n_352),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_424),
.B(n_426),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_407),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_385),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_385),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_407),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_391),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_394),
.B(n_328),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_424),
.B(n_365),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_434),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_434),
.Y(n_544)
);

NOR3xp33_ASAP7_75t_L g545 ( 
.A(n_379),
.B(n_266),
.C(n_235),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_408),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_385),
.A2(n_268),
.B1(n_216),
.B2(n_229),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_426),
.B(n_354),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_434),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_393),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_411),
.B(n_161),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_412),
.B(n_165),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_378),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_329),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_421),
.B(n_165),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_405),
.B(n_331),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_431),
.B(n_332),
.Y(n_558)
);

AOI21x1_ASAP7_75t_L g559 ( 
.A1(n_393),
.A2(n_291),
.B(n_285),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_434),
.B(n_220),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_408),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_405),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_384),
.B(n_220),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_408),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_384),
.B(n_274),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_429),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_429),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_408),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_429),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_409),
.Y(n_571)
);

BUFx6f_ASAP7_75t_SL g572 ( 
.A(n_433),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_408),
.Y(n_573)
);

INVx8_ASAP7_75t_L g574 ( 
.A(n_433),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_382),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_408),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_418),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_401),
.B(n_311),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_401),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_379),
.B(n_274),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_393),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_484),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_443),
.A2(n_280),
.B1(n_283),
.B2(n_288),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_462),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_448),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_463),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_462),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_448),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_451),
.B(n_461),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_470),
.A2(n_393),
.B1(n_433),
.B2(n_336),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_462),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_280),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_494),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_494),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_449),
.B(n_283),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_524),
.B(n_288),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_443),
.A2(n_314),
.B1(n_183),
.B2(n_293),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_487),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_487),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_447),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_509),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_554),
.B(n_409),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_435),
.B(n_382),
.Y(n_605)
);

OAI221xp5_ASAP7_75t_L g606 ( 
.A1(n_504),
.A2(n_231),
.B1(n_232),
.B2(n_264),
.C(n_233),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_562),
.B(n_240),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_460),
.B(n_415),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_562),
.B(n_244),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_465),
.B(n_263),
.Y(n_611)
);

INVxp33_ASAP7_75t_L g612 ( 
.A(n_458),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_460),
.B(n_415),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_513),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_519),
.B(n_168),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_435),
.B(n_455),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_578),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_513),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_519),
.B(n_171),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_435),
.B(n_172),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_455),
.B(n_1),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_435),
.B(n_173),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_535),
.B(n_174),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_439),
.B(n_456),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_531),
.B(n_564),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_531),
.B(n_176),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_177),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_557),
.B(n_179),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_535),
.B(n_1),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_477),
.A2(n_336),
.B(n_340),
.C(n_373),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_477),
.A2(n_340),
.B(n_373),
.C(n_377),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_537),
.B(n_181),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_537),
.B(n_184),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_447),
.B(n_323),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_457),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_472),
.B(n_163),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_557),
.B(n_186),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_515),
.B(n_3),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_484),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_506),
.B(n_188),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_447),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_515),
.B(n_5),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_457),
.Y(n_644)
);

NOR3xp33_ASAP7_75t_L g645 ( 
.A(n_486),
.B(n_339),
.C(n_337),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_515),
.B(n_5),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_464),
.Y(n_647)
);

INVxp33_ASAP7_75t_L g648 ( 
.A(n_458),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_R g649 ( 
.A(n_539),
.B(n_325),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_464),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_472),
.A2(n_418),
.B1(n_223),
.B2(n_221),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_466),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_443),
.A2(n_262),
.B1(n_236),
.B2(n_192),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_447),
.B(n_418),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_515),
.B(n_12),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_493),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_466),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_523),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_447),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_504),
.A2(n_254),
.B1(n_217),
.B2(n_213),
.C(n_209),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g661 ( 
.A1(n_522),
.A2(n_207),
.B1(n_273),
.B2(n_269),
.C(n_230),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_571),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_443),
.B(n_260),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_506),
.B(n_267),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_478),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_515),
.B(n_15),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_491),
.B(n_17),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_478),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_506),
.B(n_259),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_525),
.B(n_418),
.C(n_249),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_449),
.B(n_19),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_506),
.B(n_418),
.Y(n_674)
);

BUFx5_ASAP7_75t_L g675 ( 
.A(n_550),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_540),
.B(n_418),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_449),
.B(n_20),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_482),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_571),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_470),
.A2(n_433),
.B1(n_163),
.B2(n_222),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_540),
.B(n_234),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_474),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_533),
.B(n_247),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_547),
.B(n_20),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_439),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_449),
.B(n_250),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_493),
.A2(n_496),
.B1(n_479),
.B2(n_485),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_503),
.B(n_558),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_450),
.B(n_250),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_503),
.B(n_433),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_550),
.B(n_163),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_474),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_575),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_503),
.B(n_373),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_503),
.B(n_377),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_547),
.B(n_24),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_450),
.B(n_24),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_492),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_439),
.B(n_257),
.Y(n_699)
);

INVx8_ASAP7_75t_L g700 ( 
.A(n_463),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_541),
.B(n_392),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_467),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_571),
.B(n_222),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_492),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_450),
.B(n_25),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_571),
.B(n_468),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_541),
.B(n_392),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_470),
.A2(n_222),
.B1(n_257),
.B2(n_250),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_580),
.B(n_25),
.C(n_28),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_467),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_450),
.B(n_29),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_475),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_470),
.A2(n_257),
.B1(n_250),
.B2(n_222),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_545),
.B(n_30),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_493),
.B(n_250),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_453),
.B(n_30),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_453),
.B(n_250),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_453),
.B(n_250),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_474),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_442),
.B(n_31),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_550),
.A2(n_222),
.B1(n_257),
.B2(n_380),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_453),
.B(n_459),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_459),
.B(n_32),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_459),
.B(n_552),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_459),
.B(n_380),
.C(n_396),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_553),
.B(n_556),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_498),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_488),
.B(n_32),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_479),
.B(n_257),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_507),
.B(n_35),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_439),
.B(n_36),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_485),
.A2(n_380),
.B(n_396),
.C(n_40),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_489),
.B(n_257),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_498),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_490),
.B(n_512),
.C(n_501),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_489),
.B(n_257),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_456),
.B(n_257),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_499),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_499),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_496),
.A2(n_36),
.B1(n_38),
.B2(n_43),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_475),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_581),
.A2(n_380),
.B1(n_396),
.B2(n_218),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_501),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_510),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_505),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_505),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_532),
.B(n_44),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_589),
.B(n_555),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_649),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_675),
.B(n_456),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_658),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_637),
.A2(n_456),
.B1(n_469),
.B2(n_520),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_700),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_637),
.A2(n_500),
.B1(n_495),
.B2(n_581),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_585),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_602),
.B(n_469),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_700),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_613),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_588),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_589),
.B(n_469),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_700),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_600),
.B(n_548),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_617),
.B(n_469),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_668),
.B(n_508),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_636),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_644),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_668),
.B(n_611),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_675),
.B(n_508),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_611),
.B(n_512),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_649),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_647),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_675),
.B(n_516),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_601),
.B(n_527),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_675),
.B(n_516),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_666),
.B(n_529),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_587),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_650),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_652),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_587),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_682),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_635),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_676),
.B(n_518),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_675),
.B(n_642),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_708),
.A2(n_495),
.B1(n_581),
.B2(n_568),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_675),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_657),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_702),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_626),
.B(n_688),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_659),
.B(n_518),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_639),
.A2(n_520),
.B(n_476),
.C(n_471),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_722),
.B(n_582),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_693),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_SL g795 ( 
.A1(n_684),
.A2(n_495),
.B1(n_572),
.B2(n_511),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_607),
.B(n_610),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_722),
.B(n_474),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_621),
.B(n_440),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_674),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_591),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_662),
.B(n_440),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_710),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_639),
.A2(n_473),
.B(n_454),
.C(n_471),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_712),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_621),
.B(n_593),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_609),
.B(n_436),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_679),
.B(n_463),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_591),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_604),
.B(n_445),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_741),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_743),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_643),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_745),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_746),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_592),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_708),
.A2(n_568),
.B1(n_567),
.B2(n_570),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_586),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_599),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_592),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_696),
.A2(n_651),
.B1(n_646),
.B2(n_643),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_646),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_682),
.Y(n_822)
);

AND2x6_ASAP7_75t_L g823 ( 
.A(n_713),
.B(n_567),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_594),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_730),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_594),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_616),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_SL g828 ( 
.A1(n_606),
.A2(n_511),
.B1(n_570),
.B2(n_445),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_701),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_682),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_645),
.B(n_436),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_707),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_654),
.B(n_438),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_582),
.B(n_474),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_598),
.B(n_437),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_640),
.B(n_474),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_586),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_720),
.B(n_437),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_595),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_595),
.Y(n_840)
);

AND2x6_ASAP7_75t_SL g841 ( 
.A(n_714),
.B(n_655),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_640),
.A2(n_473),
.B1(n_452),
.B2(n_454),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_656),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_596),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_655),
.A2(n_560),
.B1(n_511),
.B2(n_452),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_596),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_682),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_603),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_683),
.B(n_444),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_603),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_656),
.B(n_673),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_615),
.B(n_438),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_667),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_441),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_608),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_681),
.B(n_441),
.Y(n_856)
);

INVx6_ASAP7_75t_L g857 ( 
.A(n_692),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_619),
.B(n_441),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_608),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_673),
.B(n_481),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_614),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_612),
.B(n_446),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_667),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_627),
.B(n_630),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_648),
.B(n_446),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_677),
.B(n_481),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_692),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_630),
.B(n_446),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_663),
.B(n_511),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_614),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_583),
.B(n_521),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_605),
.B(n_510),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_692),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_SL g874 ( 
.A(n_660),
.B(n_572),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_714),
.B(n_514),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_726),
.B(n_521),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_664),
.B(n_526),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_618),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_747),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_747),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_SL g881 ( 
.A1(n_680),
.A2(n_528),
.B1(n_536),
.B2(n_526),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_618),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_623),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_623),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_728),
.B(n_544),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_661),
.A2(n_528),
.B1(n_536),
.B2(n_543),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_677),
.B(n_542),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_697),
.B(n_542),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_665),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_671),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_669),
.Y(n_891)
);

BUFx10_ASAP7_75t_L g892 ( 
.A(n_697),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_705),
.B(n_517),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_692),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_680),
.B(n_544),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_705),
.B(n_711),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_711),
.B(n_517),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_669),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_670),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_719),
.B(n_563),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_590),
.A2(n_514),
.B1(n_549),
.B2(n_551),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_SL g902 ( 
.A(n_740),
.B(n_543),
.C(n_47),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_670),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_590),
.A2(n_549),
.B1(n_551),
.B2(n_574),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_678),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_678),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_698),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_719),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_629),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_704),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_SL g911 ( 
.A(n_620),
.B(n_622),
.C(n_641),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_704),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_727),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_719),
.B(n_690),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_716),
.B(n_538),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_727),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_719),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_716),
.B(n_538),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_724),
.B(n_563),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_734),
.A2(n_463),
.B1(n_574),
.B2(n_572),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_734),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_738),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_723),
.B(n_497),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_687),
.A2(n_546),
.B1(n_480),
.B2(n_534),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_738),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_723),
.B(n_628),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_694),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_731),
.B(n_497),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_739),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_731),
.B(n_497),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_597),
.B(n_497),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_685),
.B(n_538),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_739),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_757),
.B(n_703),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_768),
.B(n_638),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_760),
.A2(n_625),
.B(n_699),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_896),
.A2(n_709),
.B(n_633),
.C(n_624),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_790),
.B(n_744),
.Y(n_938)
);

AOI33xp33_ASAP7_75t_L g939 ( 
.A1(n_763),
.A2(n_653),
.A3(n_631),
.B1(n_632),
.B2(n_744),
.B3(n_51),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_748),
.B(n_691),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_765),
.B(n_691),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_749),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_812),
.B(n_672),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_758),
.B(n_695),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_853),
.B(n_794),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_821),
.B(n_634),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_765),
.A2(n_721),
.B1(n_597),
.B2(n_742),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_896),
.A2(n_732),
.B(n_686),
.C(n_689),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_751),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_796),
.A2(n_689),
.B(n_686),
.C(n_736),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_751),
.B(n_783),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_805),
.B(n_926),
.C(n_864),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_863),
.B(n_691),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_892),
.B(n_481),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_776),
.A2(n_717),
.B(n_718),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_829),
.B(n_691),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_892),
.B(n_497),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_762),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_772),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_862),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_806),
.B(n_480),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_887),
.A2(n_737),
.B(n_733),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_775),
.B(n_561),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_762),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_782),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_909),
.B(n_737),
.Y(n_966)
);

O2A1O1Ixp5_ASAP7_75t_L g967 ( 
.A1(n_860),
.A2(n_729),
.B(n_715),
.C(n_725),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_799),
.B(n_546),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_902),
.A2(n_538),
.B(n_483),
.C(n_573),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_888),
.A2(n_546),
.B(n_480),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_893),
.A2(n_546),
.B(n_480),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_799),
.B(n_483),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_792),
.A2(n_561),
.B(n_502),
.C(n_573),
.Y(n_973)
);

OAI22x1_ASAP7_75t_L g974 ( 
.A1(n_879),
.A2(n_559),
.B1(n_576),
.B2(n_577),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_890),
.B(n_791),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_825),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_897),
.A2(n_561),
.B(n_483),
.Y(n_977)
);

INVxp33_ASAP7_75t_L g978 ( 
.A(n_865),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_791),
.A2(n_481),
.B1(n_497),
.B2(n_561),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_792),
.A2(n_534),
.B(n_502),
.C(n_573),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_827),
.A2(n_483),
.B(n_502),
.C(n_530),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_880),
.B(n_573),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_791),
.A2(n_481),
.B1(n_502),
.B2(n_530),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_SL g984 ( 
.A1(n_825),
.A2(n_577),
.B1(n_576),
.B2(n_569),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_841),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_871),
.A2(n_481),
.B1(n_534),
.B2(n_530),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_R g987 ( 
.A(n_762),
.B(n_559),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_832),
.B(n_530),
.Y(n_988)
);

OA21x2_ASAP7_75t_L g989 ( 
.A1(n_928),
.A2(n_569),
.B(n_565),
.Y(n_989)
);

OAI22x1_ASAP7_75t_L g990 ( 
.A1(n_831),
.A2(n_875),
.B1(n_789),
.B2(n_788),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_838),
.B(n_565),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_860),
.A2(n_565),
.B(n_48),
.C(n_49),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_777),
.B(n_45),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_915),
.A2(n_565),
.B(n_574),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_757),
.B(n_565),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_918),
.A2(n_565),
.B(n_574),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_755),
.B(n_759),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_770),
.A2(n_774),
.B(n_750),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_766),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_784),
.B(n_574),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_787),
.A2(n_463),
.B(n_563),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_762),
.B(n_563),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_767),
.B(n_773),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_L g1004 ( 
.A(n_827),
.B(n_48),
.C(n_50),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_764),
.B(n_50),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_779),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_780),
.B(n_802),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_782),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_793),
.A2(n_563),
.B(n_396),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_833),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_804),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_891),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_810),
.B(n_52),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_793),
.A2(n_563),
.B(n_396),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_851),
.A2(n_396),
.B(n_380),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_811),
.B(n_813),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_814),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_851),
.A2(n_57),
.B(n_58),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_SL g1019 ( 
.A1(n_752),
.A2(n_74),
.B(n_78),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_881),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_876),
.A2(n_95),
.B(n_110),
.C(n_117),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_833),
.B(n_119),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_889),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_898),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_928),
.A2(n_930),
.B(n_770),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_872),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_930),
.A2(n_133),
.B(n_138),
.Y(n_1027)
);

BUFx8_ASAP7_75t_SL g1028 ( 
.A(n_782),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_843),
.B(n_876),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_843),
.B(n_854),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_911),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_L g1032 ( 
.A(n_828),
.B(n_931),
.C(n_803),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_927),
.B(n_895),
.Y(n_1033)
);

AO32x1_ASAP7_75t_L g1034 ( 
.A1(n_924),
.A2(n_842),
.A3(n_861),
.B1(n_870),
.B2(n_878),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_895),
.B(n_756),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_774),
.A2(n_923),
.B(n_866),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_782),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_754),
.A2(n_798),
.B1(n_786),
.B2(n_868),
.Y(n_1038)
);

CKINVDCx14_ASAP7_75t_R g1039 ( 
.A(n_857),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_807),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_761),
.B(n_769),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_866),
.A2(n_923),
.B(n_750),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_761),
.B(n_769),
.Y(n_1043)
);

AND2x4_ASAP7_75t_SL g1044 ( 
.A(n_807),
.B(n_756),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_931),
.A2(n_797),
.B(n_803),
.C(n_834),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_807),
.B(n_914),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_877),
.A2(n_845),
.B(n_809),
.C(n_869),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_877),
.A2(n_856),
.B(n_801),
.C(n_849),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_778),
.B(n_781),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_795),
.A2(n_754),
.B1(n_786),
.B2(n_904),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_899),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_835),
.A2(n_858),
.B(n_852),
.C(n_797),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_903),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_895),
.B(n_756),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_904),
.A2(n_816),
.B1(n_886),
.B2(n_932),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_885),
.B(n_854),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_905),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_906),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_834),
.A2(n_836),
.B(n_817),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_914),
.B(n_856),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_836),
.A2(n_817),
.B(n_837),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_837),
.A2(n_785),
.B(n_822),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_907),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_785),
.A2(n_826),
.B(n_778),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_753),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_822),
.A2(n_908),
.B(n_894),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_816),
.A2(n_857),
.B1(n_901),
.B2(n_885),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_922),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_857),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_847),
.B(n_867),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_856),
.A2(n_874),
.B(n_885),
.C(n_882),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_873),
.A2(n_859),
.B(n_848),
.C(n_846),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_952),
.A2(n_936),
.B(n_941),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_994),
.A2(n_824),
.B(n_781),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_1028),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_976),
.Y(n_1076)
);

AO21x2_ASAP7_75t_L g1077 ( 
.A1(n_1038),
.A2(n_883),
.B(n_884),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_1035),
.B(n_914),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_935),
.A2(n_873),
.B(n_840),
.C(n_847),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_1040),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_1038),
.A2(n_844),
.A3(n_800),
.B(n_808),
.Y(n_1081)
);

AOI221x1_ASAP7_75t_L g1082 ( 
.A1(n_1020),
.A2(n_933),
.B1(n_910),
.B2(n_912),
.C(n_913),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_942),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_941),
.A2(n_830),
.B(n_908),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1029),
.B(n_946),
.Y(n_1085)
);

AOI211x1_ASAP7_75t_L g1086 ( 
.A1(n_1007),
.A2(n_925),
.B(n_916),
.C(n_921),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_996),
.A2(n_844),
.B(n_800),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_SL g1088 ( 
.A1(n_1020),
.A2(n_850),
.B(n_808),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_937),
.A2(n_867),
.B(n_815),
.C(n_819),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1003),
.B(n_850),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_938),
.B(n_823),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1047),
.A2(n_908),
.B(n_894),
.Y(n_1092)
);

AO21x1_ASAP7_75t_L g1093 ( 
.A1(n_947),
.A2(n_855),
.B(n_815),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1016),
.B(n_819),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_965),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_955),
.A2(n_947),
.B(n_940),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_949),
.B(n_894),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1042),
.A2(n_824),
.B(n_826),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_940),
.A2(n_901),
.B(n_823),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_1040),
.B(n_822),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1025),
.A2(n_839),
.B(n_929),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_998),
.A2(n_839),
.B(n_929),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_962),
.A2(n_1048),
.B(n_1052),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1026),
.B(n_823),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1045),
.A2(n_920),
.B(n_823),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_974),
.A2(n_823),
.A3(n_919),
.B(n_920),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_960),
.B(n_822),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_1039),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1004),
.A2(n_753),
.B(n_919),
.C(n_900),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_951),
.B(n_830),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1036),
.A2(n_830),
.B(n_894),
.Y(n_1111)
);

NAND2x1_ASAP7_75t_L g1112 ( 
.A(n_965),
.B(n_908),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_SL g1113 ( 
.A1(n_1071),
.A2(n_917),
.B(n_900),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_L g1114 ( 
.A(n_1032),
.B(n_917),
.C(n_1005),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_999),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_950),
.A2(n_917),
.B(n_1000),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1031),
.B(n_945),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_948),
.A2(n_980),
.B(n_973),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1000),
.A2(n_1055),
.B(n_938),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_978),
.B(n_959),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_944),
.B(n_1006),
.Y(n_1121)
);

NAND2x1p5_ASAP7_75t_L g1122 ( 
.A(n_1046),
.B(n_1060),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1013),
.A2(n_1055),
.B(n_993),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1061),
.A2(n_1059),
.B(n_970),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_L g1125 ( 
.A1(n_943),
.A2(n_954),
.B(n_957),
.C(n_992),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_939),
.B(n_1019),
.C(n_1021),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_SL g1127 ( 
.A1(n_963),
.A2(n_988),
.B(n_961),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1011),
.B(n_1017),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1023),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_989),
.A2(n_1062),
.B(n_977),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_968),
.B(n_972),
.Y(n_1131)
);

XOR2xp5_ASAP7_75t_L g1132 ( 
.A(n_985),
.B(n_990),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1067),
.A2(n_1022),
.B(n_1072),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_SL g1134 ( 
.A1(n_1066),
.A2(n_988),
.B(n_969),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_965),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1054),
.B(n_1046),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_989),
.A2(n_971),
.B(n_956),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_SL g1138 ( 
.A(n_1008),
.B(n_1037),
.Y(n_1138)
);

AOI211x1_ASAP7_75t_L g1139 ( 
.A1(n_975),
.A2(n_1057),
.B(n_1063),
.C(n_1058),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1064),
.A2(n_967),
.B(n_1015),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1010),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1024),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1030),
.A2(n_966),
.B1(n_1044),
.B2(n_1050),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1051),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_956),
.A2(n_953),
.B(n_995),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1053),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1069),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_982),
.B(n_972),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_968),
.B(n_1008),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_981),
.A2(n_1018),
.B(n_1027),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1009),
.A2(n_1014),
.B(n_1041),
.Y(n_1151)
);

INVx6_ASAP7_75t_L g1152 ( 
.A(n_958),
.Y(n_1152)
);

NAND3x1_ASAP7_75t_L g1153 ( 
.A(n_1070),
.B(n_964),
.C(n_1033),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_986),
.A2(n_979),
.B(n_983),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_958),
.Y(n_1155)
);

AO32x2_ASAP7_75t_L g1156 ( 
.A1(n_984),
.A2(n_1034),
.A3(n_987),
.B1(n_1056),
.B2(n_1068),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1034),
.A2(n_1001),
.B(n_1049),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_SL g1158 ( 
.A1(n_991),
.A2(n_1065),
.B1(n_1049),
.B2(n_1043),
.C(n_1041),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1012),
.A2(n_1002),
.B(n_1065),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_934),
.A2(n_996),
.B(n_994),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1037),
.B(n_934),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_935),
.B(n_617),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_997),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_997),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_935),
.B(n_617),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_951),
.B(n_539),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_952),
.B(n_790),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1038),
.A2(n_974),
.A3(n_1047),
.B(n_947),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_935),
.B(n_617),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_941),
.A2(n_768),
.B(n_926),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_949),
.Y(n_1171)
);

AO32x2_ASAP7_75t_L g1172 ( 
.A1(n_1050),
.A2(n_1038),
.A3(n_1055),
.B1(n_1020),
.B2(n_1067),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_947),
.A2(n_768),
.B(n_896),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_SL g1174 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1071),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_994),
.A2(n_996),
.B(n_1042),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1028),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_935),
.B(n_617),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_997),
.Y(n_1178)
);

AOI211x1_ASAP7_75t_L g1179 ( 
.A1(n_1007),
.A2(n_606),
.B(n_696),
.C(n_684),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_935),
.B(n_617),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_947),
.A2(n_768),
.B(n_896),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_SL g1182 ( 
.A1(n_941),
.A2(n_768),
.B(n_926),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_947),
.A2(n_768),
.B(n_896),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_1045),
.A2(n_1036),
.B(n_1042),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_997),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_952),
.B(n_768),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_952),
.A2(n_896),
.B(n_768),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_947),
.A2(n_768),
.B(n_896),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1038),
.A2(n_974),
.A3(n_1047),
.B(n_947),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_935),
.B(n_617),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_947),
.A2(n_768),
.B(n_896),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_935),
.A2(n_768),
.B1(n_637),
.B2(n_820),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_SL g1193 ( 
.A1(n_1020),
.A2(n_937),
.B(n_1062),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_935),
.B(n_617),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_951),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_947),
.A2(n_768),
.B(n_896),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_994),
.A2(n_996),
.B(n_1042),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_997),
.B(n_758),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_997),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1031),
.A2(n_768),
.B1(n_820),
.B2(n_447),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_L g1201 ( 
.A(n_1004),
.B(n_768),
.C(n_765),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_SL g1202 ( 
.A1(n_943),
.A2(n_896),
.B(n_866),
.C(n_860),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_994),
.A2(n_996),
.B(n_1042),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1028),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1045),
.A2(n_1036),
.B(n_1042),
.Y(n_1205)
);

AOI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_941),
.A2(n_768),
.B(n_926),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1038),
.A2(n_974),
.A3(n_1047),
.B(n_947),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_994),
.A2(n_996),
.B(n_1042),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_997),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_935),
.B(n_617),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_L g1211 ( 
.A(n_951),
.B(n_539),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_994),
.A2(n_996),
.B(n_1042),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1192),
.A2(n_1201),
.B1(n_1188),
.B2(n_1173),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1128),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1192),
.A2(n_1172),
.B1(n_1201),
.B2(n_1126),
.Y(n_1215)
);

INVx8_ASAP7_75t_L g1216 ( 
.A(n_1075),
.Y(n_1216)
);

OAI211xp5_ASAP7_75t_L g1217 ( 
.A1(n_1123),
.A2(n_1180),
.B(n_1210),
.C(n_1177),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1077),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1130),
.A2(n_1140),
.B(n_1175),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1173),
.A2(n_1183),
.B(n_1181),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1115),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1197),
.A2(n_1208),
.B(n_1203),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1167),
.B(n_1123),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1179),
.B(n_1186),
.C(n_1114),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1198),
.B(n_1163),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1129),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1164),
.B(n_1178),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1075),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1093),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1167),
.B(n_1187),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1212),
.A2(n_1160),
.B(n_1124),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1090),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1181),
.A2(n_1191),
.B(n_1183),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1188),
.B(n_1191),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1137),
.A2(n_1151),
.B(n_1103),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1185),
.B(n_1199),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1157),
.A2(n_1088),
.B(n_1077),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1073),
.A2(n_1111),
.B(n_1096),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1075),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1200),
.A2(n_1194),
.B1(n_1190),
.B2(n_1165),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1136),
.B(n_1110),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1126),
.A2(n_1132),
.B1(n_1114),
.B2(n_1196),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1196),
.B(n_1169),
.C(n_1162),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1074),
.A2(n_1087),
.B(n_1150),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1142),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1116),
.A2(n_1102),
.B(n_1101),
.Y(n_1246)
);

BUFx2_ASAP7_75t_SL g1247 ( 
.A(n_1083),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1091),
.B(n_1119),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1085),
.B(n_1117),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1209),
.B(n_1195),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1108),
.B(n_1147),
.Y(n_1251)
);

AOI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1082),
.A2(n_1092),
.B(n_1193),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1195),
.B(n_1121),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1144),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1146),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1143),
.A2(n_1172),
.B1(n_1091),
.B2(n_1099),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1104),
.B(n_1136),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1098),
.A2(n_1127),
.B(n_1134),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1174),
.A2(n_1118),
.B(n_1133),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1204),
.Y(n_1260)
);

BUFx2_ASAP7_75t_R g1261 ( 
.A(n_1148),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1202),
.A2(n_1118),
.B(n_1125),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1094),
.B(n_1158),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1120),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1139),
.Y(n_1265)
);

AOI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1145),
.A2(n_1084),
.B(n_1097),
.Y(n_1266)
);

OAI211xp5_ASAP7_75t_L g1267 ( 
.A1(n_1166),
.A2(n_1211),
.B(n_1154),
.C(n_1176),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1158),
.B(n_1078),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1078),
.B(n_1168),
.Y(n_1269)
);

AO21x1_ASAP7_75t_L g1270 ( 
.A1(n_1079),
.A2(n_1099),
.B(n_1159),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1095),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1204),
.Y(n_1272)
);

AOI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1154),
.A2(n_1105),
.B(n_1109),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1089),
.A2(n_1131),
.B(n_1107),
.C(n_1149),
.Y(n_1274)
);

AND2x4_ASAP7_75t_SL g1275 ( 
.A(n_1135),
.B(n_1095),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1086),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1161),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1152),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1172),
.A2(n_1105),
.B1(n_1122),
.B2(n_1159),
.Y(n_1279)
);

INVx8_ASAP7_75t_L g1280 ( 
.A(n_1155),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1122),
.A2(n_1152),
.B1(n_1205),
.B2(n_1184),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1170),
.A2(n_1182),
.B(n_1206),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1138),
.A2(n_1155),
.B(n_1189),
.C(n_1168),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1153),
.A2(n_1100),
.B1(n_1135),
.B2(n_1112),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1113),
.A2(n_1205),
.B(n_1184),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1081),
.A2(n_1168),
.B(n_1189),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1081),
.A2(n_1189),
.B(n_1207),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1207),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1207),
.A2(n_1156),
.B(n_1106),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1156),
.A2(n_1093),
.A3(n_1082),
.B(n_1038),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1106),
.A2(n_1130),
.B(n_1140),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1156),
.A2(n_768),
.B(n_1192),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1077),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1128),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1200),
.A2(n_1192),
.B1(n_818),
.B2(n_768),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1130),
.A2(n_1140),
.B(n_1175),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1192),
.A2(n_637),
.B1(n_820),
.B2(n_768),
.Y(n_1297)
);

AOI221x1_ASAP7_75t_L g1298 ( 
.A1(n_1192),
.A2(n_1004),
.B1(n_1201),
.B2(n_768),
.C(n_1020),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1093),
.A2(n_1082),
.A3(n_1038),
.B(n_1157),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_SL g1300 ( 
.A1(n_1173),
.A2(n_1183),
.B(n_1181),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1141),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1200),
.A2(n_1192),
.B1(n_818),
.B2(n_768),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1192),
.A2(n_768),
.B(n_1201),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1167),
.B(n_1123),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1192),
.A2(n_637),
.B1(n_820),
.B2(n_768),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1157),
.A2(n_1088),
.B(n_1093),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1186),
.A2(n_768),
.B(n_1201),
.C(n_1165),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1075),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1173),
.A2(n_896),
.B(n_1181),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1082),
.A2(n_1096),
.B(n_1175),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1075),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1200),
.A2(n_637),
.B1(n_1050),
.B2(n_648),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1128),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1192),
.A2(n_637),
.B1(n_820),
.B2(n_768),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1141),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1075),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1171),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1130),
.A2(n_1140),
.B(n_1175),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1130),
.A2(n_1140),
.B(n_1175),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1130),
.A2(n_1140),
.B(n_1175),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1171),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1200),
.A2(n_637),
.B1(n_1050),
.B2(n_648),
.Y(n_1322)
);

INVx3_ASAP7_75t_SL g1323 ( 
.A(n_1076),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1080),
.B(n_1040),
.Y(n_1324)
);

NAND2xp33_ASAP7_75t_R g1325 ( 
.A(n_1076),
.B(n_649),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1171),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1082),
.A2(n_1137),
.B(n_1130),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1075),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1082),
.A2(n_1137),
.B(n_1130),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1083),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_SL g1331 ( 
.A1(n_1186),
.A2(n_768),
.B(n_1201),
.C(n_1165),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1288),
.B(n_1223),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1214),
.B(n_1294),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1221),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1288),
.B(n_1223),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1230),
.A2(n_1304),
.B(n_1263),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1278),
.Y(n_1337)
);

OR2x6_ASAP7_75t_L g1338 ( 
.A(n_1259),
.B(n_1269),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1259),
.A2(n_1305),
.B(n_1297),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1313),
.B(n_1304),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1297),
.A2(n_1305),
.B(n_1314),
.C(n_1302),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1267),
.B(n_1243),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1253),
.B(n_1250),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1330),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1301),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1295),
.A2(n_1215),
.B1(n_1242),
.B2(n_1217),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1215),
.A2(n_1217),
.B1(n_1314),
.B2(n_1312),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1267),
.B(n_1301),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1235),
.A2(n_1238),
.B(n_1222),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1240),
.A2(n_1292),
.B1(n_1256),
.B2(n_1224),
.C(n_1331),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1226),
.B(n_1245),
.Y(n_1351)
);

O2A1O1Ixp5_ASAP7_75t_L g1352 ( 
.A1(n_1213),
.A2(n_1303),
.B(n_1292),
.C(n_1220),
.Y(n_1352)
);

O2A1O1Ixp5_ASAP7_75t_L g1353 ( 
.A1(n_1213),
.A2(n_1303),
.B(n_1220),
.C(n_1240),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1232),
.B(n_1315),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1315),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1254),
.B(n_1227),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1257),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1322),
.A2(n_1234),
.B1(n_1233),
.B2(n_1309),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1307),
.A2(n_1233),
.B(n_1262),
.C(n_1300),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1234),
.A2(n_1309),
.B1(n_1249),
.B2(n_1256),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1325),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1230),
.A2(n_1263),
.B(n_1248),
.Y(n_1362)
);

O2A1O1Ixp5_ASAP7_75t_L g1363 ( 
.A1(n_1270),
.A2(n_1262),
.B(n_1273),
.C(n_1283),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1248),
.A2(n_1268),
.B(n_1298),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1236),
.B(n_1264),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1317),
.A2(n_1321),
.B1(n_1326),
.B2(n_1251),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1311),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1289),
.A2(n_1285),
.B(n_1296),
.Y(n_1368)
);

O2A1O1Ixp5_ASAP7_75t_L g1369 ( 
.A1(n_1273),
.A2(n_1252),
.B(n_1265),
.C(n_1276),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1279),
.A2(n_1261),
.B1(n_1247),
.B2(n_1281),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1255),
.B(n_1271),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1289),
.B(n_1286),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1287),
.B(n_1290),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1219),
.A2(n_1318),
.B(n_1319),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1274),
.A2(n_1228),
.B(n_1328),
.C(n_1323),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1277),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1274),
.A2(n_1284),
.B(n_1241),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1290),
.B(n_1299),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1299),
.B(n_1237),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1310),
.A2(n_1229),
.B(n_1231),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1306),
.A2(n_1293),
.B(n_1218),
.Y(n_1381)
);

O2A1O1Ixp5_ASAP7_75t_L g1382 ( 
.A1(n_1266),
.A2(n_1329),
.B(n_1327),
.C(n_1282),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1275),
.B(n_1258),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1239),
.B(n_1272),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1291),
.A2(n_1280),
.B(n_1244),
.C(n_1246),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1239),
.B(n_1260),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1239),
.B(n_1316),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1260),
.B(n_1316),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1324),
.A2(n_1216),
.B(n_1272),
.C(n_1260),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1320),
.B(n_1308),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1308),
.B(n_1261),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1235),
.A2(n_1238),
.B(n_1222),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1235),
.A2(n_1238),
.B(n_1222),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1259),
.A2(n_768),
.B(n_1174),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1301),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1295),
.A2(n_768),
.B1(n_1302),
.B2(n_1215),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1295),
.A2(n_768),
.B1(n_1302),
.B2(n_1215),
.Y(n_1397)
);

O2A1O1Ixp5_ASAP7_75t_L g1398 ( 
.A1(n_1259),
.A2(n_1213),
.B(n_1303),
.C(n_1292),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1221),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1259),
.A2(n_768),
.B(n_1174),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1288),
.B(n_1223),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1259),
.A2(n_1213),
.B(n_1303),
.C(n_1292),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1253),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1221),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1221),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1225),
.B(n_1250),
.Y(n_1406)
);

OA22x2_ASAP7_75t_L g1407 ( 
.A1(n_1295),
.A2(n_1302),
.B1(n_1123),
.B2(n_1217),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1221),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1259),
.A2(n_768),
.B(n_1174),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1221),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1214),
.B(n_1294),
.Y(n_1411)
);

O2A1O1Ixp5_ASAP7_75t_L g1412 ( 
.A1(n_1259),
.A2(n_1213),
.B(n_1303),
.C(n_1292),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1373),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1407),
.B(n_1396),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1373),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1372),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1380),
.A2(n_1363),
.B(n_1381),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1332),
.B(n_1335),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1345),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1401),
.B(n_1378),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1340),
.B(n_1401),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1368),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1339),
.A2(n_1379),
.B(n_1341),
.Y(n_1423)
);

CKINVDCx8_ASAP7_75t_R g1424 ( 
.A(n_1338),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1379),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1407),
.B(n_1397),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1338),
.B(n_1372),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1382),
.A2(n_1353),
.B(n_1352),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1390),
.B(n_1338),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1334),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1360),
.B(n_1355),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1383),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1395),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1376),
.B(n_1351),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1346),
.A2(n_1347),
.B(n_1341),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1399),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1398),
.A2(n_1412),
.B(n_1402),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1374),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1368),
.B(n_1351),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1404),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1368),
.B(n_1390),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1350),
.B(n_1394),
.C(n_1409),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1362),
.A2(n_1364),
.B(n_1336),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1374),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1405),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1408),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1410),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1385),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1406),
.B(n_1392),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1371),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1400),
.A2(n_1358),
.B1(n_1342),
.B2(n_1348),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1354),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1359),
.A2(n_1366),
.B1(n_1370),
.B2(n_1375),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1391),
.A2(n_1403),
.B1(n_1361),
.B2(n_1365),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1349),
.Y(n_1455)
);

AO21x2_ASAP7_75t_L g1456 ( 
.A1(n_1385),
.A2(n_1411),
.B(n_1333),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1369),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1445),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1445),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1414),
.A2(n_1344),
.B1(n_1367),
.B2(n_1361),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1430),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1439),
.B(n_1393),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1416),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1430),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1430),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1420),
.B(n_1343),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1436),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1456),
.B(n_1356),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1436),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1429),
.B(n_1383),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1424),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1414),
.A2(n_1391),
.B1(n_1344),
.B2(n_1357),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1422),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1416),
.B(n_1441),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1456),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1416),
.B(n_1441),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1441),
.B(n_1383),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1426),
.B(n_1387),
.Y(n_1479)
);

NAND2x1_ASAP7_75t_L g1480 ( 
.A(n_1432),
.B(n_1377),
.Y(n_1480)
);

OR2x6_ASAP7_75t_SL g1481 ( 
.A(n_1451),
.B(n_1367),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1426),
.B(n_1337),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1476),
.A2(n_1435),
.B1(n_1451),
.B2(n_1457),
.C(n_1431),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1461),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1475),
.B(n_1450),
.Y(n_1485)
);

NOR4xp25_ASAP7_75t_SL g1486 ( 
.A(n_1463),
.B(n_1481),
.C(n_1457),
.D(n_1458),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1479),
.A2(n_1442),
.B1(n_1423),
.B2(n_1453),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1461),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1464),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1475),
.B(n_1450),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1465),
.Y(n_1491)
);

OAI31xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1475),
.A2(n_1442),
.A3(n_1453),
.B(n_1448),
.Y(n_1492)
);

NAND2xp33_ASAP7_75t_SL g1493 ( 
.A(n_1463),
.B(n_1431),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1465),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1481),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_R g1496 ( 
.A(n_1463),
.B(n_1437),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1482),
.A2(n_1442),
.B1(n_1423),
.B2(n_1454),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1466),
.B(n_1421),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1460),
.B(n_1337),
.Y(n_1500)
);

AND2x2_ASAP7_75t_SL g1501 ( 
.A(n_1477),
.B(n_1432),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1476),
.B(n_1457),
.C(n_1448),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_R g1503 ( 
.A(n_1482),
.B(n_1388),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1480),
.A2(n_1422),
.B(n_1455),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1473),
.A2(n_1454),
.B1(n_1448),
.B2(n_1425),
.C(n_1452),
.Y(n_1505)
);

OAI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1473),
.A2(n_1454),
.B1(n_1425),
.B2(n_1452),
.C(n_1415),
.Y(n_1506)
);

AOI33xp33_ASAP7_75t_L g1507 ( 
.A1(n_1462),
.A2(n_1415),
.A3(n_1413),
.B1(n_1440),
.B2(n_1446),
.B3(n_1447),
.Y(n_1507)
);

OR2x6_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1377),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1458),
.Y(n_1509)
);

AOI31xp33_ASAP7_75t_L g1510 ( 
.A1(n_1481),
.A2(n_1433),
.A3(n_1419),
.B(n_1434),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1478),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1460),
.Y(n_1512)
);

OAI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1462),
.A2(n_1418),
.B(n_1415),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1427),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1432),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1479),
.A2(n_1443),
.B(n_1437),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1459),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1472),
.A2(n_1424),
.B1(n_1434),
.B2(n_1437),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1472),
.A2(n_1424),
.B1(n_1437),
.B2(n_1428),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1507),
.B(n_1459),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1497),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1509),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1492),
.A2(n_1423),
.B(n_1437),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_SL g1525 ( 
.A(n_1487),
.B(n_1483),
.C(n_1486),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1519),
.A2(n_1423),
.B(n_1437),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1495),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1507),
.B(n_1462),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1493),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1517),
.B(n_1467),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1504),
.A2(n_1502),
.B(n_1516),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1501),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1484),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1510),
.A2(n_1423),
.B(n_1417),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1477),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1495),
.B(n_1474),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1501),
.B(n_1493),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1488),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1513),
.A2(n_1438),
.B(n_1444),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1505),
.A2(n_1443),
.B(n_1428),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1489),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1491),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1515),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1533),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1532),
.B(n_1512),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1524),
.A2(n_1522),
.B(n_1525),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1533),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1532),
.B(n_1512),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1522),
.B(n_1467),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1538),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1529),
.B(n_1532),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1469),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1532),
.B(n_1514),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1532),
.B(n_1514),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1539),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1528),
.B(n_1419),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1521),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1539),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1433),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1532),
.B(n_1511),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1538),
.Y(n_1565)
);

A2O1A1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1526),
.A2(n_1506),
.B(n_1500),
.C(n_1518),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1511),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1538),
.Y(n_1568)
);

AND2x4_ASAP7_75t_SL g1569 ( 
.A(n_1544),
.B(n_1515),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1527),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1541),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1529),
.B(n_1471),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1472),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1466),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1485),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1539),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1541),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1485),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1530),
.B(n_1466),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1537),
.B(n_1503),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1523),
.B(n_1469),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1526),
.A2(n_1496),
.B1(n_1508),
.B2(n_1468),
.C(n_1428),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1543),
.B(n_1490),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1539),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1577),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1570),
.B(n_1523),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1561),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1546),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1569),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1570),
.B(n_1527),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1527),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1548),
.B(n_1525),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1549),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1546),
.B(n_1537),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1551),
.B(n_1540),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1552),
.B(n_1535),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1547),
.B(n_1536),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1577),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1553),
.B(n_1540),
.Y(n_1603)
);

NAND2x1_ASAP7_75t_SL g1604 ( 
.A(n_1552),
.B(n_1555),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1547),
.B(n_1534),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1549),
.B(n_1542),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1555),
.B(n_1535),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1553),
.B(n_1535),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1565),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1565),
.Y(n_1610)
);

NOR2x1_ASAP7_75t_L g1611 ( 
.A(n_1581),
.B(n_1536),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1568),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1545),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1575),
.B(n_1542),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1568),
.Y(n_1615)
);

OAI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1566),
.A2(n_1583),
.B(n_1556),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1555),
.B(n_1544),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1577),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1583),
.A2(n_1531),
.B1(n_1539),
.B2(n_1544),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1571),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1575),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1580),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1600),
.B(n_1576),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1601),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1576),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1605),
.A2(n_1531),
.B(n_1577),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1591),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1605),
.B(n_1567),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1597),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1599),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1604),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1591),
.B(n_1579),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1586),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1586),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1591),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1590),
.B(n_1569),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1584),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1604),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1584),
.Y(n_1641)
);

INVxp67_ASAP7_75t_SL g1642 ( 
.A(n_1593),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1590),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1592),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1645)
);

AOI31xp33_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_1593),
.A3(n_1611),
.B(n_1595),
.Y(n_1646)
);

NAND2x1_ASAP7_75t_L g1647 ( 
.A(n_1637),
.B(n_1595),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1642),
.A2(n_1619),
.B1(n_1598),
.B2(n_1585),
.Y(n_1648)
);

OAI21xp33_ASAP7_75t_L g1649 ( 
.A1(n_1639),
.A2(n_1613),
.B(n_1617),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1621),
.B(n_1587),
.Y(n_1650)
);

NAND3xp33_ASAP7_75t_SL g1651 ( 
.A(n_1640),
.B(n_1617),
.C(n_1574),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1623),
.B(n_1607),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1626),
.A2(n_1585),
.B1(n_1562),
.B2(n_1559),
.C(n_1531),
.Y(n_1653)
);

NAND4xp25_ASAP7_75t_L g1654 ( 
.A(n_1640),
.B(n_1588),
.C(n_1596),
.D(n_1615),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1637),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1636),
.B(n_1606),
.Y(n_1656)
);

CKINVDCx16_ASAP7_75t_R g1657 ( 
.A(n_1643),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

AOI21xp33_ASAP7_75t_L g1659 ( 
.A1(n_1631),
.A2(n_1606),
.B(n_1609),
.Y(n_1659)
);

OAI322xp33_ASAP7_75t_L g1660 ( 
.A1(n_1624),
.A2(n_1550),
.A3(n_1545),
.B1(n_1620),
.B2(n_1612),
.C1(n_1610),
.C2(n_1563),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1624),
.A2(n_1574),
.B1(n_1608),
.B2(n_1531),
.Y(n_1661)
);

AOI21xp33_ASAP7_75t_L g1662 ( 
.A1(n_1645),
.A2(n_1618),
.B(n_1602),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1621),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1632),
.A2(n_1567),
.B(n_1572),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1657),
.B(n_1644),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1652),
.B(n_1637),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_L g1667 ( 
.A(n_1655),
.B(n_1650),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1622),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1663),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1637),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_R g1671 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1664),
.B(n_1623),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1646),
.B(n_1624),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1660),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1659),
.B1(n_1660),
.B2(n_1654),
.C(n_1648),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1673),
.A2(n_1662),
.B(n_1651),
.C(n_1661),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1673),
.A2(n_1653),
.B1(n_1671),
.B2(n_1674),
.C(n_1665),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1679)
);

NAND4xp25_ASAP7_75t_L g1680 ( 
.A(n_1670),
.B(n_1628),
.C(n_1633),
.D(n_1635),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1668),
.B(n_1638),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1667),
.B(n_1635),
.C(n_1633),
.Y(n_1682)
);

AOI211xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1669),
.A2(n_1638),
.B(n_1630),
.C(n_1629),
.Y(n_1683)
);

NAND4xp75_ASAP7_75t_L g1684 ( 
.A(n_1672),
.B(n_1635),
.C(n_1633),
.D(n_1625),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1671),
.Y(n_1685)
);

A2O1A1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1675),
.A2(n_1585),
.B(n_1562),
.C(n_1559),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1676),
.A2(n_1562),
.B1(n_1559),
.B2(n_1618),
.C(n_1602),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1679),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1682),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1678),
.A2(n_1531),
.B1(n_1630),
.B2(n_1634),
.Y(n_1690)
);

NOR2x1_ASAP7_75t_L g1691 ( 
.A(n_1680),
.B(n_1684),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1641),
.Y(n_1692)
);

INVxp33_ASAP7_75t_SL g1693 ( 
.A(n_1691),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1692),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1689),
.B(n_1681),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1688),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1687),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1690),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1695),
.A2(n_1693),
.B(n_1677),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1694),
.B(n_1614),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1698),
.A2(n_1683),
.B(n_1686),
.Y(n_1701)
);

BUFx8_ASAP7_75t_SL g1702 ( 
.A(n_1697),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1697),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1696),
.B1(n_1550),
.B2(n_1572),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1702),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1701),
.A2(n_1531),
.B1(n_1557),
.B2(n_1558),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1705),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1706),
.B1(n_1699),
.B2(n_1704),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1700),
.B1(n_1558),
.B2(n_1557),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1708),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1709),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1710),
.A2(n_1573),
.B(n_1571),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1711),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1712),
.A2(n_1560),
.B1(n_1563),
.B2(n_1578),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1713),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1715),
.B(n_1714),
.Y(n_1716)
);

NOR2xp67_ASAP7_75t_L g1717 ( 
.A(n_1716),
.B(n_1573),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1717),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1718),
.A2(n_1578),
.B1(n_1582),
.B2(n_1574),
.C(n_1564),
.Y(n_1719)
);

AOI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1386),
.B(n_1389),
.C(n_1384),
.Y(n_1720)
);


endmodule