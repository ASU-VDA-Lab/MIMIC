module fake_jpeg_11215_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_2),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_51),
.Y(n_149)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_52),
.Y(n_114)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_75),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_14),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_40),
.B1(n_39),
.B2(n_46),
.Y(n_98)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_23),
.B(n_14),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_84),
.B(n_85),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_92),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_96),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_13),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_98),
.A2(n_29),
.B1(n_16),
.B2(n_38),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_101),
.B(n_117),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_27),
.B1(n_39),
.B2(n_26),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_103),
.A2(n_104),
.B1(n_33),
.B2(n_16),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_32),
.B1(n_22),
.B2(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_33),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_82),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_49),
.A2(n_28),
.B1(n_36),
.B2(n_42),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_65),
.B1(n_72),
.B2(n_71),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_135),
.B(n_143),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_48),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_38),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_36),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_157),
.Y(n_219)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_111),
.B(n_150),
.C(n_152),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_160),
.A2(n_34),
.B(n_13),
.C(n_145),
.Y(n_243)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_165),
.Y(n_224)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_103),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_179),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_120),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_29),
.B1(n_148),
.B2(n_108),
.Y(n_210)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_182),
.Y(n_217)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_112),
.A2(n_28),
.B1(n_36),
.B2(n_48),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_203),
.B(n_134),
.Y(n_205)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_185),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_187),
.Y(n_233)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_190),
.Y(n_235)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_192),
.Y(n_204)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_197),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_238)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_131),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_124),
.A2(n_48),
.B1(n_105),
.B2(n_116),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_205),
.A2(n_239),
.B(n_168),
.C(n_166),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_210),
.A2(n_218),
.B1(n_237),
.B2(n_179),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_131),
.B1(n_149),
.B2(n_110),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_146),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_230),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_155),
.B(n_111),
.C(n_124),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_137),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_155),
.B(n_139),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_155),
.A2(n_149),
.B1(n_115),
.B2(n_108),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_122),
.B1(n_116),
.B2(n_181),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_160),
.A2(n_114),
.B(n_31),
.C(n_30),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_148),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_154),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_247),
.B(n_249),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_164),
.B(n_203),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_255),
.B(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_267),
.B1(n_216),
.B2(n_217),
.Y(n_304)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_256),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_161),
.B(n_177),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_270),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_212),
.A2(n_180),
.B1(n_122),
.B2(n_95),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_258),
.A2(n_266),
.B1(n_237),
.B2(n_218),
.Y(n_286)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_212),
.A2(n_180),
.B1(n_94),
.B2(n_88),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_279),
.B1(n_252),
.B2(n_222),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_261),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_228),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_275),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_205),
.A2(n_193),
.B(n_173),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_83),
.B1(n_86),
.B2(n_70),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_176),
.B(n_184),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_221),
.B(n_233),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_220),
.B(n_185),
.Y(n_270)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_271),
.A2(n_273),
.B1(n_276),
.B2(n_222),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_208),
.B(n_158),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_274),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_225),
.A2(n_192),
.B1(n_187),
.B2(n_159),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_208),
.B(n_178),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_215),
.B(n_59),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_48),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_225),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_232),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_241),
.A2(n_56),
.B1(n_68),
.B2(n_67),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_282),
.B1(n_295),
.B2(n_296),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_238),
.B1(n_204),
.B2(n_243),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_231),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_292),
.C(n_267),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_307),
.B1(n_279),
.B2(n_278),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_18),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_231),
.C(n_211),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_223),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_293),
.B(n_309),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_219),
.B1(n_215),
.B2(n_209),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_248),
.A2(n_219),
.B1(n_209),
.B2(n_232),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_236),
.B(n_229),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_301),
.A2(n_240),
.B(n_271),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_308),
.B1(n_312),
.B2(n_197),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_258),
.A2(n_211),
.B1(n_229),
.B2(n_236),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_244),
.B(n_249),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_267),
.A2(n_226),
.B(n_222),
.C(n_242),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_269),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_263),
.A2(n_226),
.B1(n_51),
.B2(n_64),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_316),
.A2(n_319),
.B1(n_325),
.B2(n_312),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_299),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_323),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_286),
.A2(n_255),
.B1(n_267),
.B2(n_253),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_320),
.A2(n_327),
.B(n_291),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_295),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_266),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_256),
.B1(n_251),
.B2(n_276),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_257),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_305),
.A2(n_246),
.B1(n_213),
.B2(n_242),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_328),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_240),
.B1(n_271),
.B2(n_197),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_296),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_18),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_337),
.Y(n_349)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_48),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_336),
.B(n_302),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_303),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_282),
.A2(n_313),
.B1(n_280),
.B2(n_290),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_339),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_310),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_301),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_340),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_280),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_342),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_290),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_1),
.Y(n_343)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_368),
.B1(n_329),
.B2(n_283),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_321),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_342),
.Y(n_372)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_315),
.Y(n_355)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_311),
.B(n_297),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_356),
.A2(n_366),
.B(n_331),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_314),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_315),
.Y(n_361)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_343),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_289),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_335),
.C(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_367),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_300),
.B1(n_294),
.B2(n_292),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_317),
.B(n_291),
.Y(n_370)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_370),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_379),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_366),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_346),
.B(n_339),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_337),
.Y(n_380)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_389),
.Y(n_404)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_324),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_391),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_323),
.B1(n_316),
.B2(n_325),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_353),
.B1(n_348),
.B2(n_349),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_335),
.C(n_318),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_386),
.C(n_387),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_294),
.C(n_328),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_288),
.C(n_306),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_369),
.C(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g391 ( 
.A1(n_351),
.A2(n_327),
.B(n_341),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_392),
.A2(n_393),
.B1(n_355),
.B2(n_361),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_396),
.A2(n_409),
.B1(n_410),
.B2(n_382),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_397),
.B(n_398),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_373),
.B(n_349),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_356),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_387),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_373),
.B(n_348),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_405),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_345),
.Y(n_405)
);

NOR3xp33_ASAP7_75t_SL g408 ( 
.A(n_380),
.B(n_372),
.C(n_346),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_408),
.B(n_378),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_352),
.B1(n_345),
.B2(n_360),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_352),
.B1(n_358),
.B2(n_363),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_406),
.A2(n_389),
.B(n_386),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_412),
.A2(n_425),
.B(n_376),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_423),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_381),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_SL g439 ( 
.A(n_414),
.B(n_421),
.Y(n_439)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_392),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_420),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_371),
.C(n_350),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_377),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_358),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_378),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_424),
.A2(n_347),
.B1(n_285),
.B2(n_6),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_394),
.A2(n_388),
.B(n_375),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_350),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_376),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_418),
.A2(n_400),
.B1(n_395),
.B2(n_401),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_430),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_429),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_405),
.C(n_404),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_397),
.B(n_403),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_434),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_437),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_423),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_367),
.C(n_347),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_435),
.B(n_438),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_413),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_444),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_417),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_417),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_446),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_285),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_432),
.B(n_419),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_6),
.Y(n_458)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_419),
.C(n_426),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_450),
.A2(n_438),
.B(n_5),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_427),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_458),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_439),
.B(n_431),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_454),
.A2(n_455),
.B(n_456),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_12),
.B(n_6),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_1),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_457),
.Y(n_462)
);

INVx6_ASAP7_75t_L g459 ( 
.A(n_451),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_459),
.A2(n_463),
.B(n_7),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_447),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_460),
.A2(n_449),
.B(n_450),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_464),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_461),
.A2(n_7),
.B(n_9),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_465),
.A2(n_466),
.B(n_462),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_467),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_468),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_10),
.Y(n_472)
);


endmodule