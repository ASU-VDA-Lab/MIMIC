module fake_ibex_1953_n_4028 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_848, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4028);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4028;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_2979;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_2333;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3766;
wire n_2822;
wire n_3022;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3667;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3719;
wire n_3390;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_3070;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_3398;
wire n_3718;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3682;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3434;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3746;
wire n_2758;
wire n_3480;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_3506;
wire n_2845;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3349;
wire n_3928;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_1622;
wire n_897;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_1542;
wire n_1586;
wire n_1362;
wire n_946;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3919;
wire n_3683;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_2928;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_3557;
wire n_3596;
wire n_3207;
wire n_3067;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_3873;
wire n_2917;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_205),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_843),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_20),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_384),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_568),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_131),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_573),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_552),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_202),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_370),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_366),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_841),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_377),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_65),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_842),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_826),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_845),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_755),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_775),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_148),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_526),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_42),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_548),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_281),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_645),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_235),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_390),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_47),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_32),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_515),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_282),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_266),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_644),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_422),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_827),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_205),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_406),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_369),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_181),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_614),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_587),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_271),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_689),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_342),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_313),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_745),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_524),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_682),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_776),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_652),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_136),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_407),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_373),
.Y(n_901)
);

INVxp33_ASAP7_75t_SL g902 ( 
.A(n_220),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_293),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_788),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_400),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_396),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_76),
.Y(n_907)
);

CKINVDCx14_ASAP7_75t_R g908 ( 
.A(n_50),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_58),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_116),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_197),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_590),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_805),
.Y(n_913)
);

BUFx5_ASAP7_75t_L g914 ( 
.A(n_819),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_362),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_43),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_247),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_57),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_563),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_352),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_756),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_34),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_193),
.Y(n_923)
);

CKINVDCx14_ASAP7_75t_R g924 ( 
.A(n_749),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_174),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_492),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_830),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_63),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_411),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_672),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_30),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_130),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_405),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_445),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_406),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_49),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_714),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_523),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_445),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_117),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_34),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_174),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_44),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_712),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_466),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_292),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_255),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_708),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_653),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_186),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_799),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_624),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_786),
.Y(n_953)
);

CKINVDCx14_ASAP7_75t_R g954 ( 
.A(n_834),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_252),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_292),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_630),
.Y(n_957)
);

INVx4_ASAP7_75t_R g958 ( 
.A(n_368),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_835),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_376),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_150),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_838),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_635),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_77),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_132),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_837),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_198),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_338),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_92),
.Y(n_969)
);

BUFx8_ASAP7_75t_SL g970 ( 
.A(n_544),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_294),
.Y(n_971)
);

CKINVDCx14_ASAP7_75t_R g972 ( 
.A(n_320),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_313),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_521),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_468),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_197),
.Y(n_976)
);

CKINVDCx16_ASAP7_75t_R g977 ( 
.A(n_284),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_477),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_629),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_597),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_332),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_217),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_607),
.Y(n_983)
);

CKINVDCx14_ASAP7_75t_R g984 ( 
.A(n_743),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_137),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_575),
.Y(n_986)
);

BUFx5_ASAP7_75t_L g987 ( 
.A(n_160),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_341),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_162),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_756),
.Y(n_990)
);

CKINVDCx14_ASAP7_75t_R g991 ( 
.A(n_46),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_547),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_752),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_216),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_392),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_369),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_249),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_74),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_575),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_709),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_754),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_267),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_720),
.Y(n_1003)
);

BUFx5_ASAP7_75t_L g1004 ( 
.A(n_97),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_405),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_599),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_376),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_13),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_247),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_137),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_632),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_823),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_471),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_599),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_784),
.Y(n_1015)
);

BUFx8_ASAP7_75t_SL g1016 ( 
.A(n_231),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_161),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_845),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_800),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_158),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_169),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_137),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_95),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_745),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_453),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_799),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_124),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_763),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_538),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_307),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_37),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_709),
.Y(n_1032)
);

INVxp33_ASAP7_75t_L g1033 ( 
.A(n_444),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_715),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_337),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_329),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_217),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_167),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_683),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_238),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_698),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_253),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_567),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_309),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_737),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_674),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_823),
.Y(n_1047)
);

BUFx2_ASAP7_75t_R g1048 ( 
.A(n_211),
.Y(n_1048)
);

BUFx8_ASAP7_75t_SL g1049 ( 
.A(n_822),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_697),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_587),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_116),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_209),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_276),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_75),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_747),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_404),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_267),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_322),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_510),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_638),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_320),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_833),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_253),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_690),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_81),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_433),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_515),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_614),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_106),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_181),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_291),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_151),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_590),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_228),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_501),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_836),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_847),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_613),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_510),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_6),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_508),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_152),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_428),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_307),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_473),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_319),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_367),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_759),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_60),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_645),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_30),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_480),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_329),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_383),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_66),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_505),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_753),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_780),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_817),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_200),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_763),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_724),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_603),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_341),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_318),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_150),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_767),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_120),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_431),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_0),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_473),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_566),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_97),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_319),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_115),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_621),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_3),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_12),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_240),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_173),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_123),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_658),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_32),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_556),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_312),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_68),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_593),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_819),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_97),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_7),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_43),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_827),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_413),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_232),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_108),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_673),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_11),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_509),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_425),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_806),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_39),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_758),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_433),
.Y(n_1144)
);

BUFx5_ASAP7_75t_L g1145 ( 
.A(n_615),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_509),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_558),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_39),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_486),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_659),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_0),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_121),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_623),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_701),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_832),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_791),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_800),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_480),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_514),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_588),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_400),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_227),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_825),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_228),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_836),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_277),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_583),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_804),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_42),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_92),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_555),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_828),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_262),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_808),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_550),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_235),
.Y(n_1176)
);

CKINVDCx14_ASAP7_75t_R g1177 ( 
.A(n_491),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_219),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_375),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_296),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_569),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_518),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_166),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_766),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_431),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_676),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_628),
.Y(n_1187)
);

CKINVDCx12_ASAP7_75t_R g1188 ( 
.A(n_797),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_829),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_767),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_8),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_55),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_88),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_3),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_128),
.Y(n_1195)
);

BUFx5_ASAP7_75t_L g1196 ( 
.A(n_327),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_224),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_552),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_89),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_297),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_618),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_189),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_788),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_747),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_455),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_194),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_28),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_525),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_345),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_2),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_499),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_154),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_44),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_41),
.Y(n_1214)
);

CKINVDCx16_ASAP7_75t_R g1215 ( 
.A(n_163),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_150),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_629),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_182),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_180),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_462),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_208),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_94),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_557),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_360),
.Y(n_1224)
);

BUFx10_ASAP7_75t_L g1225 ( 
.A(n_276),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_840),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_472),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_469),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_573),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_12),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_166),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_534),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_336),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_95),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_286),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_124),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_681),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_752),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_57),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_560),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_328),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_260),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_605),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_372),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_192),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_308),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_844),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_757),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_595),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_69),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_499),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_85),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_392),
.Y(n_1253)
);

BUFx10_ASAP7_75t_L g1254 ( 
.A(n_514),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_145),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_824),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_467),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_343),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_340),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_843),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_622),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_839),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_182),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_666),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_92),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_701),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_42),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_790),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_438),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_551),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_401),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_361),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_177),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_172),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_32),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_842),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_831),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_380),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_839),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_908),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_991),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_876),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_862),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_965),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_970),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_965),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_L g1287 ( 
.A(n_965),
.B(n_0),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_868),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_985),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_914),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1053),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1033),
.B(n_1),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1048),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_R g1294 ( 
.A(n_924),
.B(n_1),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_989),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1092),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_926),
.B(n_1),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1092),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_899),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1109),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1002),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1109),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_970),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_914),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_857),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1016),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1111),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_876),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1111),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1016),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1102),
.B(n_2),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1049),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_950),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_880),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_950),
.Y(n_1315)
);

CKINVDCx16_ASAP7_75t_R g1316 ( 
.A(n_910),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_880),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_944),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1216),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_916),
.B(n_2),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_893),
.B(n_3),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1049),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_857),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_944),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1058),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1058),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_899),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_935),
.B(n_4),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1105),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1216),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1252),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_954),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1252),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1105),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1071),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_972),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1147),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1078),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1215),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_984),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1147),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1144),
.B(n_4),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1197),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1177),
.B(n_4),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_1204),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1204),
.Y(n_1346)
);

CKINVDCx16_ASAP7_75t_R g1347 ( 
.A(n_1081),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1272),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_907),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_849),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_977),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_854),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1261),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_870),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_877),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_884),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_887),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_918),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_872),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_923),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1037),
.B(n_5),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_872),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_874),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_874),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_875),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_931),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_875),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_932),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_913),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_909),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_936),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1096),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_987),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_911),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_913),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_925),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_928),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_940),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_941),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_967),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_929),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_942),
.Y(n_1382)
);

CKINVDCx16_ASAP7_75t_R g1383 ( 
.A(n_1225),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_943),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1096),
.Y(n_1385)
);

CKINVDCx16_ASAP7_75t_R g1386 ( 
.A(n_1225),
.Y(n_1386)
);

INVxp33_ASAP7_75t_SL g1387 ( 
.A(n_961),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_964),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_969),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1275),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_976),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_914),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1010),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1335),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1304),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1392),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1373),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1345),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1373),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1284),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1287),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1296),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1286),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1293),
.A2(n_1308),
.B1(n_1313),
.B2(n_1282),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1327),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1387),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1298),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1288),
.B(n_1289),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1385),
.B(n_994),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1300),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1302),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1307),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1295),
.B(n_898),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1309),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1314),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1305),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1390),
.B(n_998),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1317),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1339),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1349),
.A2(n_1022),
.B(n_851),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1350),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1323),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1372),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1345),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1318),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1393),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1324),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1325),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1326),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1329),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1291),
.A2(n_1008),
.B1(n_1027),
.B2(n_1020),
.Y(n_1431)
);

AND2x6_ASAP7_75t_L g1432 ( 
.A(n_1297),
.B(n_1275),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1283),
.B(n_987),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1338),
.B(n_1142),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1334),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1337),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1281),
.B(n_987),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1348),
.B(n_987),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1352),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1299),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1341),
.B(n_898),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1343),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1358),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1346),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1360),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1376),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1366),
.Y(n_1447)
);

NAND2xp33_ASAP7_75t_L g1448 ( 
.A(n_1280),
.B(n_987),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1377),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1368),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1371),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1301),
.B(n_902),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1380),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1389),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1354),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1342),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1321),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1328),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1315),
.A2(n_966),
.B1(n_975),
.B2(n_968),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1355),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1361),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1356),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1361),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1292),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1357),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1320),
.B(n_973),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1370),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1311),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1311),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1292),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1374),
.B(n_1077),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1378),
.A2(n_1022),
.B(n_851),
.Y(n_1472)
);

CKINVDCx8_ASAP7_75t_R g1473 ( 
.A(n_1316),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1379),
.B(n_1038),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1294),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1344),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1382),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1384),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1388),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1391),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1383),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1386),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1332),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1336),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1340),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1285),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1303),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1306),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1310),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1312),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1351),
.B(n_1066),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1322),
.A2(n_1148),
.B(n_1021),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1353),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1319),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1330),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1331),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1333),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1359),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1362),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_L g1500 ( 
.A(n_1363),
.B(n_1083),
.C(n_1073),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1364),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1365),
.B(n_1004),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1367),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1369),
.B(n_1090),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1375),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1381),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1286),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1286),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1286),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1299),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1286),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1291),
.A2(n_1114),
.B1(n_1116),
.B2(n_1101),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1286),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1286),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1299),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_SL g1516 ( 
.A(n_1347),
.B(n_1118),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1286),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1286),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1327),
.Y(n_1519)
);

BUFx8_ASAP7_75t_L g1520 ( 
.A(n_1283),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1286),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1283),
.B(n_1004),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1335),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1345),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1345),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1286),
.Y(n_1526)
);

INVx5_ASAP7_75t_L g1527 ( 
.A(n_1345),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1335),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1335),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1345),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1290),
.Y(n_1531)
);

AND2x4_ASAP7_75t_SL g1532 ( 
.A(n_1281),
.B(n_1225),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1327),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1335),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1281),
.B(n_902),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1345),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1283),
.B(n_1004),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1335),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1335),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1283),
.B(n_1004),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1345),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1288),
.B(n_1077),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1347),
.B(n_1004),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1345),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1373),
.A2(n_1148),
.B(n_1023),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1286),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1345),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1385),
.B(n_1121),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1290),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1290),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1288),
.B(n_1095),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1373),
.A2(n_1031),
.B(n_1017),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1286),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1299),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1286),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1281),
.B(n_1124),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1290),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1345),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1425),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1527),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1452),
.A2(n_1274),
.B1(n_1273),
.B2(n_1130),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1420),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1421),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1523),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1398),
.B(n_1127),
.Y(n_1567)
);

AO22x2_ASAP7_75t_L g1568 ( 
.A1(n_1459),
.A2(n_968),
.B1(n_975),
.B2(n_966),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1427),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1427),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1429),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_974),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1456),
.B(n_1131),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1398),
.B(n_1132),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1429),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1402),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1407),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_L g1578 ( 
.A(n_1432),
.B(n_914),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1419),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1414),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1434),
.B(n_1254),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1439),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1462),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1406),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1552),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1410),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1410),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1446),
.Y(n_1588)
);

CKINVDCx16_ASAP7_75t_R g1589 ( 
.A(n_1516),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1424),
.B(n_1152),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1558),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1449),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1411),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1440),
.B(n_1254),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1464),
.B(n_1170),
.Y(n_1595)
);

AND2x4_ASAP7_75t_SL g1596 ( 
.A(n_1482),
.B(n_1254),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1533),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1411),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1524),
.B(n_1095),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1520),
.Y(n_1600)
);

AND2x2_ASAP7_75t_SL g1601 ( 
.A(n_1532),
.B(n_1070),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1415),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1529),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1464),
.B(n_1183),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1520),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1529),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1418),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1524),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1428),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1525),
.B(n_1097),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1525),
.B(n_1191),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1510),
.B(n_895),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1504),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1552),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1530),
.B(n_1536),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1470),
.B(n_1267),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1442),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1451),
.B(n_1403),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1403),
.B(n_1192),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1470),
.B(n_1193),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1412),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1515),
.B(n_895),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1409),
.B(n_1195),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1482),
.B(n_889),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1545),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1408),
.A2(n_1206),
.B1(n_1210),
.B2(n_1202),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1417),
.B(n_1212),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1473),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1558),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1470),
.B(n_1213),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1545),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1430),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1435),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1538),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1468),
.A2(n_1119),
.B1(n_1136),
.B2(n_1107),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1538),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1394),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1472),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1457),
.B(n_1218),
.Y(n_1639)
);

OR2x6_ASAP7_75t_L g1640 ( 
.A(n_1493),
.B(n_986),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1436),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_L g1642 ( 
.A(n_1432),
.B(n_914),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1472),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1548),
.B(n_1221),
.Y(n_1644)
);

NOR3xp33_ASAP7_75t_L g1645 ( 
.A(n_1404),
.B(n_885),
.C(n_852),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1444),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1441),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1441),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1400),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1400),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1493),
.B(n_986),
.Y(n_1651)
);

BUFx10_ASAP7_75t_L g1652 ( 
.A(n_1481),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1457),
.B(n_1222),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1426),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1426),
.Y(n_1655)
);

AND2x2_ASAP7_75t_SL g1656 ( 
.A(n_1455),
.B(n_1151),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1541),
.B(n_1097),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1544),
.B(n_1239),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1544),
.B(n_1123),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1495),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1443),
.Y(n_1661)
);

BUFx10_ASAP7_75t_L g1662 ( 
.A(n_1481),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1528),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1466),
.B(n_1546),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1554),
.B(n_900),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1443),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1547),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1475),
.B(n_1250),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_SL g1669 ( 
.A(n_1493),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1489),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1431),
.B(n_900),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1450),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1512),
.B(n_889),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1507),
.B(n_1255),
.Y(n_1674)
);

BUFx8_ASAP7_75t_SL g1675 ( 
.A(n_1499),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1508),
.B(n_1169),
.Y(n_1676)
);

AND2x6_ASAP7_75t_L g1677 ( 
.A(n_1458),
.B(n_922),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1453),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1494),
.B(n_1003),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1489),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1509),
.B(n_1194),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1461),
.B(n_850),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1511),
.B(n_1199),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1433),
.B(n_1279),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1513),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1494),
.B(n_1003),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1463),
.B(n_853),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1514),
.B(n_1207),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1556),
.B(n_892),
.C(n_890),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1460),
.B(n_1123),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1517),
.B(n_1214),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1460),
.Y(n_1692)
);

INVx8_ASAP7_75t_L g1693 ( 
.A(n_1490),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1534),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1477),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1518),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1522),
.B(n_896),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1465),
.B(n_1228),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1471),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1471),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1521),
.B(n_1219),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1539),
.Y(n_1702)
);

INVxp33_ASAP7_75t_SL g1703 ( 
.A(n_1479),
.Y(n_1703)
);

AND2x6_ASAP7_75t_L g1704 ( 
.A(n_1465),
.B(n_922),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1469),
.A2(n_1231),
.B1(n_1234),
.B2(n_1230),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1526),
.B(n_1236),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1467),
.B(n_1228),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1490),
.Y(n_1708)
);

BUFx4f_ASAP7_75t_L g1709 ( 
.A(n_1490),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1553),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1555),
.Y(n_1711)
);

CKINVDCx20_ASAP7_75t_R g1712 ( 
.A(n_1405),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1537),
.B(n_1279),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1416),
.B(n_1422),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1423),
.B(n_1438),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1401),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1437),
.B(n_1245),
.Y(n_1717)
);

AO22x2_ASAP7_75t_L g1718 ( 
.A1(n_1496),
.A2(n_1025),
.B1(n_1043),
.B2(n_1012),
.Y(n_1718)
);

NAND3x1_ASAP7_75t_L g1719 ( 
.A(n_1498),
.B(n_1497),
.C(n_1503),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1408),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1540),
.B(n_1263),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1519),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1467),
.B(n_1251),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1413),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1480),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1474),
.B(n_892),
.C(n_890),
.Y(n_1726)
);

CKINVDCx11_ASAP7_75t_R g1727 ( 
.A(n_1494),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1445),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1535),
.B(n_859),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1492),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1432),
.A2(n_1476),
.B1(n_1492),
.B2(n_1502),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1447),
.B(n_1265),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1432),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1413),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1480),
.B(n_1063),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1454),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1491),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1498),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1501),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1478),
.A2(n_1551),
.B1(n_1542),
.B2(n_1483),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1484),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1483),
.B(n_861),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1551),
.Y(n_1743)
);

BUFx10_ASAP7_75t_L g1744 ( 
.A(n_1488),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1506),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1484),
.B(n_894),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1486),
.B(n_1487),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1486),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1395),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1485),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1543),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1505),
.B(n_894),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1396),
.B(n_1052),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1531),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1755)
);

BUFx10_ASAP7_75t_L g1756 ( 
.A(n_1549),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1550),
.Y(n_1757)
);

INVx5_ASAP7_75t_L g1758 ( 
.A(n_1550),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1500),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1557),
.Y(n_1760)
);

AO22x2_ASAP7_75t_L g1761 ( 
.A1(n_1722),
.A2(n_1025),
.B1(n_1043),
.B2(n_1012),
.Y(n_1761)
);

AO22x2_ASAP7_75t_L g1762 ( 
.A1(n_1673),
.A2(n_1046),
.B1(n_1051),
.B2(n_1044),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1664),
.B(n_1448),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1588),
.B(n_1044),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1618),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1586),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1587),
.Y(n_1767)
);

AO22x2_ASAP7_75t_L g1768 ( 
.A1(n_1718),
.A2(n_1051),
.B1(n_1057),
.B2(n_1046),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1593),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1598),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1685),
.B(n_1277),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1584),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1696),
.B(n_1278),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1592),
.B(n_1057),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1710),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1563),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1711),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1778)
);

AO22x2_ASAP7_75t_L g1779 ( 
.A1(n_1718),
.A2(n_1062),
.B1(n_1065),
.B2(n_1061),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1695),
.B(n_1597),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1647),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1648),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1573),
.B(n_1619),
.Y(n_1783)
);

AO22x2_ASAP7_75t_L g1784 ( 
.A1(n_1730),
.A2(n_1062),
.B1(n_1065),
.B2(n_1061),
.Y(n_1784)
);

AO22x2_ASAP7_75t_L g1785 ( 
.A1(n_1600),
.A2(n_1076),
.B1(n_1079),
.B2(n_1067),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1737),
.B(n_1278),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1720),
.A2(n_1188),
.B1(n_865),
.B2(n_866),
.Y(n_1787)
);

AND2x6_ASAP7_75t_L g1788 ( 
.A(n_1733),
.B(n_1052),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1715),
.B(n_863),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1596),
.B(n_1067),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1621),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1656),
.B(n_1076),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1675),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1581),
.B(n_1079),
.Y(n_1794)
);

XOR2x2_ASAP7_75t_L g1795 ( 
.A(n_1703),
.B(n_7),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1626),
.A2(n_934),
.B1(n_937),
.B2(n_901),
.C(n_891),
.Y(n_1796)
);

XNOR2xp5_ASAP7_75t_L g1797 ( 
.A(n_1601),
.B(n_1082),
.Y(n_1797)
);

AO22x2_ASAP7_75t_L g1798 ( 
.A1(n_1730),
.A2(n_1087),
.B1(n_1115),
.B2(n_1082),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1632),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1735),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1633),
.Y(n_1801)
);

AO22x2_ASAP7_75t_L g1802 ( 
.A1(n_1613),
.A2(n_1645),
.B1(n_1568),
.B2(n_1740),
.Y(n_1802)
);

NAND2x1p5_ASAP7_75t_L g1803 ( 
.A(n_1566),
.B(n_990),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1641),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1624),
.Y(n_1805)
);

AO22x2_ASAP7_75t_L g1806 ( 
.A1(n_1568),
.A2(n_1115),
.B1(n_1150),
.B2(n_1087),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1646),
.Y(n_1807)
);

AO22x2_ASAP7_75t_L g1808 ( 
.A1(n_1671),
.A2(n_1153),
.B1(n_1158),
.B2(n_1150),
.Y(n_1808)
);

AO22x2_ASAP7_75t_L g1809 ( 
.A1(n_1759),
.A2(n_1158),
.B1(n_1179),
.B2(n_1153),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1649),
.Y(n_1810)
);

AND2x2_ASAP7_75t_SL g1811 ( 
.A(n_1589),
.B(n_1179),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1650),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1736),
.Y(n_1813)
);

NOR2xp67_ASAP7_75t_L g1814 ( 
.A(n_1605),
.B(n_7),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1612),
.A2(n_1622),
.B1(n_1665),
.B2(n_1594),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1724),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1566),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1652),
.Y(n_1818)
);

AO22x2_ASAP7_75t_L g1819 ( 
.A1(n_1690),
.A2(n_1189),
.B1(n_1262),
.B2(n_1238),
.Y(n_1819)
);

AO22x2_ASAP7_75t_L g1820 ( 
.A1(n_1690),
.A2(n_1189),
.B1(n_1262),
.B2(n_1238),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1734),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1728),
.Y(n_1822)
);

NAND2x1p5_ASAP7_75t_L g1823 ( 
.A(n_1692),
.B(n_1181),
.Y(n_1823)
);

NAND2x1p5_ASAP7_75t_L g1824 ( 
.A(n_1692),
.B(n_1251),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1729),
.A2(n_873),
.B1(n_878),
.B2(n_869),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1591),
.Y(n_1826)
);

AO22x2_ASAP7_75t_L g1827 ( 
.A1(n_1698),
.A2(n_856),
.B1(n_871),
.B2(n_867),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1662),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1576),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1635),
.A2(n_883),
.B1(n_886),
.B2(n_882),
.C(n_879),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1577),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1580),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1602),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1640),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1746),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1607),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1684),
.B(n_903),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1628),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1756),
.B(n_1741),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1609),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1617),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1623),
.B(n_906),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1714),
.Y(n_1843)
);

AO22x2_ASAP7_75t_L g1844 ( 
.A1(n_1698),
.A2(n_897),
.B1(n_904),
.B2(n_881),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1755),
.Y(n_1845)
);

XNOR2xp5_ASAP7_75t_L g1846 ( 
.A(n_1579),
.B(n_8),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1712),
.B(n_905),
.Y(n_1847)
);

AO22x2_ASAP7_75t_L g1848 ( 
.A1(n_1707),
.A2(n_1723),
.B1(n_1651),
.B2(n_1640),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1627),
.B(n_912),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1749),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1749),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1757),
.Y(n_1852)
);

NOR2xp67_ASAP7_75t_L g1853 ( 
.A(n_1726),
.B(n_8),
.Y(n_1853)
);

AND2x6_ASAP7_75t_SL g1854 ( 
.A(n_1651),
.B(n_920),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1697),
.B(n_915),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1699),
.B(n_917),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1682),
.A2(n_1122),
.B1(n_1138),
.B2(n_1055),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1757),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1679),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1679),
.Y(n_1860)
);

OAI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1705),
.A2(n_927),
.B1(n_939),
.B2(n_938),
.C(n_919),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1725),
.B(n_921),
.Y(n_1862)
);

AO22x2_ASAP7_75t_L g1863 ( 
.A1(n_1707),
.A2(n_933),
.B1(n_953),
.B2(n_930),
.Y(n_1863)
);

AO22x2_ASAP7_75t_L g1864 ( 
.A1(n_1723),
.A2(n_962),
.B1(n_963),
.B2(n_960),
.Y(n_1864)
);

OR2x6_ASAP7_75t_L g1865 ( 
.A(n_1686),
.B(n_855),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1693),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1559),
.Y(n_1867)
);

AO22x2_ASAP7_75t_L g1868 ( 
.A1(n_1686),
.A2(n_978),
.B1(n_983),
.B2(n_971),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1731),
.A2(n_1000),
.B1(n_1005),
.B2(n_997),
.Y(n_1869)
);

AO22x2_ASAP7_75t_L g1870 ( 
.A1(n_1745),
.A2(n_1007),
.B1(n_1009),
.B2(n_1006),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1569),
.Y(n_1871)
);

AO22x2_ASAP7_75t_L g1872 ( 
.A1(n_1743),
.A2(n_1013),
.B1(n_1019),
.B2(n_1011),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1570),
.Y(n_1873)
);

AO22x2_ASAP7_75t_L g1874 ( 
.A1(n_1700),
.A2(n_1028),
.B1(n_1032),
.B2(n_1026),
.Y(n_1874)
);

NAND2x1p5_ASAP7_75t_L g1875 ( 
.A(n_1608),
.B(n_1629),
.Y(n_1875)
);

AO22x2_ASAP7_75t_L g1876 ( 
.A1(n_1752),
.A2(n_1035),
.B1(n_1036),
.B2(n_1034),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1571),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1575),
.Y(n_1878)
);

OR2x2_ASAP7_75t_SL g1879 ( 
.A(n_1689),
.B(n_958),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1754),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1760),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1733),
.A2(n_1040),
.B1(n_1041),
.B2(n_1039),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1716),
.Y(n_1883)
);

NAND2x1p5_ASAP7_75t_L g1884 ( 
.A(n_1608),
.B(n_1055),
.Y(n_1884)
);

AND2x6_ASAP7_75t_L g1885 ( 
.A(n_1733),
.B(n_1055),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1676),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1644),
.B(n_945),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1758),
.B(n_946),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1681),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1629),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1567),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1585),
.Y(n_1892)
);

AO22x2_ASAP7_75t_L g1893 ( 
.A1(n_1599),
.A2(n_1050),
.B1(n_1056),
.B2(n_1045),
.Y(n_1893)
);

BUFx8_ASAP7_75t_L g1894 ( 
.A(n_1669),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1747),
.B(n_947),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1683),
.Y(n_1896)
);

OAI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1561),
.A2(n_951),
.B1(n_952),
.B2(n_949),
.C(n_948),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1585),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1688),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1585),
.Y(n_1900)
);

AO22x2_ASAP7_75t_L g1901 ( 
.A1(n_1599),
.A2(n_1610),
.B1(n_1659),
.B2(n_1657),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1691),
.Y(n_1902)
);

NOR2xp67_ASAP7_75t_L g1903 ( 
.A(n_1660),
.B(n_9),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1701),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1667),
.B(n_1122),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1739),
.A2(n_957),
.B1(n_959),
.B2(n_956),
.C(n_955),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1706),
.Y(n_1907)
);

BUFx8_ASAP7_75t_L g1908 ( 
.A(n_1750),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1674),
.B(n_1687),
.Y(n_1909)
);

AO22x2_ASAP7_75t_L g1910 ( 
.A1(n_1610),
.A2(n_1060),
.B1(n_1064),
.B2(n_1059),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1732),
.Y(n_1911)
);

AO22x2_ASAP7_75t_L g1912 ( 
.A1(n_1657),
.A2(n_1069),
.B1(n_1072),
.B2(n_1068),
.Y(n_1912)
);

NAND2xp33_ASAP7_75t_L g1913 ( 
.A(n_1704),
.B(n_1196),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1727),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1614),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1667),
.B(n_1122),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1738),
.Y(n_1917)
);

NAND2x1p5_ASAP7_75t_L g1918 ( 
.A(n_1709),
.B(n_1138),
.Y(n_1918)
);

AO22x2_ASAP7_75t_L g1919 ( 
.A1(n_1572),
.A2(n_1091),
.B1(n_1094),
.B2(n_1075),
.Y(n_1919)
);

AO22x2_ASAP7_75t_L g1920 ( 
.A1(n_1572),
.A2(n_1120),
.B1(n_1128),
.B2(n_1103),
.Y(n_1920)
);

NAND2x1p5_ASAP7_75t_L g1921 ( 
.A(n_1670),
.B(n_1680),
.Y(n_1921)
);

NOR2xp67_ASAP7_75t_L g1922 ( 
.A(n_1560),
.B(n_9),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1717),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1637),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1614),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1748),
.B(n_1159),
.Y(n_1926)
);

NAND2x1p5_ASAP7_75t_L g1927 ( 
.A(n_1708),
.B(n_1138),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1614),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1574),
.B(n_1590),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1615),
.B(n_1163),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1713),
.B(n_979),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1625),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1611),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1758),
.B(n_980),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1663),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1662),
.B(n_981),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1693),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1702),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1658),
.B(n_988),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1638),
.A2(n_1176),
.B1(n_1184),
.B2(n_1178),
.Y(n_1940)
);

AO22x2_ASAP7_75t_L g1941 ( 
.A1(n_1751),
.A2(n_1190),
.B1(n_1203),
.B2(n_1187),
.Y(n_1941)
);

AO22x2_ASAP7_75t_L g1942 ( 
.A1(n_1562),
.A2(n_1208),
.B1(n_1211),
.B2(n_1205),
.Y(n_1942)
);

AO22x2_ASAP7_75t_L g1943 ( 
.A1(n_1639),
.A2(n_1226),
.B1(n_1227),
.B2(n_1224),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1721),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1742),
.B(n_992),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1595),
.A2(n_995),
.B1(n_996),
.B2(n_993),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1604),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1616),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1620),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1630),
.Y(n_1950)
);

AO22x2_ASAP7_75t_L g1951 ( 
.A1(n_1653),
.A2(n_1247),
.B1(n_1249),
.B2(n_1237),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1758),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1668),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1631),
.Y(n_1954)
);

AO22x2_ASAP7_75t_L g1955 ( 
.A1(n_1638),
.A2(n_1257),
.B1(n_1264),
.B2(n_1256),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1578),
.A2(n_1001),
.B1(n_1014),
.B2(n_999),
.Y(n_1956)
);

NAND2xp33_ASAP7_75t_L g1957 ( 
.A(n_1704),
.B(n_1643),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1744),
.Y(n_1958)
);

NAND2x1p5_ASAP7_75t_L g1959 ( 
.A(n_1603),
.B(n_1269),
.Y(n_1959)
);

OAI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1642),
.A2(n_1024),
.B1(n_1029),
.B2(n_1018),
.C(n_1015),
.Y(n_1960)
);

AO22x2_ASAP7_75t_L g1961 ( 
.A1(n_1719),
.A2(n_1276),
.B1(n_860),
.B2(n_888),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_R g1962 ( 
.A(n_1744),
.B(n_1030),
.Y(n_1962)
);

AO22x2_ASAP7_75t_L g1963 ( 
.A1(n_1606),
.A2(n_860),
.B1(n_888),
.B2(n_855),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1694),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1655),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1654),
.B(n_1042),
.Y(n_1966)
);

BUFx8_ASAP7_75t_L g1967 ( 
.A(n_1677),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1636),
.B(n_1047),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1661),
.Y(n_1969)
);

AO22x2_ASAP7_75t_L g1970 ( 
.A1(n_1564),
.A2(n_1108),
.B1(n_1137),
.B2(n_1104),
.Y(n_1970)
);

OR2x2_ASAP7_75t_SL g1971 ( 
.A(n_1565),
.B(n_1104),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1654),
.B(n_1054),
.Y(n_1972)
);

AND2x2_ASAP7_75t_SL g1973 ( 
.A(n_1634),
.B(n_1146),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1672),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_R g1975 ( 
.A(n_1666),
.B(n_1074),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1677),
.A2(n_1196),
.B1(n_1145),
.B2(n_864),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1666),
.B(n_1080),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1678),
.Y(n_1978)
);

OAI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1753),
.A2(n_1086),
.B1(n_1088),
.B2(n_1085),
.C(n_1084),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1618),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1618),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1845),
.B(n_1954),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1962),
.B(n_1270),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1843),
.B(n_1089),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1818),
.B(n_1093),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1828),
.B(n_1235),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1805),
.B(n_1098),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1780),
.B(n_1241),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1958),
.B(n_1242),
.Y(n_1989)
);

NAND2xp33_ASAP7_75t_SL g1990 ( 
.A(n_1765),
.B(n_858),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_SL g1991 ( 
.A(n_1981),
.B(n_858),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1772),
.B(n_1243),
.Y(n_1992)
);

NAND2xp33_ASAP7_75t_SL g1993 ( 
.A(n_1980),
.B(n_858),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1936),
.B(n_1246),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_SL g1995 ( 
.A(n_1766),
.B(n_1767),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1886),
.B(n_1099),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1776),
.B(n_1253),
.Y(n_1997)
);

NAND2xp33_ASAP7_75t_SL g1998 ( 
.A(n_1769),
.B(n_1200),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1778),
.B(n_1258),
.Y(n_1999)
);

NAND2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1770),
.B(n_1200),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1823),
.B(n_1259),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1975),
.B(n_1260),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1803),
.B(n_1266),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1891),
.B(n_1268),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1889),
.B(n_1896),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1792),
.B(n_1100),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1933),
.B(n_1106),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1764),
.B(n_1110),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1973),
.B(n_1209),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1899),
.B(n_1112),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1902),
.B(n_1113),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1904),
.B(n_1117),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1907),
.B(n_1223),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_SL g2014 ( 
.A(n_1810),
.B(n_864),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1815),
.B(n_1229),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1911),
.B(n_1232),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1923),
.B(n_1233),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1944),
.B(n_1240),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1790),
.B(n_1244),
.Y(n_2019)
);

NAND2xp33_ASAP7_75t_SL g2020 ( 
.A(n_1812),
.B(n_1929),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1783),
.B(n_1125),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1959),
.B(n_1800),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1835),
.B(n_1126),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1908),
.B(n_1185),
.Y(n_2024)
);

NAND2xp33_ASAP7_75t_SL g2025 ( 
.A(n_1791),
.B(n_864),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1875),
.B(n_1186),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1774),
.B(n_1937),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1775),
.B(n_1129),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1786),
.B(n_1248),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1917),
.B(n_1271),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_SL g2031 ( 
.A(n_1839),
.B(n_1133),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1784),
.B(n_1134),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1799),
.B(n_10),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1784),
.B(n_1135),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1903),
.B(n_1201),
.Y(n_2035)
);

NAND2xp33_ASAP7_75t_SL g2036 ( 
.A(n_1909),
.B(n_1139),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1895),
.B(n_1217),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1866),
.B(n_1220),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1968),
.B(n_1168),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1837),
.B(n_1171),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1801),
.B(n_10),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1855),
.B(n_1173),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1931),
.B(n_1174),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1918),
.B(n_1175),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1777),
.B(n_1140),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1804),
.B(n_1141),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1826),
.B(n_1890),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1787),
.B(n_1143),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1946),
.B(n_1198),
.Y(n_2049)
);

NAND2xp33_ASAP7_75t_SL g2050 ( 
.A(n_1797),
.B(n_1149),
.Y(n_2050)
);

NAND2xp33_ASAP7_75t_SL g2051 ( 
.A(n_1952),
.B(n_1154),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1794),
.B(n_1155),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1789),
.B(n_1160),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1811),
.B(n_1161),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1922),
.B(n_1162),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1926),
.B(n_1164),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1807),
.B(n_1813),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1884),
.B(n_1165),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1905),
.B(n_1166),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1916),
.B(n_1167),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_SL g2061 ( 
.A(n_1822),
.B(n_1156),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1862),
.B(n_1180),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1956),
.B(n_1182),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1883),
.B(n_1157),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1825),
.B(n_1172),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1814),
.B(n_1824),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1880),
.B(n_1881),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1771),
.B(n_1145),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1773),
.B(n_1145),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_SL g2070 ( 
.A(n_1850),
.B(n_864),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_1851),
.B(n_982),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1798),
.B(n_11),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1945),
.B(n_1856),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1874),
.B(n_13),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1842),
.B(n_14),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1859),
.B(n_13),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1849),
.B(n_15),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1887),
.B(n_15),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1874),
.B(n_14),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1967),
.B(n_16),
.Y(n_2080)
);

NAND2xp33_ASAP7_75t_SL g2081 ( 
.A(n_1852),
.B(n_14),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1781),
.B(n_16),
.Y(n_2082)
);

NAND2xp33_ASAP7_75t_SL g2083 ( 
.A(n_1858),
.B(n_16),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1782),
.B(n_17),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1817),
.B(n_18),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1930),
.B(n_18),
.Y(n_2086)
);

NAND2xp33_ASAP7_75t_SL g2087 ( 
.A(n_1892),
.B(n_17),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1939),
.B(n_1763),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1853),
.B(n_19),
.Y(n_2089)
);

NAND2xp33_ASAP7_75t_SL g2090 ( 
.A(n_1898),
.B(n_17),
.Y(n_2090)
);

NAND2xp33_ASAP7_75t_SL g2091 ( 
.A(n_1900),
.B(n_19),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1847),
.B(n_21),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1947),
.B(n_20),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1816),
.B(n_20),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1948),
.B(n_21),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1940),
.B(n_23),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1829),
.B(n_1831),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1832),
.B(n_23),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1833),
.B(n_23),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1836),
.B(n_24),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1840),
.B(n_24),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1834),
.B(n_22),
.Y(n_2102)
);

NAND2xp33_ASAP7_75t_SL g2103 ( 
.A(n_1915),
.B(n_22),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1841),
.B(n_25),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1821),
.B(n_24),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1798),
.B(n_25),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1882),
.B(n_27),
.Y(n_2107)
);

NAND2xp33_ASAP7_75t_SL g2108 ( 
.A(n_1925),
.B(n_26),
.Y(n_2108)
);

NAND2xp33_ASAP7_75t_SL g2109 ( 
.A(n_1928),
.B(n_26),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_1865),
.B(n_26),
.Y(n_2110)
);

NAND2xp33_ASAP7_75t_SL g2111 ( 
.A(n_1932),
.B(n_27),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1870),
.B(n_28),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1949),
.B(n_28),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_1950),
.B(n_29),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1921),
.B(n_30),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1927),
.B(n_31),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1901),
.B(n_29),
.Y(n_2117)
);

NAND2xp33_ASAP7_75t_SL g2118 ( 
.A(n_1860),
.B(n_31),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1966),
.B(n_1972),
.Y(n_2119)
);

XNOR2x2_ASAP7_75t_L g2120 ( 
.A(n_1870),
.B(n_33),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_SL g2121 ( 
.A(n_1924),
.B(n_33),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1901),
.B(n_33),
.Y(n_2122)
);

AND2x2_ASAP7_75t_SL g2123 ( 
.A(n_1957),
.B(n_35),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1977),
.B(n_1869),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1953),
.B(n_36),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1872),
.B(n_35),
.Y(n_2126)
);

AND2x4_ASAP7_75t_L g2127 ( 
.A(n_1867),
.B(n_35),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1876),
.B(n_36),
.Y(n_2128)
);

NAND2xp33_ASAP7_75t_SL g2129 ( 
.A(n_1935),
.B(n_38),
.Y(n_2129)
);

XNOR2x2_ASAP7_75t_L g2130 ( 
.A(n_1768),
.B(n_40),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1938),
.B(n_44),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_1871),
.B(n_43),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1897),
.B(n_45),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1876),
.B(n_45),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1838),
.B(n_46),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1964),
.B(n_47),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1872),
.B(n_45),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1857),
.B(n_49),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1827),
.B(n_48),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1873),
.B(n_50),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_SL g2141 ( 
.A(n_1955),
.B(n_48),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1877),
.B(n_50),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_SL g2143 ( 
.A(n_1955),
.B(n_48),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1878),
.B(n_52),
.Y(n_2144)
);

NAND2xp33_ASAP7_75t_SL g2145 ( 
.A(n_1888),
.B(n_51),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_1865),
.B(n_51),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_1795),
.B(n_53),
.Y(n_2147)
);

NAND2xp33_ASAP7_75t_SL g2148 ( 
.A(n_1934),
.B(n_53),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1965),
.B(n_54),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_SL g2150 ( 
.A(n_1793),
.B(n_53),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1827),
.B(n_54),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1844),
.B(n_55),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1844),
.B(n_55),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1969),
.B(n_57),
.Y(n_2154)
);

NAND2xp33_ASAP7_75t_SL g2155 ( 
.A(n_1914),
.B(n_56),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_SL g2156 ( 
.A(n_1846),
.B(n_56),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1974),
.B(n_59),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1978),
.B(n_59),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1863),
.B(n_58),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1863),
.B(n_1864),
.Y(n_2160)
);

NAND2xp33_ASAP7_75t_SL g2161 ( 
.A(n_1848),
.B(n_58),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1864),
.B(n_60),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1941),
.B(n_61),
.Y(n_2163)
);

NAND2xp33_ASAP7_75t_SL g2164 ( 
.A(n_1848),
.B(n_61),
.Y(n_2164)
);

NAND2xp33_ASAP7_75t_SL g2165 ( 
.A(n_1976),
.B(n_61),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1894),
.B(n_63),
.Y(n_2166)
);

NAND2xp33_ASAP7_75t_SL g2167 ( 
.A(n_1963),
.B(n_62),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_SL g2168 ( 
.A(n_1963),
.B(n_62),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1942),
.B(n_1868),
.Y(n_2169)
);

NAND2xp33_ASAP7_75t_SL g2170 ( 
.A(n_1868),
.B(n_62),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1942),
.B(n_65),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1970),
.B(n_65),
.Y(n_2172)
);

NAND2xp33_ASAP7_75t_SL g2173 ( 
.A(n_1788),
.B(n_64),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1941),
.B(n_66),
.Y(n_2174)
);

NAND2xp33_ASAP7_75t_SL g2175 ( 
.A(n_1788),
.B(n_66),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1919),
.B(n_67),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1919),
.B(n_1920),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1854),
.B(n_70),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1920),
.B(n_1893),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1893),
.B(n_70),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1910),
.B(n_71),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1910),
.B(n_71),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1912),
.B(n_72),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_1912),
.B(n_72),
.Y(n_2184)
);

NAND2xp33_ASAP7_75t_SL g2185 ( 
.A(n_1788),
.B(n_67),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1943),
.B(n_73),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1943),
.B(n_75),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1951),
.B(n_75),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1951),
.B(n_76),
.Y(n_2189)
);

NAND2xp33_ASAP7_75t_SL g2190 ( 
.A(n_1885),
.B(n_73),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1906),
.B(n_76),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1971),
.B(n_77),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1879),
.B(n_78),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1762),
.B(n_73),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1885),
.B(n_79),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1885),
.B(n_80),
.Y(n_2196)
);

NAND2xp33_ASAP7_75t_SL g2197 ( 
.A(n_1819),
.B(n_78),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1960),
.B(n_80),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_1819),
.B(n_81),
.Y(n_2199)
);

NAND2xp33_ASAP7_75t_SL g2200 ( 
.A(n_1820),
.B(n_78),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1796),
.B(n_1830),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_1820),
.B(n_82),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1979),
.B(n_82),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_1861),
.B(n_82),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_1802),
.B(n_83),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1761),
.B(n_83),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1785),
.B(n_84),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1809),
.B(n_84),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1809),
.B(n_84),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1808),
.B(n_85),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1808),
.B(n_85),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_1961),
.B(n_81),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1762),
.B(n_87),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1768),
.B(n_88),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1779),
.B(n_88),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_SL g2216 ( 
.A(n_1806),
.B(n_86),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_1806),
.B(n_1913),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1962),
.B(n_90),
.Y(n_2218)
);

NAND2xp33_ASAP7_75t_SL g2219 ( 
.A(n_1962),
.B(n_89),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_1962),
.B(n_90),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_1962),
.B(n_90),
.Y(n_2221)
);

NAND2xp33_ASAP7_75t_SL g2222 ( 
.A(n_1962),
.B(n_89),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1962),
.B(n_93),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1843),
.B(n_91),
.Y(n_2224)
);

AND2x2_ASAP7_75t_SL g2225 ( 
.A(n_1973),
.B(n_91),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1962),
.B(n_93),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_SL g2227 ( 
.A(n_1962),
.B(n_91),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1962),
.B(n_94),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_1962),
.B(n_94),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1843),
.B(n_93),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1958),
.B(n_95),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1962),
.B(n_98),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1962),
.B(n_98),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_1962),
.B(n_98),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1843),
.B(n_96),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1962),
.B(n_99),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1843),
.B(n_96),
.Y(n_2237)
);

NAND2xp33_ASAP7_75t_SL g2238 ( 
.A(n_1962),
.B(n_99),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1843),
.B(n_99),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_1962),
.B(n_101),
.Y(n_2240)
);

NAND2xp33_ASAP7_75t_SL g2241 ( 
.A(n_1962),
.B(n_100),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1962),
.B(n_101),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1962),
.B(n_101),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_SL g2244 ( 
.A(n_1962),
.B(n_102),
.Y(n_2244)
);

NAND2xp33_ASAP7_75t_SL g2245 ( 
.A(n_1962),
.B(n_100),
.Y(n_2245)
);

NAND2xp33_ASAP7_75t_SL g2246 ( 
.A(n_1962),
.B(n_100),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1843),
.B(n_102),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1843),
.B(n_102),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1843),
.B(n_103),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_1962),
.B(n_104),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1962),
.B(n_104),
.Y(n_2251)
);

NAND2xp33_ASAP7_75t_SL g2252 ( 
.A(n_1962),
.B(n_103),
.Y(n_2252)
);

NAND2xp33_ASAP7_75t_SL g2253 ( 
.A(n_1962),
.B(n_104),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_1962),
.B(n_106),
.Y(n_2254)
);

NAND2xp33_ASAP7_75t_SL g2255 ( 
.A(n_1962),
.B(n_105),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_1962),
.B(n_106),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_1843),
.B(n_105),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_1962),
.B(n_107),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_1794),
.B(n_105),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1843),
.B(n_107),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_SL g2261 ( 
.A(n_1845),
.B(n_107),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_1962),
.B(n_109),
.Y(n_2262)
);

NAND2xp33_ASAP7_75t_SL g2263 ( 
.A(n_1845),
.B(n_108),
.Y(n_2263)
);

NAND2xp33_ASAP7_75t_SL g2264 ( 
.A(n_1845),
.B(n_108),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1962),
.B(n_110),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1962),
.B(n_110),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_SL g2267 ( 
.A(n_1845),
.B(n_109),
.Y(n_2267)
);

NAND2xp33_ASAP7_75t_SL g2268 ( 
.A(n_1845),
.B(n_109),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_1962),
.B(n_111),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_1962),
.B(n_111),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_1962),
.B(n_111),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_1962),
.B(n_112),
.Y(n_2272)
);

NAND2xp33_ASAP7_75t_SL g2273 ( 
.A(n_1845),
.B(n_110),
.Y(n_2273)
);

NAND2xp33_ASAP7_75t_SL g2274 ( 
.A(n_1845),
.B(n_112),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1843),
.B(n_112),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1843),
.B(n_113),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1843),
.B(n_113),
.Y(n_2277)
);

NAND2xp33_ASAP7_75t_SL g2278 ( 
.A(n_1845),
.B(n_113),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_1962),
.B(n_115),
.Y(n_2279)
);

NAND2xp33_ASAP7_75t_SL g2280 ( 
.A(n_1845),
.B(n_114),
.Y(n_2280)
);

AND2x4_ASAP7_75t_L g2281 ( 
.A(n_1958),
.B(n_114),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_1958),
.B(n_115),
.Y(n_2282)
);

OR2x2_ASAP7_75t_L g2283 ( 
.A(n_1764),
.B(n_116),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1962),
.B(n_118),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1843),
.B(n_117),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_1962),
.B(n_119),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_1962),
.B(n_119),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_1962),
.B(n_119),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1962),
.B(n_120),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_1962),
.B(n_120),
.Y(n_2290)
);

NAND2xp33_ASAP7_75t_SL g2291 ( 
.A(n_1845),
.B(n_118),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_1958),
.B(n_118),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_1962),
.B(n_122),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_1962),
.B(n_122),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_1962),
.B(n_122),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_1962),
.B(n_123),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_SL g2297 ( 
.A(n_1845),
.B(n_121),
.Y(n_2297)
);

AND2x2_ASAP7_75t_SL g2298 ( 
.A(n_1973),
.B(n_121),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_SL g2299 ( 
.A(n_1845),
.B(n_123),
.Y(n_2299)
);

NAND2xp33_ASAP7_75t_SL g2300 ( 
.A(n_1845),
.B(n_124),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_1962),
.B(n_126),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_1962),
.B(n_126),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_1962),
.B(n_126),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_1962),
.B(n_127),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_1962),
.B(n_127),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_1962),
.B(n_128),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1843),
.B(n_125),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_1962),
.B(n_128),
.Y(n_2308)
);

NAND2xp33_ASAP7_75t_SL g2309 ( 
.A(n_1845),
.B(n_125),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1962),
.B(n_129),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1843),
.B(n_125),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1843),
.B(n_129),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1843),
.B(n_129),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_1962),
.B(n_131),
.Y(n_2314)
);

NAND2xp33_ASAP7_75t_SL g2315 ( 
.A(n_1845),
.B(n_130),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1843),
.B(n_130),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_1843),
.B(n_131),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_1843),
.B(n_132),
.Y(n_2318)
);

NAND2xp33_ASAP7_75t_SL g2319 ( 
.A(n_1845),
.B(n_132),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1843),
.B(n_133),
.Y(n_2320)
);

NAND2xp33_ASAP7_75t_SL g2321 ( 
.A(n_1845),
.B(n_133),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_1962),
.B(n_134),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1843),
.B(n_133),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1962),
.B(n_135),
.Y(n_2324)
);

NAND2xp33_ASAP7_75t_SL g2325 ( 
.A(n_1845),
.B(n_134),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1962),
.B(n_135),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_1962),
.B(n_135),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_1958),
.B(n_134),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_1962),
.B(n_138),
.Y(n_2329)
);

NAND2xp33_ASAP7_75t_SL g2330 ( 
.A(n_1845),
.B(n_136),
.Y(n_2330)
);

NAND2xp33_ASAP7_75t_SL g2331 ( 
.A(n_1845),
.B(n_136),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_1962),
.B(n_139),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_1962),
.B(n_139),
.Y(n_2333)
);

AND2x2_ASAP7_75t_SL g2334 ( 
.A(n_1973),
.B(n_138),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_1962),
.B(n_140),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_1962),
.B(n_140),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1962),
.B(n_140),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1843),
.B(n_139),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_1962),
.B(n_142),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1962),
.B(n_142),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_1962),
.B(n_142),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_1962),
.B(n_143),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1962),
.B(n_143),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_1962),
.B(n_143),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_1843),
.B(n_141),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1843),
.B(n_141),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_1962),
.B(n_144),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_1962),
.B(n_144),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_1962),
.B(n_144),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_1962),
.B(n_145),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_1962),
.B(n_145),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_1845),
.B(n_141),
.Y(n_2352)
);

NAND2xp33_ASAP7_75t_SL g2353 ( 
.A(n_1845),
.B(n_146),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_SL g2354 ( 
.A(n_1845),
.B(n_146),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_1962),
.B(n_147),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1843),
.B(n_146),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1962),
.B(n_148),
.Y(n_2357)
);

NAND2xp33_ASAP7_75t_SL g2358 ( 
.A(n_1845),
.B(n_147),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_SL g2359 ( 
.A(n_1845),
.B(n_147),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_1962),
.B(n_149),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_1962),
.B(n_149),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1962),
.B(n_149),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_1962),
.B(n_151),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_1962),
.B(n_151),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_1962),
.B(n_152),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1843),
.B(n_148),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_1962),
.B(n_153),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_1962),
.B(n_153),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_1962),
.B(n_153),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_1962),
.B(n_154),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_1843),
.B(n_152),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1843),
.B(n_155),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_1843),
.B(n_155),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_SL g2374 ( 
.A(n_1845),
.B(n_155),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_1962),
.B(n_157),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_1962),
.B(n_157),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_1962),
.B(n_157),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1843),
.B(n_156),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_1962),
.B(n_158),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_1962),
.B(n_158),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_1962),
.B(n_159),
.Y(n_2381)
);

NAND2xp33_ASAP7_75t_SL g2382 ( 
.A(n_1845),
.B(n_156),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_1962),
.B(n_160),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_1962),
.B(n_160),
.Y(n_2384)
);

NAND2xp33_ASAP7_75t_SL g2385 ( 
.A(n_1845),
.B(n_159),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_1843),
.B(n_159),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_1962),
.B(n_162),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_1962),
.B(n_162),
.Y(n_2388)
);

NAND2xp33_ASAP7_75t_SL g2389 ( 
.A(n_1845),
.B(n_161),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_1962),
.B(n_163),
.Y(n_2390)
);

NAND2xp33_ASAP7_75t_SL g2391 ( 
.A(n_1845),
.B(n_161),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_1843),
.B(n_163),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1843),
.B(n_164),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_1962),
.B(n_165),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_1962),
.B(n_165),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_1962),
.B(n_165),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_1962),
.B(n_166),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_1962),
.B(n_167),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_1962),
.B(n_167),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_1962),
.B(n_168),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_1962),
.B(n_168),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_1962),
.B(n_168),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_1843),
.B(n_164),
.Y(n_2403)
);

OAI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2225),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2005),
.B(n_169),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2156),
.Y(n_2406)
);

NAND2x1_ASAP7_75t_L g2407 ( 
.A(n_2005),
.B(n_170),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2033),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2005),
.B(n_170),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2201),
.B(n_171),
.Y(n_2410)
);

NOR4xp25_ASAP7_75t_L g2411 ( 
.A(n_2214),
.B(n_2215),
.C(n_2209),
.D(n_2208),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2128),
.B(n_171),
.Y(n_2412)
);

AOI221x1_ASAP7_75t_L g2413 ( 
.A1(n_2141),
.A2(n_2143),
.B1(n_2167),
.B2(n_2168),
.C(n_2216),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2225),
.B(n_218),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2033),
.Y(n_2415)
);

A2O1A1Ixp33_ASAP7_75t_L g2416 ( 
.A1(n_2020),
.A2(n_175),
.B(n_172),
.C(n_173),
.Y(n_2416)
);

AOI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_1990),
.A2(n_172),
.B(n_173),
.Y(n_2417)
);

INVxp67_ASAP7_75t_L g2418 ( 
.A(n_2231),
.Y(n_2418)
);

OAI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2124),
.A2(n_2088),
.B(n_2021),
.Y(n_2419)
);

INVx3_ASAP7_75t_SL g2420 ( 
.A(n_2024),
.Y(n_2420)
);

O2A1O1Ixp5_ASAP7_75t_L g2421 ( 
.A1(n_1990),
.A2(n_178),
.B(n_176),
.C(n_177),
.Y(n_2421)
);

NAND2x1p5_ASAP7_75t_L g2422 ( 
.A(n_2169),
.B(n_177),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2231),
.Y(n_2423)
);

AOI22xp33_ASAP7_75t_L g2424 ( 
.A1(n_2298),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2298),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2425)
);

CKINVDCx20_ASAP7_75t_R g2426 ( 
.A(n_2197),
.Y(n_2426)
);

O2A1O1Ixp5_ASAP7_75t_L g2427 ( 
.A1(n_1991),
.A2(n_1993),
.B(n_2000),
.C(n_1998),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2033),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2008),
.B(n_183),
.Y(n_2429)
);

AOI221xp5_ASAP7_75t_L g2430 ( 
.A1(n_2200),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.C(n_186),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2067),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2057),
.B(n_184),
.Y(n_2432)
);

AO32x2_ASAP7_75t_L g2433 ( 
.A1(n_2120),
.A2(n_187),
.A3(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2334),
.A2(n_188),
.B1(n_185),
.B2(n_187),
.Y(n_2434)
);

INVx4_ASAP7_75t_L g2435 ( 
.A(n_2212),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2134),
.B(n_189),
.Y(n_2436)
);

AOI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2334),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2259),
.B(n_190),
.Y(n_2438)
);

AND3x4_ASAP7_75t_L g2439 ( 
.A(n_2212),
.B(n_191),
.C(n_193),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2130),
.Y(n_2440)
);

NAND3xp33_ASAP7_75t_L g2441 ( 
.A(n_2020),
.B(n_191),
.C(n_194),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2230),
.B(n_194),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_1991),
.A2(n_195),
.B(n_196),
.Y(n_2443)
);

O2A1O1Ixp33_ASAP7_75t_L g2444 ( 
.A1(n_2207),
.A2(n_2073),
.B(n_2211),
.C(n_2210),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2257),
.B(n_195),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2123),
.A2(n_199),
.B1(n_196),
.B2(n_198),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2041),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_1993),
.A2(n_198),
.B(n_199),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2025),
.B(n_221),
.Y(n_2449)
);

NAND3x1_ASAP7_75t_L g2450 ( 
.A(n_2194),
.B(n_199),
.C(n_200),
.Y(n_2450)
);

OAI22x1_ASAP7_75t_L g2451 ( 
.A1(n_2212),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2451)
);

INVx4_ASAP7_75t_L g2452 ( 
.A(n_2041),
.Y(n_2452)
);

OAI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_1996),
.A2(n_203),
.B(n_204),
.Y(n_2453)
);

BUFx12f_ASAP7_75t_L g2454 ( 
.A(n_2147),
.Y(n_2454)
);

NOR2x1_ASAP7_75t_SL g2455 ( 
.A(n_2172),
.B(n_204),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2019),
.B(n_206),
.Y(n_2456)
);

AOI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_1998),
.A2(n_206),
.B(n_207),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2051),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2123),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2041),
.Y(n_2460)
);

INVx1_ASAP7_75t_SL g2461 ( 
.A(n_2231),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_2050),
.Y(n_2462)
);

OAI21xp5_ASAP7_75t_SL g2463 ( 
.A1(n_2112),
.A2(n_208),
.B(n_209),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_2054),
.B(n_209),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2317),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2345),
.B(n_210),
.Y(n_2466)
);

AOI221xp5_ASAP7_75t_SL g2467 ( 
.A1(n_2205),
.A2(n_2187),
.B1(n_2189),
.B2(n_2188),
.C(n_2213),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2000),
.A2(n_212),
.B(n_213),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2027),
.B(n_212),
.Y(n_2469)
);

OR2x6_ASAP7_75t_L g2470 ( 
.A(n_2281),
.B(n_213),
.Y(n_2470)
);

NAND3xp33_ASAP7_75t_SL g2471 ( 
.A(n_2150),
.B(n_214),
.C(n_215),
.Y(n_2471)
);

OAI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2010),
.A2(n_214),
.B(n_215),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2373),
.B(n_216),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_SL g2474 ( 
.A1(n_2127),
.A2(n_216),
.B(n_222),
.Y(n_2474)
);

OAI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2011),
.A2(n_222),
.B(n_223),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2386),
.Y(n_2476)
);

BUFx10_ASAP7_75t_L g2477 ( 
.A(n_2281),
.Y(n_2477)
);

A2O1A1Ixp33_ASAP7_75t_L g2478 ( 
.A1(n_2025),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2392),
.Y(n_2479)
);

AOI21xp33_ASAP7_75t_L g2480 ( 
.A1(n_2052),
.A2(n_225),
.B(n_226),
.Y(n_2480)
);

AOI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2170),
.A2(n_2006),
.B1(n_2160),
.B2(n_2179),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2127),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2133),
.B(n_229),
.Y(n_2483)
);

AO31x2_ASAP7_75t_L g2484 ( 
.A1(n_2074),
.A2(n_233),
.A3(n_230),
.B(n_232),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2127),
.Y(n_2485)
);

INVxp67_ASAP7_75t_SL g2486 ( 
.A(n_2132),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2012),
.A2(n_233),
.B(n_234),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2132),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_2177),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2132),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2281),
.Y(n_2491)
);

AO31x2_ASAP7_75t_L g2492 ( 
.A1(n_2079),
.A2(n_2137),
.A3(n_2126),
.B(n_2186),
.Y(n_2492)
);

AOI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_2014),
.A2(n_239),
.B(n_241),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2224),
.B(n_242),
.Y(n_2494)
);

INVx4_ASAP7_75t_L g2495 ( 
.A(n_2282),
.Y(n_2495)
);

NAND2xp33_ASAP7_75t_R g2496 ( 
.A(n_2282),
.B(n_242),
.Y(n_2496)
);

OAI22x1_ASAP7_75t_L g2497 ( 
.A1(n_2199),
.A2(n_245),
.B1(n_246),
.B2(n_244),
.Y(n_2497)
);

OAI22x1_ASAP7_75t_L g2498 ( 
.A1(n_2202),
.A2(n_245),
.B1(n_246),
.B2(n_244),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2022),
.B(n_243),
.Y(n_2499)
);

BUFx3_ASAP7_75t_L g2500 ( 
.A(n_2282),
.Y(n_2500)
);

NAND3x1_ASAP7_75t_L g2501 ( 
.A(n_2072),
.B(n_248),
.C(n_250),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2235),
.B(n_250),
.Y(n_2502)
);

OR2x6_ASAP7_75t_L g2503 ( 
.A(n_2292),
.B(n_251),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2292),
.Y(n_2504)
);

AO22x1_ASAP7_75t_L g2505 ( 
.A1(n_2106),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_2505)
);

AOI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2014),
.A2(n_254),
.B(n_256),
.Y(n_2506)
);

OAI22xp5_ASAP7_75t_L g2507 ( 
.A1(n_2093),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_2507)
);

O2A1O1Ixp33_ASAP7_75t_L g2508 ( 
.A1(n_2206),
.A2(n_261),
.B(n_258),
.C(n_260),
.Y(n_2508)
);

AOI22xp33_ASAP7_75t_L g2509 ( 
.A1(n_2032),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2283),
.B(n_263),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_SL g2511 ( 
.A1(n_2093),
.A2(n_2113),
.B(n_2095),
.Y(n_2511)
);

BUFx6f_ASAP7_75t_L g2512 ( 
.A(n_2292),
.Y(n_2512)
);

AOI21xp5_ASAP7_75t_L g2513 ( 
.A1(n_2070),
.A2(n_2071),
.B(n_2119),
.Y(n_2513)
);

BUFx2_ASAP7_75t_L g2514 ( 
.A(n_2061),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2237),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_2155),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2328),
.Y(n_2517)
);

AOI21xp5_ASAP7_75t_L g2518 ( 
.A1(n_1995),
.A2(n_2069),
.B(n_2068),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2239),
.Y(n_2519)
);

OAI22xp33_ASAP7_75t_L g2520 ( 
.A1(n_2110),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2247),
.B(n_268),
.Y(n_2521)
);

OAI21x1_ASAP7_75t_SL g2522 ( 
.A1(n_2163),
.A2(n_2174),
.B(n_2122),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2328),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2328),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2093),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2219),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2248),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_1987),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2528)
);

NOR2xp67_ASAP7_75t_L g2529 ( 
.A(n_2003),
.B(n_275),
.Y(n_2529)
);

BUFx2_ASAP7_75t_L g2530 ( 
.A(n_2222),
.Y(n_2530)
);

AO31x2_ASAP7_75t_L g2531 ( 
.A1(n_2117),
.A2(n_278),
.A3(n_275),
.B(n_277),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2403),
.B(n_278),
.Y(n_2532)
);

OAI22x1_ASAP7_75t_L g2533 ( 
.A1(n_2217),
.A2(n_2180),
.B1(n_2182),
.B2(n_2181),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2249),
.B(n_279),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2260),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2275),
.B(n_280),
.Y(n_2536)
);

AO21x2_ASAP7_75t_L g2537 ( 
.A1(n_2171),
.A2(n_281),
.B(n_282),
.Y(n_2537)
);

OAI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_1984),
.A2(n_283),
.B(n_284),
.Y(n_2538)
);

BUFx6f_ASAP7_75t_L g2539 ( 
.A(n_2095),
.Y(n_2539)
);

NOR2xp67_ASAP7_75t_L g2540 ( 
.A(n_2001),
.B(n_285),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2276),
.B(n_285),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2113),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2277),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2113),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2097),
.Y(n_2545)
);

INVx3_ASAP7_75t_SL g2546 ( 
.A(n_2166),
.Y(n_2546)
);

A2O1A1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2261),
.A2(n_2264),
.B(n_2267),
.C(n_2263),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2285),
.B(n_287),
.Y(n_2548)
);

OAI21x1_ASAP7_75t_SL g2549 ( 
.A1(n_2139),
.A2(n_288),
.B(n_289),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2307),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2311),
.Y(n_2551)
);

NOR2xp67_ASAP7_75t_SL g2552 ( 
.A(n_2183),
.B(n_290),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2312),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2313),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2316),
.Y(n_2555)
);

A2O1A1Ixp33_ASAP7_75t_L g2556 ( 
.A1(n_2263),
.A2(n_298),
.B(n_295),
.C(n_297),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2318),
.B(n_299),
.Y(n_2557)
);

NAND3xp33_ASAP7_75t_L g2558 ( 
.A(n_2264),
.B(n_300),
.C(n_301),
.Y(n_2558)
);

AOI221x1_ASAP7_75t_L g2559 ( 
.A1(n_2161),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.C(n_305),
.Y(n_2559)
);

AO32x2_ASAP7_75t_L g2560 ( 
.A1(n_2164),
.A2(n_305),
.A3(n_303),
.B1(n_304),
.B2(n_306),
.Y(n_2560)
);

BUFx3_ASAP7_75t_L g2561 ( 
.A(n_2114),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2320),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2075),
.A2(n_2078),
.B(n_2077),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2323),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2338),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2114),
.Y(n_2566)
);

INVx1_ASAP7_75t_SL g2567 ( 
.A(n_2114),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2056),
.B(n_310),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2346),
.B(n_2356),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2047),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2366),
.B(n_311),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2371),
.Y(n_2572)
);

AO32x2_ASAP7_75t_L g2573 ( 
.A1(n_2267),
.A2(n_316),
.A3(n_314),
.B1(n_315),
.B2(n_317),
.Y(n_2573)
);

OAI21x1_ASAP7_75t_SL g2574 ( 
.A1(n_2151),
.A2(n_314),
.B(n_315),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2372),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2378),
.A2(n_316),
.B(n_317),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2393),
.B(n_318),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2066),
.B(n_2058),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2082),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2015),
.B(n_321),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2084),
.Y(n_2581)
);

BUFx10_ASAP7_75t_L g2582 ( 
.A(n_2146),
.Y(n_2582)
);

NOR3xp33_ASAP7_75t_SL g2583 ( 
.A(n_2227),
.B(n_323),
.C(n_324),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2094),
.B(n_323),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2105),
.B(n_324),
.Y(n_2585)
);

NAND3xp33_ASAP7_75t_L g2586 ( 
.A(n_2268),
.B(n_2274),
.C(n_2273),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2116),
.Y(n_2587)
);

AO21x1_ASAP7_75t_L g2588 ( 
.A1(n_2268),
.A2(n_325),
.B(n_326),
.Y(n_2588)
);

OR2x2_ASAP7_75t_L g2589 ( 
.A(n_2034),
.B(n_326),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_2178),
.Y(n_2590)
);

OAI21xp5_ASAP7_75t_L g2591 ( 
.A1(n_2204),
.A2(n_330),
.B(n_331),
.Y(n_2591)
);

OA21x2_ASAP7_75t_L g2592 ( 
.A1(n_2089),
.A2(n_332),
.B(n_333),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2152),
.Y(n_2593)
);

INVx2_ASAP7_75t_SL g2594 ( 
.A(n_2026),
.Y(n_2594)
);

BUFx4_ASAP7_75t_SL g2595 ( 
.A(n_2080),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2086),
.B(n_334),
.Y(n_2596)
);

INVxp67_ASAP7_75t_L g2597 ( 
.A(n_2102),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2092),
.B(n_335),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2153),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2238),
.Y(n_2600)
);

INVx1_ASAP7_75t_SL g2601 ( 
.A(n_2241),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2184),
.B(n_339),
.Y(n_2602)
);

AOI21x1_ASAP7_75t_SL g2603 ( 
.A1(n_2176),
.A2(n_2162),
.B(n_2159),
.Y(n_2603)
);

INVxp67_ASAP7_75t_L g2604 ( 
.A(n_2118),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2028),
.B(n_340),
.Y(n_2605)
);

OAI22x1_ASAP7_75t_L g2606 ( 
.A1(n_2193),
.A2(n_346),
.B1(n_347),
.B2(n_345),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2045),
.B(n_344),
.Y(n_2607)
);

BUFx3_ASAP7_75t_L g2608 ( 
.A(n_2076),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2036),
.A2(n_347),
.B1(n_344),
.B2(n_346),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2198),
.A2(n_348),
.B(n_349),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_1988),
.B(n_350),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_L g2612 ( 
.A(n_2062),
.B(n_351),
.Y(n_2612)
);

NOR2xp67_ASAP7_75t_L g2613 ( 
.A(n_1983),
.B(n_351),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2273),
.B(n_2274),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2046),
.B(n_353),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2039),
.B(n_354),
.Y(n_2616)
);

OA22x2_ASAP7_75t_L g2617 ( 
.A1(n_2218),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_2617)
);

OAI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2192),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_2618)
);

A2O1A1Ixp33_ASAP7_75t_L g2619 ( 
.A1(n_2278),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2098),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2085),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_R g2622 ( 
.A(n_2245),
.B(n_370),
.Y(n_2622)
);

NOR2xp67_ASAP7_75t_SL g2623 ( 
.A(n_2195),
.B(n_371),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2064),
.B(n_2191),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2135),
.B(n_374),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2280),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2029),
.B(n_378),
.Y(n_2627)
);

AO31x2_ASAP7_75t_L g2628 ( 
.A1(n_2280),
.A2(n_380),
.A3(n_378),
.B(n_379),
.Y(n_2628)
);

AND2x2_ASAP7_75t_L g2629 ( 
.A(n_2402),
.B(n_381),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2291),
.B(n_382),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2291),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2099),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2297),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2220),
.B(n_386),
.Y(n_2634)
);

OAI21x1_ASAP7_75t_SL g2635 ( 
.A1(n_2297),
.A2(n_387),
.B(n_388),
.Y(n_2635)
);

AOI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_1982),
.A2(n_388),
.B(n_389),
.Y(n_2636)
);

AO31x2_ASAP7_75t_L g2637 ( 
.A1(n_2299),
.A2(n_391),
.A3(n_389),
.B(n_390),
.Y(n_2637)
);

OAI21xp5_ASAP7_75t_L g2638 ( 
.A1(n_2203),
.A2(n_391),
.B(n_393),
.Y(n_2638)
);

AO21x2_ASAP7_75t_L g2639 ( 
.A1(n_2131),
.A2(n_393),
.B(n_394),
.Y(n_2639)
);

BUFx12f_ASAP7_75t_L g2640 ( 
.A(n_2246),
.Y(n_2640)
);

OAI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2096),
.A2(n_394),
.B(n_395),
.Y(n_2641)
);

INVx4_ASAP7_75t_SL g2642 ( 
.A(n_2252),
.Y(n_2642)
);

AOI21xp5_ASAP7_75t_SL g2643 ( 
.A1(n_2196),
.A2(n_395),
.B(n_396),
.Y(n_2643)
);

A2O1A1Ixp33_ASAP7_75t_L g2644 ( 
.A1(n_2299),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_2644)
);

AOI21xp33_ASAP7_75t_L g2645 ( 
.A1(n_2035),
.A2(n_397),
.B(n_398),
.Y(n_2645)
);

AND2x4_ASAP7_75t_L g2646 ( 
.A(n_2059),
.B(n_399),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_1994),
.B(n_401),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2100),
.Y(n_2648)
);

A2O1A1Ixp33_ASAP7_75t_L g2649 ( 
.A1(n_2300),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_2649)
);

INVx6_ASAP7_75t_L g2650 ( 
.A(n_2253),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2017),
.B(n_408),
.Y(n_2651)
);

AO31x2_ASAP7_75t_L g2652 ( 
.A1(n_2300),
.A2(n_411),
.A3(n_409),
.B(n_410),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2060),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2221),
.B(n_412),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2018),
.B(n_414),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2101),
.Y(n_2656)
);

AO31x2_ASAP7_75t_L g2657 ( 
.A1(n_2309),
.A2(n_417),
.A3(n_415),
.B(n_416),
.Y(n_2657)
);

AOI21xp5_ASAP7_75t_L g2658 ( 
.A1(n_2309),
.A2(n_416),
.B(n_418),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2009),
.A2(n_2104),
.B1(n_2142),
.B2(n_2140),
.Y(n_2659)
);

AOI21xp5_ASAP7_75t_L g2660 ( 
.A1(n_2315),
.A2(n_418),
.B(n_419),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2149),
.Y(n_2661)
);

A2O1A1Ixp33_ASAP7_75t_L g2662 ( 
.A1(n_2315),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2013),
.B(n_420),
.Y(n_2663)
);

INVxp67_ASAP7_75t_SL g2664 ( 
.A(n_2107),
.Y(n_2664)
);

INVx4_ASAP7_75t_L g2665 ( 
.A(n_2319),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2223),
.B(n_423),
.Y(n_2666)
);

AOI21xp5_ASAP7_75t_L g2667 ( 
.A1(n_2319),
.A2(n_424),
.B(n_426),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2154),
.Y(n_2668)
);

CKINVDCx20_ASAP7_75t_R g2669 ( 
.A(n_2255),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2157),
.Y(n_2670)
);

INVx4_ASAP7_75t_L g2671 ( 
.A(n_2321),
.Y(n_2671)
);

AOI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2321),
.A2(n_427),
.B(n_428),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2144),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2158),
.A2(n_429),
.B(n_430),
.Y(n_2674)
);

OAI22x1_ASAP7_75t_L g2675 ( 
.A1(n_2226),
.A2(n_434),
.B1(n_430),
.B2(n_432),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_1999),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2115),
.Y(n_2677)
);

OAI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2125),
.A2(n_435),
.B(n_436),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2030),
.Y(n_2679)
);

AOI221xp5_ASAP7_75t_L g2680 ( 
.A1(n_2325),
.A2(n_439),
.B1(n_436),
.B2(n_437),
.C(n_440),
.Y(n_2680)
);

AO31x2_ASAP7_75t_L g2681 ( 
.A1(n_2325),
.A2(n_440),
.A3(n_437),
.B(n_439),
.Y(n_2681)
);

AO31x2_ASAP7_75t_L g2682 ( 
.A1(n_2330),
.A2(n_443),
.A3(n_441),
.B(n_442),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2048),
.B(n_441),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2044),
.B(n_2016),
.Y(n_2684)
);

BUFx12f_ASAP7_75t_L g2685 ( 
.A(n_2038),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2040),
.B(n_442),
.Y(n_2686)
);

NAND2x1_ASAP7_75t_L g2687 ( 
.A(n_2173),
.B(n_443),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2330),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2331),
.A2(n_444),
.B(n_446),
.Y(n_2689)
);

OR2x6_ASAP7_75t_L g2690 ( 
.A(n_2228),
.B(n_446),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2352),
.B(n_447),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2136),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2138),
.Y(n_2693)
);

BUFx10_ASAP7_75t_L g2694 ( 
.A(n_2031),
.Y(n_2694)
);

AOI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2353),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_2695)
);

AO31x2_ASAP7_75t_L g2696 ( 
.A1(n_2353),
.A2(n_451),
.A3(n_449),
.B(n_450),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2354),
.Y(n_2697)
);

NAND3xp33_ASAP7_75t_SL g2698 ( 
.A(n_2229),
.B(n_452),
.C(n_453),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2354),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2358),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2037),
.B(n_454),
.Y(n_2701)
);

A2O1A1Ixp33_ASAP7_75t_L g2702 ( 
.A1(n_2359),
.A2(n_458),
.B(n_456),
.C(n_457),
.Y(n_2702)
);

INVx4_ASAP7_75t_L g2703 ( 
.A(n_2359),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2374),
.Y(n_2704)
);

NOR2x1_ASAP7_75t_L g2705 ( 
.A(n_2232),
.B(n_2233),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2374),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2065),
.B(n_2042),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2382),
.A2(n_458),
.B(n_459),
.Y(n_2708)
);

AOI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2382),
.A2(n_459),
.B(n_460),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2043),
.B(n_460),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2004),
.B(n_461),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2385),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2007),
.B(n_461),
.Y(n_2713)
);

BUFx2_ASAP7_75t_R g2714 ( 
.A(n_2234),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2053),
.B(n_2049),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2385),
.A2(n_463),
.B(n_464),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2389),
.B(n_465),
.Y(n_2717)
);

AND2x4_ASAP7_75t_L g2718 ( 
.A(n_2055),
.B(n_465),
.Y(n_2718)
);

BUFx12f_ASAP7_75t_L g2719 ( 
.A(n_2236),
.Y(n_2719)
);

OAI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2240),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_SL g2721 ( 
.A1(n_2391),
.A2(n_470),
.B(n_474),
.Y(n_2721)
);

OAI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2063),
.A2(n_475),
.B(n_476),
.Y(n_2722)
);

A2O1A1Ixp33_ASAP7_75t_L g2723 ( 
.A1(n_2081),
.A2(n_478),
.B(n_476),
.C(n_477),
.Y(n_2723)
);

NOR2x1_ASAP7_75t_L g2724 ( 
.A(n_2242),
.B(n_478),
.Y(n_2724)
);

OAI21x1_ASAP7_75t_SL g2725 ( 
.A1(n_2083),
.A2(n_479),
.B(n_481),
.Y(n_2725)
);

AOI211x1_ASAP7_75t_L g2726 ( 
.A1(n_2243),
.A2(n_2250),
.B(n_2251),
.C(n_2244),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2023),
.B(n_479),
.Y(n_2727)
);

NAND2xp33_ASAP7_75t_L g2728 ( 
.A(n_2175),
.B(n_481),
.Y(n_2728)
);

A2O1A1Ixp33_ASAP7_75t_L g2729 ( 
.A1(n_2121),
.A2(n_484),
.B(n_482),
.C(n_483),
.Y(n_2729)
);

AO21x1_ASAP7_75t_L g2730 ( 
.A1(n_2087),
.A2(n_485),
.B(n_486),
.Y(n_2730)
);

A2O1A1Ixp33_ASAP7_75t_L g2731 ( 
.A1(n_2129),
.A2(n_489),
.B(n_487),
.C(n_488),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2002),
.Y(n_2732)
);

INVx1_ASAP7_75t_SL g2733 ( 
.A(n_2090),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2254),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2091),
.A2(n_493),
.B(n_490),
.C(n_492),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2091),
.Y(n_2736)
);

AO31x2_ASAP7_75t_L g2737 ( 
.A1(n_2103),
.A2(n_495),
.A3(n_493),
.B(n_494),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_SL g2738 ( 
.A(n_2185),
.B(n_494),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_1992),
.B(n_495),
.Y(n_2739)
);

AOI22xp5_ASAP7_75t_L g2740 ( 
.A1(n_2145),
.A2(n_498),
.B1(n_496),
.B2(n_497),
.Y(n_2740)
);

CKINVDCx11_ASAP7_75t_R g2741 ( 
.A(n_2256),
.Y(n_2741)
);

OAI21xp5_ASAP7_75t_SL g2742 ( 
.A1(n_2258),
.A2(n_497),
.B(n_498),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2262),
.B(n_500),
.Y(n_2743)
);

INVx3_ASAP7_75t_L g2744 ( 
.A(n_2103),
.Y(n_2744)
);

OA21x2_ASAP7_75t_L g2745 ( 
.A1(n_2265),
.A2(n_502),
.B(n_503),
.Y(n_2745)
);

INVxp67_ASAP7_75t_SL g2746 ( 
.A(n_2266),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2108),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2165),
.A2(n_504),
.B(n_505),
.Y(n_2748)
);

NOR2x1_ASAP7_75t_SL g2749 ( 
.A(n_2269),
.B(n_504),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2270),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2271),
.Y(n_2751)
);

AO31x2_ASAP7_75t_L g2752 ( 
.A1(n_2108),
.A2(n_508),
.A3(n_506),
.B(n_507),
.Y(n_2752)
);

OAI21x1_ASAP7_75t_SL g2753 ( 
.A1(n_2109),
.A2(n_506),
.B(n_507),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2272),
.B(n_511),
.Y(n_2754)
);

INVx3_ASAP7_75t_SL g2755 ( 
.A(n_2401),
.Y(n_2755)
);

AOI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2148),
.A2(n_516),
.B1(n_512),
.B2(n_513),
.Y(n_2756)
);

BUFx8_ASAP7_75t_L g2757 ( 
.A(n_2279),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2284),
.Y(n_2758)
);

BUFx12f_ASAP7_75t_L g2759 ( 
.A(n_2685),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2688),
.Y(n_2760)
);

OA21x2_ASAP7_75t_L g2761 ( 
.A1(n_2547),
.A2(n_2287),
.B(n_2286),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_SL g2762 ( 
.A1(n_2665),
.A2(n_2190),
.B1(n_2111),
.B2(n_2109),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2700),
.Y(n_2763)
);

OAI21x1_ASAP7_75t_L g2764 ( 
.A1(n_2427),
.A2(n_2289),
.B(n_2288),
.Y(n_2764)
);

AOI21xp5_ASAP7_75t_L g2765 ( 
.A1(n_2513),
.A2(n_2111),
.B(n_2290),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2704),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2706),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2431),
.B(n_2293),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2593),
.B(n_2294),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2595),
.Y(n_2770)
);

AOI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2511),
.A2(n_2296),
.B(n_2295),
.Y(n_2771)
);

AO31x2_ASAP7_75t_L g2772 ( 
.A1(n_2413),
.A2(n_2302),
.A3(n_2303),
.B(n_2301),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2412),
.B(n_2304),
.Y(n_2773)
);

AND2x2_ASAP7_75t_SL g2774 ( 
.A(n_2435),
.B(n_2305),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2436),
.B(n_2306),
.Y(n_2775)
);

BUFx6f_ASAP7_75t_L g2776 ( 
.A(n_2504),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2470),
.B(n_2308),
.Y(n_2777)
);

OAI21x1_ASAP7_75t_L g2778 ( 
.A1(n_2603),
.A2(n_2314),
.B(n_2310),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2551),
.Y(n_2779)
);

OAI21x1_ASAP7_75t_SL g2780 ( 
.A1(n_2435),
.A2(n_2324),
.B(n_2322),
.Y(n_2780)
);

OAI21x1_ASAP7_75t_L g2781 ( 
.A1(n_2518),
.A2(n_2327),
.B(n_2326),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2459),
.B(n_2329),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_2420),
.Y(n_2783)
);

HB1xp67_ASAP7_75t_L g2784 ( 
.A(n_2470),
.Y(n_2784)
);

OAI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2496),
.A2(n_2333),
.B1(n_2335),
.B2(n_2332),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2459),
.A2(n_2400),
.B1(n_2337),
.B2(n_2339),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_SL g2787 ( 
.A(n_2503),
.Y(n_2787)
);

OAI21x1_ASAP7_75t_L g2788 ( 
.A1(n_2744),
.A2(n_2340),
.B(n_2336),
.Y(n_2788)
);

AOI22x1_ASAP7_75t_L g2789 ( 
.A1(n_2665),
.A2(n_2342),
.B1(n_2343),
.B2(n_2341),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2712),
.Y(n_2790)
);

OAI21x1_ASAP7_75t_L g2791 ( 
.A1(n_2744),
.A2(n_2347),
.B(n_2344),
.Y(n_2791)
);

BUFx4f_ASAP7_75t_SL g2792 ( 
.A(n_2454),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2459),
.A2(n_2399),
.B1(n_2349),
.B2(n_2350),
.Y(n_2793)
);

OR2x2_ASAP7_75t_L g2794 ( 
.A(n_2510),
.B(n_2348),
.Y(n_2794)
);

OAI21x1_ASAP7_75t_L g2795 ( 
.A1(n_2747),
.A2(n_2355),
.B(n_2351),
.Y(n_2795)
);

OAI21x1_ASAP7_75t_L g2796 ( 
.A1(n_2747),
.A2(n_2360),
.B(n_2357),
.Y(n_2796)
);

OAI21x1_ASAP7_75t_L g2797 ( 
.A1(n_2626),
.A2(n_2362),
.B(n_2361),
.Y(n_2797)
);

OAI21x1_ASAP7_75t_L g2798 ( 
.A1(n_2626),
.A2(n_2364),
.B(n_2363),
.Y(n_2798)
);

OAI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2503),
.A2(n_2367),
.B1(n_2368),
.B2(n_2365),
.Y(n_2799)
);

OR2x6_ASAP7_75t_L g2800 ( 
.A(n_2474),
.B(n_2369),
.Y(n_2800)
);

AO21x2_ASAP7_75t_L g2801 ( 
.A1(n_2522),
.A2(n_2375),
.B(n_2370),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2555),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2628),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2429),
.B(n_2376),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2486),
.A2(n_2379),
.B(n_2377),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2599),
.B(n_2380),
.Y(n_2806)
);

CKINVDCx20_ASAP7_75t_R g2807 ( 
.A(n_2546),
.Y(n_2807)
);

AOI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2414),
.A2(n_2398),
.B1(n_2383),
.B2(n_2384),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2406),
.B(n_2381),
.Y(n_2809)
);

OAI21x1_ASAP7_75t_L g2810 ( 
.A1(n_2631),
.A2(n_2388),
.B(n_2387),
.Y(n_2810)
);

AOI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2439),
.A2(n_2394),
.B1(n_2395),
.B2(n_2390),
.Y(n_2811)
);

INVx3_ASAP7_75t_L g2812 ( 
.A(n_2452),
.Y(n_2812)
);

AO21x2_ASAP7_75t_L g2813 ( 
.A1(n_2614),
.A2(n_2397),
.B(n_2396),
.Y(n_2813)
);

AO31x2_ASAP7_75t_L g2814 ( 
.A1(n_2533),
.A2(n_518),
.A3(n_516),
.B(n_517),
.Y(n_2814)
);

AO32x2_ASAP7_75t_L g2815 ( 
.A1(n_2446),
.A2(n_520),
.A3(n_517),
.B1(n_519),
.B2(n_521),
.Y(n_2815)
);

AO21x2_ASAP7_75t_L g2816 ( 
.A1(n_2586),
.A2(n_1986),
.B(n_1985),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2465),
.B(n_1997),
.Y(n_2817)
);

OR2x6_ASAP7_75t_L g2818 ( 
.A(n_2452),
.B(n_2640),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2572),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2728),
.A2(n_1989),
.B(n_519),
.Y(n_2820)
);

OR2x2_ASAP7_75t_SL g2821 ( 
.A(n_2471),
.B(n_520),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2476),
.B(n_522),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2504),
.Y(n_2823)
);

AO21x2_ASAP7_75t_L g2824 ( 
.A1(n_2635),
.A2(n_522),
.B(n_523),
.Y(n_2824)
);

NAND3xp33_ASAP7_75t_L g2825 ( 
.A(n_2583),
.B(n_524),
.C(n_525),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2504),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2671),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2581),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2637),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2495),
.B(n_527),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2463),
.B(n_528),
.Y(n_2831)
);

OAI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2421),
.A2(n_529),
.B(n_530),
.Y(n_2832)
);

AOI21x1_ASAP7_75t_L g2833 ( 
.A1(n_2697),
.A2(n_531),
.B(n_532),
.Y(n_2833)
);

OAI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2563),
.A2(n_532),
.B(n_533),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2637),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2637),
.Y(n_2836)
);

OAI211xp5_ASAP7_75t_L g2837 ( 
.A1(n_2622),
.A2(n_536),
.B(n_533),
.C(n_535),
.Y(n_2837)
);

OR2x2_ASAP7_75t_L g2838 ( 
.A(n_2589),
.B(n_535),
.Y(n_2838)
);

OAI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2419),
.A2(n_536),
.B(n_537),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2652),
.Y(n_2840)
);

O2A1O1Ixp33_ASAP7_75t_L g2841 ( 
.A1(n_2410),
.A2(n_540),
.B(n_538),
.C(n_539),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2679),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2652),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2495),
.B(n_541),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2449),
.A2(n_542),
.B(n_543),
.Y(n_2845)
);

BUFx12f_ASAP7_75t_L g2846 ( 
.A(n_2741),
.Y(n_2846)
);

OA21x2_ASAP7_75t_L g2847 ( 
.A1(n_2467),
.A2(n_542),
.B(n_543),
.Y(n_2847)
);

NAND2x1p5_ASAP7_75t_L g2848 ( 
.A(n_2458),
.B(n_2500),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2733),
.A2(n_545),
.B(n_546),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2569),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_2850)
);

CKINVDCx5p33_ASAP7_75t_R g2851 ( 
.A(n_2732),
.Y(n_2851)
);

OAI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2437),
.A2(n_553),
.B1(n_549),
.B2(n_551),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2652),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2515),
.Y(n_2854)
);

INVx2_ASAP7_75t_SL g2855 ( 
.A(n_2694),
.Y(n_2855)
);

AO21x2_ASAP7_75t_L g2856 ( 
.A1(n_2753),
.A2(n_553),
.B(n_554),
.Y(n_2856)
);

INVxp33_ASAP7_75t_L g2857 ( 
.A(n_2514),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_L g2858 ( 
.A(n_2755),
.B(n_555),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2694),
.Y(n_2859)
);

INVxp67_ASAP7_75t_L g2860 ( 
.A(n_2456),
.Y(n_2860)
);

AO31x2_ASAP7_75t_L g2861 ( 
.A1(n_2588),
.A2(n_558),
.A3(n_556),
.B(n_557),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2657),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2657),
.Y(n_2863)
);

O2A1O1Ixp33_ASAP7_75t_SL g2864 ( 
.A1(n_2478),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2590),
.B(n_562),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2671),
.A2(n_562),
.B(n_563),
.Y(n_2866)
);

INVx1_ASAP7_75t_SL g2867 ( 
.A(n_2676),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2479),
.B(n_848),
.Y(n_2868)
);

OAI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2441),
.A2(n_564),
.B(n_565),
.Y(n_2869)
);

A2O1A1Ixp33_ASAP7_75t_L g2870 ( 
.A1(n_2417),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_2870)
);

CKINVDCx8_ASAP7_75t_R g2871 ( 
.A(n_2516),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2519),
.B(n_567),
.Y(n_2872)
);

AO31x2_ASAP7_75t_L g2873 ( 
.A1(n_2730),
.A2(n_570),
.A3(n_568),
.B(n_569),
.Y(n_2873)
);

AOI21x1_ASAP7_75t_L g2874 ( 
.A1(n_2630),
.A2(n_570),
.B(n_571),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2527),
.B(n_2535),
.Y(n_2875)
);

AOI22xp33_ASAP7_75t_L g2876 ( 
.A1(n_2569),
.A2(n_576),
.B1(n_572),
.B2(n_574),
.Y(n_2876)
);

OAI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2624),
.A2(n_574),
.B(n_576),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_SL g2878 ( 
.A(n_2462),
.B(n_577),
.Y(n_2878)
);

NOR2xp67_ASAP7_75t_L g2879 ( 
.A(n_2703),
.B(n_578),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2451),
.Y(n_2880)
);

AOI21x1_ASAP7_75t_L g2881 ( 
.A1(n_2691),
.A2(n_579),
.B(n_580),
.Y(n_2881)
);

OAI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2591),
.A2(n_581),
.B(n_582),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_L g2883 ( 
.A(n_2523),
.Y(n_2883)
);

AOI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2717),
.A2(n_581),
.B(n_582),
.Y(n_2884)
);

OAI21x1_ASAP7_75t_SL g2885 ( 
.A1(n_2703),
.A2(n_2455),
.B(n_2725),
.Y(n_2885)
);

OR2x6_ASAP7_75t_L g2886 ( 
.A(n_2650),
.B(n_583),
.Y(n_2886)
);

NAND3xp33_ASAP7_75t_L g2887 ( 
.A(n_2559),
.B(n_584),
.C(n_585),
.Y(n_2887)
);

OR2x6_ASAP7_75t_L g2888 ( 
.A(n_2650),
.B(n_584),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2681),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2543),
.B(n_2550),
.Y(n_2890)
);

BUFx2_ASAP7_75t_L g2891 ( 
.A(n_2512),
.Y(n_2891)
);

OAI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2424),
.A2(n_591),
.B1(n_586),
.B2(n_589),
.Y(n_2892)
);

INVx3_ASAP7_75t_L g2893 ( 
.A(n_2699),
.Y(n_2893)
);

CKINVDCx12_ASAP7_75t_R g2894 ( 
.A(n_2690),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2553),
.B(n_848),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2554),
.B(n_2562),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2564),
.B(n_589),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2682),
.Y(n_2898)
);

AND2x4_ASAP7_75t_L g2899 ( 
.A(n_2642),
.B(n_592),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2597),
.B(n_594),
.Y(n_2900)
);

AO21x2_ASAP7_75t_L g2901 ( 
.A1(n_2549),
.A2(n_596),
.B(n_597),
.Y(n_2901)
);

A2O1A1Ixp33_ASAP7_75t_L g2902 ( 
.A1(n_2443),
.A2(n_601),
.B(n_598),
.C(n_600),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2565),
.Y(n_2903)
);

AND2x4_ASAP7_75t_L g2904 ( 
.A(n_2642),
.B(n_602),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2575),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2690),
.B(n_604),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2440),
.B(n_605),
.Y(n_2907)
);

INVx4_ASAP7_75t_L g2908 ( 
.A(n_2512),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2539),
.Y(n_2909)
);

OR2x2_ASAP7_75t_L g2910 ( 
.A(n_2405),
.B(n_606),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2579),
.B(n_847),
.Y(n_2911)
);

HB1xp67_ASAP7_75t_L g2912 ( 
.A(n_2524),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2545),
.Y(n_2913)
);

HB1xp67_ASAP7_75t_L g2914 ( 
.A(n_2512),
.Y(n_2914)
);

BUFx2_ASAP7_75t_L g2915 ( 
.A(n_2517),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2481),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_2916)
);

A2O1A1Ixp33_ASAP7_75t_L g2917 ( 
.A1(n_2448),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2499),
.B(n_611),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2517),
.Y(n_2919)
);

BUFx3_ASAP7_75t_L g2920 ( 
.A(n_2517),
.Y(n_2920)
);

HB1xp67_ASAP7_75t_L g2921 ( 
.A(n_2461),
.Y(n_2921)
);

NAND2x1_ASAP7_75t_L g2922 ( 
.A(n_2447),
.B(n_612),
.Y(n_2922)
);

OAI21x1_ASAP7_75t_SL g2923 ( 
.A1(n_2748),
.A2(n_616),
.B(n_617),
.Y(n_2923)
);

AND2x2_ASAP7_75t_L g2924 ( 
.A(n_2499),
.B(n_2608),
.Y(n_2924)
);

OAI211xp5_ASAP7_75t_L g2925 ( 
.A1(n_2726),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_2925)
);

OAI222xp33_ASAP7_75t_L g2926 ( 
.A1(n_2404),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.C1(n_622),
.C2(n_623),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2625),
.B(n_2598),
.Y(n_2927)
);

AOI22xp33_ASAP7_75t_SL g2928 ( 
.A1(n_2426),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2629),
.B(n_626),
.Y(n_2929)
);

AOI21xp33_ASAP7_75t_SL g2930 ( 
.A1(n_2617),
.A2(n_630),
.B(n_631),
.Y(n_2930)
);

NAND2x1p5_ASAP7_75t_L g2931 ( 
.A(n_2407),
.B(n_631),
.Y(n_2931)
);

INVx6_ASAP7_75t_L g2932 ( 
.A(n_2757),
.Y(n_2932)
);

AND2x4_ASAP7_75t_L g2933 ( 
.A(n_2447),
.B(n_633),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2634),
.B(n_633),
.Y(n_2934)
);

INVx1_ASAP7_75t_SL g2935 ( 
.A(n_2477),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2714),
.B(n_634),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2526),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2696),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2567),
.A2(n_638),
.B(n_639),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2757),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2561),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_SL g2942 ( 
.A1(n_2530),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_2942)
);

OAI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2610),
.A2(n_644),
.B(n_646),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2654),
.B(n_646),
.Y(n_2944)
);

A2O1A1Ixp33_ASAP7_75t_L g2945 ( 
.A1(n_2457),
.A2(n_649),
.B(n_647),
.C(n_648),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2432),
.B(n_2483),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2666),
.B(n_649),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2566),
.A2(n_650),
.B(n_651),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_2418),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2736),
.B(n_654),
.Y(n_2950)
);

CKINVDCx11_ASAP7_75t_R g2951 ( 
.A(n_2582),
.Y(n_2951)
);

NOR2xp33_ASAP7_75t_SL g2952 ( 
.A(n_2669),
.B(n_655),
.Y(n_2952)
);

AO21x2_ASAP7_75t_L g2953 ( 
.A1(n_2574),
.A2(n_656),
.B(n_657),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2469),
.B(n_656),
.Y(n_2954)
);

OAI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2638),
.A2(n_657),
.B(n_658),
.Y(n_2955)
);

AOI221xp5_ASAP7_75t_L g2956 ( 
.A1(n_2425),
.A2(n_659),
.B1(n_660),
.B2(n_661),
.C(n_662),
.Y(n_2956)
);

AO21x1_ASAP7_75t_L g2957 ( 
.A1(n_2422),
.A2(n_660),
.B(n_661),
.Y(n_2957)
);

BUFx6f_ASAP7_75t_L g2958 ( 
.A(n_2539),
.Y(n_2958)
);

BUFx3_ASAP7_75t_L g2959 ( 
.A(n_2719),
.Y(n_2959)
);

A2O1A1Ixp33_ASAP7_75t_L g2960 ( 
.A1(n_2468),
.A2(n_665),
.B(n_663),
.C(n_664),
.Y(n_2960)
);

AOI21x1_ASAP7_75t_L g2961 ( 
.A1(n_2552),
.A2(n_666),
.B(n_667),
.Y(n_2961)
);

OAI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2423),
.A2(n_669),
.B1(n_667),
.B2(n_668),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2525),
.A2(n_670),
.B(n_671),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2434),
.A2(n_672),
.B1(n_670),
.B2(n_671),
.Y(n_2964)
);

AND2x2_ASAP7_75t_SL g2965 ( 
.A(n_2539),
.B(n_673),
.Y(n_2965)
);

BUFx12f_ASAP7_75t_L g2966 ( 
.A(n_2477),
.Y(n_2966)
);

BUFx6f_ASAP7_75t_L g2967 ( 
.A(n_2542),
.Y(n_2967)
);

O2A1O1Ixp33_ASAP7_75t_L g2968 ( 
.A1(n_2444),
.A2(n_677),
.B(n_675),
.C(n_676),
.Y(n_2968)
);

OR2x6_ASAP7_75t_L g2969 ( 
.A(n_2721),
.B(n_675),
.Y(n_2969)
);

AOI21xp33_ASAP7_75t_SL g2970 ( 
.A1(n_2600),
.A2(n_678),
.B(n_679),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_SL g2971 ( 
.A1(n_2749),
.A2(n_680),
.B(n_681),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2409),
.B(n_2442),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2646),
.B(n_682),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2698),
.A2(n_683),
.B1(n_684),
.B2(n_685),
.Y(n_2974)
);

NAND2x1p5_ASAP7_75t_L g2975 ( 
.A(n_2491),
.B(n_846),
.Y(n_2975)
);

OAI21x1_ASAP7_75t_SL g2976 ( 
.A1(n_2749),
.A2(n_684),
.B(n_685),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2491),
.Y(n_2977)
);

NAND2xp33_ASAP7_75t_R g2978 ( 
.A(n_2646),
.B(n_2718),
.Y(n_2978)
);

AOI22x1_ASAP7_75t_L g2979 ( 
.A1(n_2493),
.A2(n_686),
.B1(n_687),
.B2(n_688),
.Y(n_2979)
);

BUFx3_ASAP7_75t_L g2980 ( 
.A(n_2542),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2582),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2445),
.B(n_687),
.Y(n_2982)
);

AO31x2_ASAP7_75t_L g2983 ( 
.A1(n_2416),
.A2(n_688),
.A3(n_689),
.B(n_690),
.Y(n_2983)
);

INVxp67_ASAP7_75t_L g2984 ( 
.A(n_2568),
.Y(n_2984)
);

OA21x2_ASAP7_75t_L g2985 ( 
.A1(n_2658),
.A2(n_691),
.B(n_692),
.Y(n_2985)
);

OR2x6_ASAP7_75t_L g2986 ( 
.A(n_2643),
.B(n_691),
.Y(n_2986)
);

AOI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2612),
.A2(n_692),
.B1(n_693),
.B2(n_694),
.Y(n_2987)
);

AOI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2705),
.A2(n_695),
.B1(n_696),
.B2(n_697),
.Y(n_2988)
);

O2A1O1Ixp33_ASAP7_75t_SL g2989 ( 
.A1(n_2556),
.A2(n_2619),
.B(n_2649),
.C(n_2644),
.Y(n_2989)
);

BUFx2_ASAP7_75t_R g2990 ( 
.A(n_2537),
.Y(n_2990)
);

OAI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2453),
.A2(n_698),
.B(n_699),
.Y(n_2991)
);

BUFx2_ASAP7_75t_L g2992 ( 
.A(n_2542),
.Y(n_2992)
);

AOI21x1_ASAP7_75t_L g2993 ( 
.A1(n_2687),
.A2(n_700),
.B(n_702),
.Y(n_2993)
);

AOI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2664),
.A2(n_703),
.B(n_704),
.Y(n_2994)
);

INVx1_ASAP7_75t_SL g2995 ( 
.A(n_2594),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2408),
.Y(n_2996)
);

NOR2x1_ASAP7_75t_SL g2997 ( 
.A(n_2544),
.B(n_705),
.Y(n_2997)
);

OA21x2_ASAP7_75t_L g2998 ( 
.A1(n_2660),
.A2(n_706),
.B(n_707),
.Y(n_2998)
);

AOI21xp33_ASAP7_75t_L g2999 ( 
.A1(n_2659),
.A2(n_706),
.B(n_707),
.Y(n_2999)
);

INVx3_ASAP7_75t_L g3000 ( 
.A(n_2544),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2415),
.Y(n_3001)
);

NOR2x1_ASAP7_75t_R g3002 ( 
.A(n_2718),
.B(n_708),
.Y(n_3002)
);

AO21x2_ASAP7_75t_L g3003 ( 
.A1(n_2411),
.A2(n_710),
.B(n_711),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2428),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2636),
.A2(n_710),
.B(n_711),
.Y(n_3005)
);

OAI221xp5_ASAP7_75t_L g3006 ( 
.A1(n_2742),
.A2(n_712),
.B1(n_713),
.B2(n_714),
.C(n_715),
.Y(n_3006)
);

NOR2xp33_ASAP7_75t_L g3007 ( 
.A(n_2601),
.B(n_713),
.Y(n_3007)
);

NAND2x1p5_ASAP7_75t_L g3008 ( 
.A(n_2544),
.B(n_2623),
.Y(n_3008)
);

AND2x4_ASAP7_75t_L g3009 ( 
.A(n_2460),
.B(n_2485),
.Y(n_3009)
);

CKINVDCx20_ASAP7_75t_R g3010 ( 
.A(n_2653),
.Y(n_3010)
);

AO31x2_ASAP7_75t_L g3011 ( 
.A1(n_2662),
.A2(n_716),
.A3(n_717),
.B(n_718),
.Y(n_3011)
);

INVx6_ASAP7_75t_L g3012 ( 
.A(n_2653),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2737),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2587),
.Y(n_3014)
);

NAND2x1p5_ASAP7_75t_L g3015 ( 
.A(n_2529),
.B(n_2540),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2488),
.Y(n_3016)
);

AND2x4_ASAP7_75t_L g3017 ( 
.A(n_2490),
.B(n_716),
.Y(n_3017)
);

O2A1O1Ixp33_ASAP7_75t_SL g3018 ( 
.A1(n_2702),
.A2(n_719),
.B(n_720),
.C(n_721),
.Y(n_3018)
);

CKINVDCx20_ASAP7_75t_R g3019 ( 
.A(n_2653),
.Y(n_3019)
);

AND2x4_ASAP7_75t_L g3020 ( 
.A(n_2661),
.B(n_721),
.Y(n_3020)
);

OAI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2472),
.A2(n_722),
.B(n_723),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2734),
.A2(n_724),
.B1(n_725),
.B2(n_726),
.Y(n_3022)
);

INVx8_ASAP7_75t_L g3023 ( 
.A(n_2578),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_SL g3024 ( 
.A(n_2604),
.B(n_2613),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2611),
.A2(n_727),
.B1(n_728),
.B2(n_729),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2578),
.Y(n_3026)
);

BUFx3_ASAP7_75t_L g3027 ( 
.A(n_2684),
.Y(n_3027)
);

INVxp67_ASAP7_75t_L g3028 ( 
.A(n_2616),
.Y(n_3028)
);

OAI21x1_ASAP7_75t_SL g3029 ( 
.A1(n_2667),
.A2(n_2689),
.B(n_2672),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2506),
.A2(n_2632),
.B(n_2620),
.Y(n_3030)
);

AOI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2464),
.A2(n_730),
.B1(n_731),
.B2(n_732),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2668),
.B(n_730),
.Y(n_3032)
);

INVx4_ASAP7_75t_L g3033 ( 
.A(n_2677),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_2587),
.Y(n_3034)
);

BUFx2_ASAP7_75t_L g3035 ( 
.A(n_2684),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2466),
.B(n_733),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2752),
.Y(n_3037)
);

BUFx3_ASAP7_75t_L g3038 ( 
.A(n_2570),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2484),
.Y(n_3039)
);

INVx4_ASAP7_75t_L g3040 ( 
.A(n_2677),
.Y(n_3040)
);

OA21x2_ASAP7_75t_L g3041 ( 
.A1(n_2708),
.A2(n_734),
.B(n_735),
.Y(n_3041)
);

AOI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_2750),
.A2(n_735),
.B1(n_736),
.B2(n_738),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_2473),
.B(n_736),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2602),
.B(n_2433),
.Y(n_3044)
);

NOR2x1_ASAP7_75t_R g3045 ( 
.A(n_2746),
.B(n_738),
.Y(n_3045)
);

INVx1_ASAP7_75t_SL g3046 ( 
.A(n_2710),
.Y(n_3046)
);

AOI221x1_ASAP7_75t_L g3047 ( 
.A1(n_2497),
.A2(n_739),
.B1(n_740),
.B2(n_741),
.C(n_742),
.Y(n_3047)
);

OAI22xp5_ASAP7_75t_L g3048 ( 
.A1(n_2695),
.A2(n_740),
.B1(n_741),
.B2(n_742),
.Y(n_3048)
);

OAI21x1_ASAP7_75t_SL g3049 ( 
.A1(n_2709),
.A2(n_743),
.B(n_744),
.Y(n_3049)
);

INVx1_ASAP7_75t_SL g3050 ( 
.A(n_2707),
.Y(n_3050)
);

BUFx12f_ASAP7_75t_L g3051 ( 
.A(n_2677),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2492),
.Y(n_3052)
);

OAI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2438),
.A2(n_746),
.B(n_748),
.Y(n_3053)
);

AND2x4_ASAP7_75t_L g3054 ( 
.A(n_2670),
.B(n_748),
.Y(n_3054)
);

OA21x2_ASAP7_75t_L g3055 ( 
.A1(n_2716),
.A2(n_749),
.B(n_750),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2492),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2492),
.Y(n_3057)
);

OR2x6_ASAP7_75t_L g3058 ( 
.A(n_2505),
.B(n_2501),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2484),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2433),
.B(n_750),
.Y(n_3060)
);

NOR2x1_ASAP7_75t_SL g3061 ( 
.A(n_2738),
.B(n_751),
.Y(n_3061)
);

AO31x2_ASAP7_75t_L g3062 ( 
.A1(n_2498),
.A2(n_751),
.A3(n_754),
.B(n_755),
.Y(n_3062)
);

INVx1_ASAP7_75t_SL g3063 ( 
.A(n_2739),
.Y(n_3063)
);

AND2x4_ASAP7_75t_L g3064 ( 
.A(n_2648),
.B(n_757),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2433),
.B(n_758),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2751),
.B(n_2615),
.Y(n_3066)
);

AOI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_2683),
.A2(n_760),
.B1(n_761),
.B2(n_762),
.Y(n_3067)
);

AOI22xp33_ASAP7_75t_L g3068 ( 
.A1(n_2758),
.A2(n_762),
.B1(n_764),
.B2(n_765),
.Y(n_3068)
);

BUFx6f_ASAP7_75t_SL g3069 ( 
.A(n_2570),
.Y(n_3069)
);

AOI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2656),
.A2(n_766),
.B(n_768),
.Y(n_3070)
);

O2A1O1Ixp33_ASAP7_75t_SL g3071 ( 
.A1(n_2723),
.A2(n_768),
.B(n_769),
.C(n_770),
.Y(n_3071)
);

AOI22xp5_ASAP7_75t_L g3072 ( 
.A1(n_2686),
.A2(n_769),
.B1(n_770),
.B2(n_771),
.Y(n_3072)
);

CKINVDCx6p67_ASAP7_75t_R g3073 ( 
.A(n_2675),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2854),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2779),
.Y(n_3075)
);

NAND2xp33_ASAP7_75t_SL g3076 ( 
.A(n_2787),
.B(n_2606),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2903),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_3058),
.A2(n_2430),
.B1(n_2680),
.B2(n_2558),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2905),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2802),
.Y(n_3080)
);

OAI221xp5_ASAP7_75t_L g3081 ( 
.A1(n_2952),
.A2(n_2509),
.B1(n_2633),
.B2(n_2528),
.C(n_2538),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_3052),
.B(n_2673),
.Y(n_3082)
);

CKINVDCx11_ASAP7_75t_R g3083 ( 
.A(n_2759),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2927),
.B(n_2773),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2819),
.Y(n_3085)
);

OR2x6_ASAP7_75t_L g3086 ( 
.A(n_2885),
.B(n_2505),
.Y(n_3086)
);

BUFx3_ASAP7_75t_L g3087 ( 
.A(n_2940),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2828),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2875),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2913),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2996),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_3001),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2890),
.Y(n_3093)
);

AOI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2978),
.A2(n_2787),
.B1(n_2894),
.B2(n_2965),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2896),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_3004),
.Y(n_3096)
);

BUFx3_ASAP7_75t_L g3097 ( 
.A(n_2932),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_3016),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2760),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2760),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2775),
.B(n_2560),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_2763),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2907),
.B(n_2560),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2973),
.B(n_2560),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2763),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2766),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2880),
.Y(n_3107)
);

HB1xp67_ASAP7_75t_L g3108 ( 
.A(n_2766),
.Y(n_3108)
);

AO21x1_ASAP7_75t_L g3109 ( 
.A1(n_2930),
.A2(n_2482),
.B(n_2507),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2785),
.B(n_2520),
.Y(n_3110)
);

BUFx4f_ASAP7_75t_SL g3111 ( 
.A(n_2783),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_2860),
.B(n_2573),
.Y(n_3112)
);

HB1xp67_ASAP7_75t_L g3113 ( 
.A(n_2767),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_3058),
.A2(n_2475),
.B1(n_2487),
.B2(n_2480),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2767),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2790),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2790),
.Y(n_3117)
);

INVx3_ASAP7_75t_L g3118 ( 
.A(n_2827),
.Y(n_3118)
);

OAI22xp5_ASAP7_75t_L g3119 ( 
.A1(n_2762),
.A2(n_2450),
.B1(n_2489),
.B2(n_2735),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_3017),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3017),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_2770),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3035),
.Y(n_3123)
);

INVx3_ASAP7_75t_L g3124 ( 
.A(n_2827),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3020),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_3020),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3032),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3032),
.Y(n_3128)
);

INVx3_ASAP7_75t_L g3129 ( 
.A(n_2812),
.Y(n_3129)
);

INVxp33_ASAP7_75t_L g3130 ( 
.A(n_3002),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2812),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3054),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2818),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3054),
.Y(n_3134)
);

BUFx2_ASAP7_75t_L g3135 ( 
.A(n_3010),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2893),
.B(n_2587),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3064),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3064),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2933),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2831),
.B(n_2573),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2933),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2868),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2906),
.B(n_2573),
.Y(n_3143)
);

OAI22xp33_ASAP7_75t_SL g3144 ( 
.A1(n_2886),
.A2(n_2609),
.B1(n_2756),
.B2(n_2740),
.Y(n_3144)
);

AOI21xp33_ASAP7_75t_L g3145 ( 
.A1(n_3029),
.A2(n_2968),
.B(n_2925),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_3050),
.B(n_772),
.Y(n_3146)
);

BUFx2_ASAP7_75t_L g3147 ( 
.A(n_3019),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2872),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_2893),
.B(n_2576),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2895),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2897),
.Y(n_3151)
);

OR2x2_ASAP7_75t_L g3152 ( 
.A(n_2838),
.B(n_2531),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2911),
.Y(n_3153)
);

NAND2x1_ASAP7_75t_L g3154 ( 
.A(n_2971),
.B(n_2592),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2919),
.B(n_2570),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3062),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2918),
.B(n_773),
.Y(n_3157)
);

OAI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_2886),
.A2(n_2729),
.B1(n_2731),
.B2(n_2745),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_3073),
.A2(n_2724),
.B1(n_2621),
.B2(n_2745),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3062),
.Y(n_3160)
);

INVx3_ASAP7_75t_L g3161 ( 
.A(n_2818),
.Y(n_3161)
);

HB1xp67_ASAP7_75t_L g3162 ( 
.A(n_3052),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_2784),
.B(n_2584),
.Y(n_3163)
);

BUFx6f_ASAP7_75t_L g3164 ( 
.A(n_2966),
.Y(n_3164)
);

BUFx2_ASAP7_75t_L g3165 ( 
.A(n_3051),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3062),
.Y(n_3166)
);

NAND2x1p5_ASAP7_75t_L g3167 ( 
.A(n_2830),
.B(n_2592),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_2776),
.Y(n_3168)
);

INVx3_ASAP7_75t_L g3169 ( 
.A(n_2830),
.Y(n_3169)
);

BUFx4f_ASAP7_75t_SL g3170 ( 
.A(n_2807),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2873),
.Y(n_3171)
);

AND2x4_ASAP7_75t_SL g3172 ( 
.A(n_2888),
.B(n_2692),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2873),
.Y(n_3173)
);

BUFx12f_ASAP7_75t_L g3174 ( 
.A(n_2932),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_2929),
.B(n_773),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2873),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2861),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_2844),
.Y(n_3178)
);

BUFx6f_ASAP7_75t_L g3179 ( 
.A(n_2776),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2861),
.Y(n_3180)
);

OAI221xp5_ASAP7_75t_L g3181 ( 
.A1(n_2811),
.A2(n_2722),
.B1(n_2674),
.B2(n_2678),
.C(n_2641),
.Y(n_3181)
);

OR2x2_ASAP7_75t_L g3182 ( 
.A(n_2883),
.B(n_2585),
.Y(n_3182)
);

BUFx2_ASAP7_75t_L g3183 ( 
.A(n_2848),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2861),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3027),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2934),
.B(n_774),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3066),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2949),
.Y(n_3188)
);

INVxp67_ASAP7_75t_L g3189 ( 
.A(n_3013),
.Y(n_3189)
);

BUFx3_ASAP7_75t_L g3190 ( 
.A(n_2959),
.Y(n_3190)
);

INVx3_ASAP7_75t_L g3191 ( 
.A(n_2844),
.Y(n_3191)
);

HB1xp67_ASAP7_75t_L g3192 ( 
.A(n_3056),
.Y(n_3192)
);

OR2x2_ASAP7_75t_L g3193 ( 
.A(n_2912),
.B(n_2494),
.Y(n_3193)
);

HB1xp67_ASAP7_75t_L g3194 ( 
.A(n_3056),
.Y(n_3194)
);

INVx3_ASAP7_75t_L g3195 ( 
.A(n_2908),
.Y(n_3195)
);

BUFx2_ASAP7_75t_L g3196 ( 
.A(n_2980),
.Y(n_3196)
);

OR2x6_ASAP7_75t_L g3197 ( 
.A(n_2888),
.B(n_2508),
.Y(n_3197)
);

HB1xp67_ASAP7_75t_L g3198 ( 
.A(n_3057),
.Y(n_3198)
);

CKINVDCx12_ASAP7_75t_R g3199 ( 
.A(n_3045),
.Y(n_3199)
);

HB1xp67_ASAP7_75t_L g3200 ( 
.A(n_3057),
.Y(n_3200)
);

OR2x2_ASAP7_75t_L g3201 ( 
.A(n_3026),
.B(n_2502),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_2969),
.A2(n_2521),
.B1(n_2557),
.B2(n_2577),
.Y(n_3202)
);

AOI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_2969),
.A2(n_2532),
.B1(n_2548),
.B2(n_2541),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3044),
.Y(n_3204)
);

AOI22xp33_ASAP7_75t_L g3205 ( 
.A1(n_2800),
.A2(n_2534),
.B1(n_2536),
.B2(n_2571),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_2944),
.B(n_774),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2924),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2947),
.B(n_775),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2822),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2768),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2983),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_2921),
.B(n_2743),
.Y(n_3212)
);

BUFx12f_ASAP7_75t_L g3213 ( 
.A(n_2846),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2983),
.Y(n_3214)
);

INVx3_ASAP7_75t_L g3215 ( 
.A(n_2908),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2983),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3037),
.Y(n_3217)
);

INVx1_ASAP7_75t_SL g3218 ( 
.A(n_2935),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_SL g3219 ( 
.A(n_2899),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2817),
.B(n_776),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_2920),
.B(n_2639),
.Y(n_3221)
);

BUFx3_ASAP7_75t_L g3222 ( 
.A(n_2951),
.Y(n_3222)
);

INVx3_ASAP7_75t_L g3223 ( 
.A(n_3033),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_2984),
.B(n_777),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_3028),
.B(n_2647),
.Y(n_3225)
);

INVx3_ASAP7_75t_L g3226 ( 
.A(n_3033),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2803),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2829),
.Y(n_3228)
);

INVx1_ASAP7_75t_SL g3229 ( 
.A(n_2992),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2829),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2835),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_2954),
.B(n_777),
.Y(n_3232)
);

INVx3_ASAP7_75t_L g3233 ( 
.A(n_3040),
.Y(n_3233)
);

BUFx3_ASAP7_75t_L g3234 ( 
.A(n_2792),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2836),
.Y(n_3235)
);

HB1xp67_ASAP7_75t_SL g3236 ( 
.A(n_2899),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2836),
.Y(n_3237)
);

AND2x2_ASAP7_75t_L g3238 ( 
.A(n_2900),
.B(n_778),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2840),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2799),
.B(n_2754),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2843),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2843),
.B(n_2853),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_2804),
.B(n_778),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2853),
.Y(n_3244)
);

BUFx2_ASAP7_75t_L g3245 ( 
.A(n_3023),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2862),
.Y(n_3246)
);

HB1xp67_ASAP7_75t_L g3247 ( 
.A(n_2862),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2863),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2863),
.Y(n_3249)
);

BUFx2_ASAP7_75t_L g3250 ( 
.A(n_3023),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_2777),
.B(n_779),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2889),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2898),
.B(n_2693),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2898),
.B(n_2693),
.Y(n_3254)
);

BUFx6f_ASAP7_75t_L g3255 ( 
.A(n_2776),
.Y(n_3255)
);

OR2x2_ASAP7_75t_L g3256 ( 
.A(n_2867),
.B(n_2596),
.Y(n_3256)
);

A2O1A1Ixp33_ASAP7_75t_L g3257 ( 
.A1(n_2837),
.A2(n_2627),
.B(n_2645),
.C(n_2618),
.Y(n_3257)
);

INVx1_ASAP7_75t_SL g3258 ( 
.A(n_3012),
.Y(n_3258)
);

AND2x4_ASAP7_75t_L g3259 ( 
.A(n_2909),
.B(n_2693),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_2823),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_2794),
.B(n_779),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_SL g3262 ( 
.A(n_2990),
.B(n_2720),
.Y(n_3262)
);

INVx3_ASAP7_75t_L g3263 ( 
.A(n_3040),
.Y(n_3263)
);

HB1xp67_ASAP7_75t_L g3264 ( 
.A(n_2938),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2833),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_2977),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3060),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3065),
.Y(n_3268)
);

BUFx2_ASAP7_75t_L g3269 ( 
.A(n_3038),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3011),
.Y(n_3270)
);

INVxp67_ASAP7_75t_L g3271 ( 
.A(n_3059),
.Y(n_3271)
);

INVx3_ASAP7_75t_L g3272 ( 
.A(n_3008),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3011),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3011),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2975),
.Y(n_3275)
);

AOI221xp5_ASAP7_75t_L g3276 ( 
.A1(n_2946),
.A2(n_2605),
.B1(n_2607),
.B2(n_2727),
.C(n_2711),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2995),
.B(n_781),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2769),
.Y(n_3278)
);

BUFx6f_ASAP7_75t_L g3279 ( 
.A(n_2823),
.Y(n_3279)
);

OR2x6_ASAP7_75t_L g3280 ( 
.A(n_2931),
.B(n_2580),
.Y(n_3280)
);

INVx2_ASAP7_75t_SL g3281 ( 
.A(n_3012),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_3046),
.B(n_781),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_2904),
.B(n_782),
.Y(n_3283)
);

OR2x2_ASAP7_75t_L g3284 ( 
.A(n_2972),
.B(n_2713),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2806),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_2800),
.A2(n_2663),
.B1(n_2655),
.B2(n_2651),
.Y(n_3286)
);

OR2x2_ASAP7_75t_L g3287 ( 
.A(n_2857),
.B(n_2701),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2815),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_2904),
.B(n_782),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2815),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2815),
.Y(n_3291)
);

INVx4_ASAP7_75t_L g3292 ( 
.A(n_2958),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3059),
.B(n_2715),
.Y(n_3293)
);

NAND2xp33_ASAP7_75t_L g3294 ( 
.A(n_2981),
.B(n_783),
.Y(n_3294)
);

INVx3_ASAP7_75t_L g3295 ( 
.A(n_2823),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_3006),
.A2(n_785),
.B1(n_786),
.B2(n_787),
.Y(n_3296)
);

INVx3_ASAP7_75t_L g3297 ( 
.A(n_2826),
.Y(n_3297)
);

HB1xp67_ASAP7_75t_L g3298 ( 
.A(n_3039),
.Y(n_3298)
);

AOI22xp33_ASAP7_75t_L g3299 ( 
.A1(n_2774),
.A2(n_785),
.B1(n_787),
.B2(n_789),
.Y(n_3299)
);

AO21x2_ASAP7_75t_L g3300 ( 
.A1(n_3030),
.A2(n_789),
.B(n_790),
.Y(n_3300)
);

OR2x2_ASAP7_75t_L g3301 ( 
.A(n_3043),
.B(n_791),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2814),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2814),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2814),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2879),
.Y(n_3305)
);

BUFx3_ASAP7_75t_L g3306 ( 
.A(n_2871),
.Y(n_3306)
);

OR2x2_ASAP7_75t_L g3307 ( 
.A(n_2910),
.B(n_792),
.Y(n_3307)
);

HB1xp67_ASAP7_75t_L g3308 ( 
.A(n_2914),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_3063),
.B(n_846),
.Y(n_3309)
);

CKINVDCx5p33_ASAP7_75t_R g3310 ( 
.A(n_2842),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_SL g3311 ( 
.A(n_3024),
.B(n_792),
.Y(n_3311)
);

AND2x4_ASAP7_75t_L g3312 ( 
.A(n_3245),
.B(n_3250),
.Y(n_3312)
);

NAND2xp33_ASAP7_75t_R g3313 ( 
.A(n_3165),
.B(n_2936),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3187),
.B(n_3009),
.Y(n_3314)
);

INVxp67_ASAP7_75t_L g3315 ( 
.A(n_3219),
.Y(n_3315)
);

NAND2xp33_ASAP7_75t_R g3316 ( 
.A(n_3133),
.B(n_2851),
.Y(n_3316)
);

AND2x4_ASAP7_75t_L g3317 ( 
.A(n_3269),
.B(n_2891),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_R g3318 ( 
.A(n_3219),
.B(n_3236),
.Y(n_3318)
);

AND2x4_ASAP7_75t_L g3319 ( 
.A(n_3196),
.B(n_2915),
.Y(n_3319)
);

CKINVDCx14_ASAP7_75t_R g3320 ( 
.A(n_3083),
.Y(n_3320)
);

XNOR2xp5_ASAP7_75t_L g3321 ( 
.A(n_3122),
.B(n_2855),
.Y(n_3321)
);

XNOR2xp5_ASAP7_75t_L g3322 ( 
.A(n_3310),
.B(n_2859),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_R g3323 ( 
.A(n_3236),
.B(n_2878),
.Y(n_3323)
);

CKINVDCx5p33_ASAP7_75t_R g3324 ( 
.A(n_3174),
.Y(n_3324)
);

NAND2xp33_ASAP7_75t_R g3325 ( 
.A(n_3133),
.B(n_2858),
.Y(n_3325)
);

BUFx10_ASAP7_75t_L g3326 ( 
.A(n_3164),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3089),
.B(n_3009),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_3190),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3074),
.Y(n_3329)
);

INVxp67_ASAP7_75t_L g3330 ( 
.A(n_3218),
.Y(n_3330)
);

XNOR2xp5_ASAP7_75t_L g3331 ( 
.A(n_3234),
.B(n_2928),
.Y(n_3331)
);

CKINVDCx5p33_ASAP7_75t_R g3332 ( 
.A(n_3213),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3077),
.Y(n_3333)
);

NAND2xp33_ASAP7_75t_R g3334 ( 
.A(n_3161),
.B(n_2986),
.Y(n_3334)
);

XOR2xp5_ASAP7_75t_L g3335 ( 
.A(n_3222),
.B(n_3015),
.Y(n_3335)
);

NOR2xp33_ASAP7_75t_R g3336 ( 
.A(n_3111),
.B(n_2865),
.Y(n_3336)
);

BUFx6f_ASAP7_75t_L g3337 ( 
.A(n_3087),
.Y(n_3337)
);

AND2x4_ASAP7_75t_L g3338 ( 
.A(n_3161),
.B(n_3000),
.Y(n_3338)
);

NAND2xp33_ASAP7_75t_R g3339 ( 
.A(n_3283),
.B(n_2986),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_R g3340 ( 
.A(n_3111),
.B(n_2961),
.Y(n_3340)
);

NAND2x1_ASAP7_75t_L g3341 ( 
.A(n_3086),
.B(n_2976),
.Y(n_3341)
);

BUFx3_ASAP7_75t_L g3342 ( 
.A(n_3097),
.Y(n_3342)
);

AND2x4_ASAP7_75t_L g3343 ( 
.A(n_3094),
.B(n_3000),
.Y(n_3343)
);

AND2x4_ASAP7_75t_L g3344 ( 
.A(n_3094),
.B(n_2958),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3093),
.B(n_3007),
.Y(n_3345)
);

AND2x4_ASAP7_75t_L g3346 ( 
.A(n_3195),
.B(n_3215),
.Y(n_3346)
);

AND2x4_ASAP7_75t_L g3347 ( 
.A(n_3195),
.B(n_2958),
.Y(n_3347)
);

OR2x4_ASAP7_75t_L g3348 ( 
.A(n_3164),
.B(n_2809),
.Y(n_3348)
);

INVx8_ASAP7_75t_L g3349 ( 
.A(n_3164),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3130),
.B(n_2782),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_3084),
.B(n_3003),
.Y(n_3351)
);

NAND2xp33_ASAP7_75t_R g3352 ( 
.A(n_3289),
.B(n_2761),
.Y(n_3352)
);

OR2x6_ASAP7_75t_L g3353 ( 
.A(n_3183),
.B(n_2771),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_L g3354 ( 
.A(n_3135),
.B(n_2982),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3075),
.Y(n_3355)
);

INVxp67_ASAP7_75t_L g3356 ( 
.A(n_3218),
.Y(n_3356)
);

BUFx24_ASAP7_75t_SL g3357 ( 
.A(n_3202),
.Y(n_3357)
);

BUFx3_ASAP7_75t_L g3358 ( 
.A(n_3170),
.Y(n_3358)
);

NAND2xp33_ASAP7_75t_R g3359 ( 
.A(n_3169),
.B(n_2761),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3207),
.B(n_3014),
.Y(n_3360)
);

NAND2xp33_ASAP7_75t_R g3361 ( 
.A(n_3169),
.B(n_2970),
.Y(n_3361)
);

NAND2xp33_ASAP7_75t_R g3362 ( 
.A(n_3178),
.B(n_2985),
.Y(n_3362)
);

NAND2xp33_ASAP7_75t_R g3363 ( 
.A(n_3178),
.B(n_2985),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_3076),
.B(n_2957),
.Y(n_3364)
);

CKINVDCx5p33_ASAP7_75t_R g3365 ( 
.A(n_3170),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3107),
.B(n_3014),
.Y(n_3366)
);

NAND2xp33_ASAP7_75t_R g3367 ( 
.A(n_3191),
.B(n_2998),
.Y(n_3367)
);

BUFx3_ASAP7_75t_L g3368 ( 
.A(n_3147),
.Y(n_3368)
);

BUFx3_ASAP7_75t_L g3369 ( 
.A(n_3306),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_R g3370 ( 
.A(n_3199),
.B(n_2993),
.Y(n_3370)
);

BUFx24_ASAP7_75t_SL g3371 ( 
.A(n_3202),
.Y(n_3371)
);

NAND2xp33_ASAP7_75t_R g3372 ( 
.A(n_3191),
.B(n_3223),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3095),
.B(n_2916),
.Y(n_3373)
);

BUFx10_ASAP7_75t_L g3374 ( 
.A(n_3172),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_3225),
.B(n_3036),
.Y(n_3375)
);

NAND2xp33_ASAP7_75t_R g3376 ( 
.A(n_3223),
.B(n_2998),
.Y(n_3376)
);

XNOR2xp5_ASAP7_75t_L g3377 ( 
.A(n_3251),
.B(n_2789),
.Y(n_3377)
);

INVxp67_ASAP7_75t_L g3378 ( 
.A(n_3225),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3188),
.B(n_3034),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_3266),
.Y(n_3380)
);

NAND2xp33_ASAP7_75t_R g3381 ( 
.A(n_3226),
.B(n_3233),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_3226),
.Y(n_3382)
);

AND2x4_ASAP7_75t_L g3383 ( 
.A(n_3215),
.B(n_2967),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3079),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_R g3385 ( 
.A(n_3294),
.B(n_3069),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3233),
.B(n_3263),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_3266),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_R g3388 ( 
.A(n_3262),
.B(n_3069),
.Y(n_3388)
);

INVxp67_ASAP7_75t_L g3389 ( 
.A(n_3308),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_R g3390 ( 
.A(n_3262),
.B(n_2874),
.Y(n_3390)
);

NAND2xp33_ASAP7_75t_R g3391 ( 
.A(n_3263),
.B(n_3041),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3159),
.B(n_3034),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3091),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_R g3394 ( 
.A(n_3129),
.B(n_2881),
.Y(n_3394)
);

INVxp67_ASAP7_75t_L g3395 ( 
.A(n_3308),
.Y(n_3395)
);

OR2x6_ASAP7_75t_L g3396 ( 
.A(n_3311),
.B(n_2922),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3204),
.B(n_2967),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3143),
.B(n_2967),
.Y(n_3398)
);

BUFx6f_ASAP7_75t_L g3399 ( 
.A(n_3168),
.Y(n_3399)
);

NAND2xp33_ASAP7_75t_R g3400 ( 
.A(n_3086),
.B(n_3041),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_3281),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3278),
.B(n_3053),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3092),
.Y(n_3403)
);

CKINVDCx20_ASAP7_75t_R g3404 ( 
.A(n_3220),
.Y(n_3404)
);

NAND2xp33_ASAP7_75t_R g3405 ( 
.A(n_3086),
.B(n_3055),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_R g3406 ( 
.A(n_3131),
.B(n_3055),
.Y(n_3406)
);

BUFx3_ASAP7_75t_L g3407 ( 
.A(n_3155),
.Y(n_3407)
);

OR2x6_ASAP7_75t_L g3408 ( 
.A(n_3311),
.B(n_2780),
.Y(n_3408)
);

INVxp67_ASAP7_75t_L g3409 ( 
.A(n_3224),
.Y(n_3409)
);

OR2x6_ASAP7_75t_L g3410 ( 
.A(n_3280),
.B(n_2866),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_R g3411 ( 
.A(n_3118),
.B(n_2884),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_R g3412 ( 
.A(n_3118),
.B(n_793),
.Y(n_3412)
);

CKINVDCx11_ASAP7_75t_R g3413 ( 
.A(n_3258),
.Y(n_3413)
);

AND2x4_ASAP7_75t_L g3414 ( 
.A(n_3229),
.B(n_2997),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_SL g3415 ( 
.A(n_3159),
.B(n_2942),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_R g3416 ( 
.A(n_3124),
.B(n_793),
.Y(n_3416)
);

CKINVDCx12_ASAP7_75t_R g3417 ( 
.A(n_3256),
.Y(n_3417)
);

OR2x6_ASAP7_75t_L g3418 ( 
.A(n_3280),
.B(n_2834),
.Y(n_3418)
);

NAND2xp33_ASAP7_75t_R g3419 ( 
.A(n_3103),
.B(n_794),
.Y(n_3419)
);

INVxp67_ASAP7_75t_L g3420 ( 
.A(n_3175),
.Y(n_3420)
);

INVx8_ASAP7_75t_L g3421 ( 
.A(n_3155),
.Y(n_3421)
);

AND2x4_ASAP7_75t_L g3422 ( 
.A(n_3229),
.B(n_2997),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_3292),
.Y(n_3423)
);

OR2x6_ASAP7_75t_L g3424 ( 
.A(n_3280),
.B(n_2923),
.Y(n_3424)
);

NAND2xp33_ASAP7_75t_R g3425 ( 
.A(n_3124),
.B(n_3238),
.Y(n_3425)
);

BUFx3_ASAP7_75t_L g3426 ( 
.A(n_3292),
.Y(n_3426)
);

INVxp67_ASAP7_75t_L g3427 ( 
.A(n_3186),
.Y(n_3427)
);

NAND2xp33_ASAP7_75t_R g3428 ( 
.A(n_3206),
.B(n_794),
.Y(n_3428)
);

BUFx10_ASAP7_75t_L g3429 ( 
.A(n_3275),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_R g3430 ( 
.A(n_3272),
.B(n_795),
.Y(n_3430)
);

INVxp67_ASAP7_75t_L g3431 ( 
.A(n_3208),
.Y(n_3431)
);

NAND2xp33_ASAP7_75t_SL g3432 ( 
.A(n_3114),
.B(n_2856),
.Y(n_3432)
);

NAND2xp33_ASAP7_75t_R g3433 ( 
.A(n_3232),
.B(n_3272),
.Y(n_3433)
);

XNOR2xp5_ASAP7_75t_L g3434 ( 
.A(n_3157),
.B(n_3243),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_R g3435 ( 
.A(n_3299),
.B(n_796),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3285),
.B(n_2772),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_R g3437 ( 
.A(n_3299),
.B(n_796),
.Y(n_3437)
);

XNOR2xp5_ASAP7_75t_L g3438 ( 
.A(n_3261),
.B(n_2789),
.Y(n_3438)
);

NAND2xp33_ASAP7_75t_SL g3439 ( 
.A(n_3114),
.B(n_2824),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_R g3440 ( 
.A(n_3295),
.B(n_797),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_R g3441 ( 
.A(n_3295),
.B(n_3297),
.Y(n_3441)
);

NAND2xp33_ASAP7_75t_R g3442 ( 
.A(n_3277),
.B(n_798),
.Y(n_3442)
);

AND2x4_ASAP7_75t_L g3443 ( 
.A(n_3137),
.B(n_2801),
.Y(n_3443)
);

NAND2xp33_ASAP7_75t_SL g3444 ( 
.A(n_3152),
.B(n_2901),
.Y(n_3444)
);

AND2x4_ASAP7_75t_L g3445 ( 
.A(n_3138),
.B(n_3061),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3301),
.B(n_2821),
.Y(n_3446)
);

AND2x4_ASAP7_75t_L g3447 ( 
.A(n_3185),
.B(n_3061),
.Y(n_3447)
);

AND2x4_ASAP7_75t_L g3448 ( 
.A(n_3120),
.B(n_2788),
.Y(n_3448)
);

XNOR2xp5_ASAP7_75t_L g3449 ( 
.A(n_3282),
.B(n_3031),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3210),
.B(n_2772),
.Y(n_3450)
);

INVx1_ASAP7_75t_SL g3451 ( 
.A(n_3258),
.Y(n_3451)
);

XOR2xp5_ASAP7_75t_L g3452 ( 
.A(n_3307),
.B(n_2987),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3102),
.Y(n_3453)
);

NAND2xp33_ASAP7_75t_R g3454 ( 
.A(n_3140),
.B(n_798),
.Y(n_3454)
);

AND2x4_ASAP7_75t_L g3455 ( 
.A(n_3121),
.B(n_2791),
.Y(n_3455)
);

CKINVDCx20_ASAP7_75t_R g3456 ( 
.A(n_3309),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3080),
.B(n_2772),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3102),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_R g3459 ( 
.A(n_3297),
.B(n_801),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3108),
.Y(n_3460)
);

NAND2xp33_ASAP7_75t_R g3461 ( 
.A(n_3197),
.B(n_801),
.Y(n_3461)
);

CKINVDCx12_ASAP7_75t_R g3462 ( 
.A(n_3197),
.Y(n_3462)
);

AND2x4_ASAP7_75t_L g3463 ( 
.A(n_3139),
.B(n_2795),
.Y(n_3463)
);

NAND2xp33_ASAP7_75t_R g3464 ( 
.A(n_3197),
.B(n_802),
.Y(n_3464)
);

AND2x4_ASAP7_75t_L g3465 ( 
.A(n_3141),
.B(n_2796),
.Y(n_3465)
);

AND2x4_ASAP7_75t_L g3466 ( 
.A(n_3085),
.B(n_2797),
.Y(n_3466)
);

AND2x4_ASAP7_75t_L g3467 ( 
.A(n_3088),
.B(n_2798),
.Y(n_3467)
);

BUFx10_ASAP7_75t_L g3468 ( 
.A(n_3305),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3112),
.B(n_3072),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3101),
.B(n_2953),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3108),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_R g3472 ( 
.A(n_3168),
.B(n_802),
.Y(n_3472)
);

NAND2xp33_ASAP7_75t_R g3473 ( 
.A(n_3146),
.B(n_803),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3113),
.Y(n_3474)
);

AND2x4_ASAP7_75t_L g3475 ( 
.A(n_3123),
.B(n_2810),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3267),
.B(n_3025),
.Y(n_3476)
);

NAND2xp33_ASAP7_75t_R g3477 ( 
.A(n_3110),
.B(n_804),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3096),
.B(n_2813),
.Y(n_3478)
);

NAND2xp33_ASAP7_75t_R g3479 ( 
.A(n_3110),
.B(n_805),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_3179),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3268),
.B(n_2852),
.Y(n_3481)
);

XOR2xp5_ASAP7_75t_L g3482 ( 
.A(n_3163),
.B(n_2825),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3098),
.B(n_2847),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3104),
.B(n_2847),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3090),
.B(n_2816),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3148),
.B(n_2839),
.Y(n_3486)
);

NOR2xp33_ASAP7_75t_R g3487 ( 
.A(n_3179),
.B(n_806),
.Y(n_3487)
);

NOR2xp33_ASAP7_75t_R g3488 ( 
.A(n_3255),
.B(n_807),
.Y(n_3488)
);

NAND2xp33_ASAP7_75t_R g3489 ( 
.A(n_3287),
.B(n_807),
.Y(n_3489)
);

OR2x4_ASAP7_75t_L g3490 ( 
.A(n_3240),
.B(n_2926),
.Y(n_3490)
);

HB1xp67_ASAP7_75t_L g3491 ( 
.A(n_3212),
.Y(n_3491)
);

AND2x4_ASAP7_75t_L g3492 ( 
.A(n_3136),
.B(n_3047),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3150),
.B(n_2956),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3151),
.B(n_2850),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3113),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3144),
.B(n_2887),
.Y(n_3496)
);

INVxp67_ASAP7_75t_L g3497 ( 
.A(n_3142),
.Y(n_3497)
);

NOR2xp33_ASAP7_75t_R g3498 ( 
.A(n_3260),
.B(n_808),
.Y(n_3498)
);

NAND2xp33_ASAP7_75t_SL g3499 ( 
.A(n_3119),
.B(n_2950),
.Y(n_3499)
);

XOR2xp5_ASAP7_75t_L g3500 ( 
.A(n_3284),
.B(n_2786),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3099),
.Y(n_3501)
);

INVxp67_ASAP7_75t_L g3502 ( 
.A(n_3153),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3116),
.B(n_2876),
.Y(n_3503)
);

XOR2xp5_ASAP7_75t_L g3504 ( 
.A(n_3119),
.B(n_2793),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3209),
.B(n_2877),
.Y(n_3505)
);

INVxp67_ASAP7_75t_L g3506 ( 
.A(n_3182),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3125),
.B(n_3005),
.Y(n_3507)
);

OR2x6_ASAP7_75t_L g3508 ( 
.A(n_3136),
.B(n_2991),
.Y(n_3508)
);

XNOR2xp5_ASAP7_75t_L g3509 ( 
.A(n_3203),
.B(n_2808),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_R g3510 ( 
.A(n_3260),
.B(n_809),
.Y(n_3510)
);

OR2x2_ASAP7_75t_L g3511 ( 
.A(n_3293),
.B(n_2941),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_R g3512 ( 
.A(n_3260),
.B(n_809),
.Y(n_3512)
);

NAND2xp33_ASAP7_75t_R g3513 ( 
.A(n_3240),
.B(n_810),
.Y(n_3513)
);

XNOR2xp5_ASAP7_75t_L g3514 ( 
.A(n_3203),
.B(n_2962),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3100),
.B(n_3021),
.Y(n_3515)
);

NAND2xp33_ASAP7_75t_R g3516 ( 
.A(n_3201),
.B(n_810),
.Y(n_3516)
);

NOR2xp33_ASAP7_75t_L g3517 ( 
.A(n_3193),
.B(n_811),
.Y(n_3517)
);

NAND2xp33_ASAP7_75t_R g3518 ( 
.A(n_3288),
.B(n_811),
.Y(n_3518)
);

CKINVDCx9p33_ASAP7_75t_R g3519 ( 
.A(n_3253),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3105),
.B(n_2964),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_SL g3521 ( 
.A(n_3144),
.B(n_2882),
.Y(n_3521)
);

AND2x4_ASAP7_75t_L g3522 ( 
.A(n_3126),
.B(n_2764),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_R g3523 ( 
.A(n_3279),
.B(n_812),
.Y(n_3523)
);

OR2x6_ASAP7_75t_L g3524 ( 
.A(n_3167),
.B(n_2849),
.Y(n_3524)
);

OR2x6_ASAP7_75t_L g3525 ( 
.A(n_3167),
.B(n_2820),
.Y(n_3525)
);

NAND2xp33_ASAP7_75t_R g3526 ( 
.A(n_3290),
.B(n_812),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_3279),
.Y(n_3527)
);

NAND2xp33_ASAP7_75t_R g3528 ( 
.A(n_3291),
.B(n_813),
.Y(n_3528)
);

AND2x4_ASAP7_75t_L g3529 ( 
.A(n_3127),
.B(n_3128),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_3132),
.B(n_2781),
.Y(n_3530)
);

INVxp67_ASAP7_75t_L g3531 ( 
.A(n_3293),
.Y(n_3531)
);

AND2x4_ASAP7_75t_L g3532 ( 
.A(n_3134),
.B(n_2778),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_3109),
.B(n_2955),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3531),
.B(n_3217),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3380),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3355),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3393),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3453),
.B(n_3227),
.Y(n_3538)
);

HB1xp67_ASAP7_75t_L g3539 ( 
.A(n_3387),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3329),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3491),
.B(n_3106),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3458),
.B(n_3228),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3403),
.Y(n_3543)
);

INVxp67_ASAP7_75t_L g3544 ( 
.A(n_3381),
.Y(n_3544)
);

NAND2x1p5_ASAP7_75t_L g3545 ( 
.A(n_3382),
.B(n_3149),
.Y(n_3545)
);

BUFx2_ASAP7_75t_L g3546 ( 
.A(n_3318),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3333),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3499),
.A2(n_3081),
.B1(n_3078),
.B2(n_3181),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3501),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_3389),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3398),
.B(n_3115),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3460),
.B(n_3471),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3474),
.Y(n_3553)
);

BUFx2_ASAP7_75t_L g3554 ( 
.A(n_3423),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3495),
.Y(n_3555)
);

OR2x2_ASAP7_75t_L g3556 ( 
.A(n_3395),
.B(n_3117),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3384),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3330),
.B(n_3156),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3497),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3356),
.B(n_3160),
.Y(n_3560)
);

AND2x4_ASAP7_75t_L g3561 ( 
.A(n_3443),
.B(n_3271),
.Y(n_3561)
);

OR2x2_ASAP7_75t_L g3562 ( 
.A(n_3506),
.B(n_3082),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3451),
.B(n_3166),
.Y(n_3563)
);

BUFx3_ASAP7_75t_L g3564 ( 
.A(n_3426),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3502),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3397),
.B(n_3162),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3436),
.B(n_3470),
.Y(n_3567)
);

OR2x2_ASAP7_75t_L g3568 ( 
.A(n_3450),
.B(n_3082),
.Y(n_3568)
);

OAI21xp5_ASAP7_75t_SL g3569 ( 
.A1(n_3315),
.A2(n_3078),
.B(n_3296),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3351),
.B(n_3230),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3379),
.B(n_3366),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3327),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3478),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3378),
.B(n_3162),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3314),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3346),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3386),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3529),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3420),
.B(n_3192),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3485),
.Y(n_3580)
);

AND2x4_ASAP7_75t_L g3581 ( 
.A(n_3530),
.B(n_3475),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3427),
.B(n_3431),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3507),
.B(n_3231),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3468),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3417),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3409),
.B(n_3192),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3457),
.B(n_3235),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3360),
.B(n_3194),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3368),
.B(n_3194),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3317),
.B(n_3198),
.Y(n_3590)
);

OR2x2_ASAP7_75t_L g3591 ( 
.A(n_3469),
.B(n_3253),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3484),
.B(n_3237),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3522),
.B(n_3239),
.Y(n_3593)
);

NAND2x1p5_ASAP7_75t_L g3594 ( 
.A(n_3328),
.B(n_3149),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3462),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3319),
.B(n_3198),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3345),
.Y(n_3597)
);

AND2x4_ASAP7_75t_L g3598 ( 
.A(n_3448),
.B(n_3271),
.Y(n_3598)
);

AND2x4_ASAP7_75t_SL g3599 ( 
.A(n_3337),
.B(n_3259),
.Y(n_3599)
);

INVxp67_ASAP7_75t_L g3600 ( 
.A(n_3376),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3407),
.Y(n_3601)
);

INVx2_ASAP7_75t_SL g3602 ( 
.A(n_3337),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3519),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_3323),
.Y(n_3604)
);

OR2x2_ASAP7_75t_L g3605 ( 
.A(n_3511),
.B(n_3254),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3483),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3429),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3354),
.B(n_3200),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3401),
.B(n_3200),
.Y(n_3609)
);

HB1xp67_ASAP7_75t_L g3610 ( 
.A(n_3372),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3466),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3515),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3455),
.B(n_3241),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3463),
.B(n_3244),
.Y(n_3614)
);

INVx3_ASAP7_75t_L g3615 ( 
.A(n_3414),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3467),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3465),
.B(n_3246),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3532),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3422),
.B(n_3248),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3343),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3402),
.B(n_3249),
.Y(n_3621)
);

AOI22xp33_ASAP7_75t_L g3622 ( 
.A1(n_3504),
.A2(n_3081),
.B1(n_3181),
.B2(n_3205),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3312),
.B(n_3252),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3347),
.Y(n_3624)
);

OR2x2_ASAP7_75t_L g3625 ( 
.A(n_3421),
.B(n_3254),
.Y(n_3625)
);

INVx3_ASAP7_75t_L g3626 ( 
.A(n_3374),
.Y(n_3626)
);

INVx3_ASAP7_75t_L g3627 ( 
.A(n_3341),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3447),
.Y(n_3628)
);

INVxp67_ASAP7_75t_SL g3629 ( 
.A(n_3391),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3445),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3505),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_L g3632 ( 
.A(n_3490),
.B(n_3205),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3344),
.Y(n_3633)
);

BUFx2_ASAP7_75t_L g3634 ( 
.A(n_3441),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3383),
.Y(n_3635)
);

INVxp67_ASAP7_75t_SL g3636 ( 
.A(n_3406),
.Y(n_3636)
);

NOR2xp33_ASAP7_75t_SL g3637 ( 
.A(n_3418),
.B(n_3158),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3392),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3492),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3486),
.Y(n_3640)
);

INVxp67_ASAP7_75t_L g3641 ( 
.A(n_3362),
.Y(n_3641)
);

BUFx3_ASAP7_75t_L g3642 ( 
.A(n_3564),
.Y(n_3642)
);

OR2x2_ASAP7_75t_L g3643 ( 
.A(n_3567),
.B(n_3247),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3631),
.B(n_3496),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3535),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3571),
.B(n_3413),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3535),
.Y(n_3647)
);

AND2x4_ASAP7_75t_L g3648 ( 
.A(n_3639),
.B(n_3353),
.Y(n_3648)
);

INVxp67_ASAP7_75t_SL g3649 ( 
.A(n_3539),
.Y(n_3649)
);

OR2x2_ASAP7_75t_L g3650 ( 
.A(n_3567),
.B(n_3247),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3539),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3564),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3640),
.B(n_3612),
.Y(n_3653)
);

OAI221xp5_ASAP7_75t_SL g3654 ( 
.A1(n_3548),
.A2(n_3509),
.B1(n_3514),
.B2(n_3418),
.C(n_3482),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3574),
.B(n_3521),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3541),
.Y(n_3656)
);

OAI22xp5_ASAP7_75t_L g3657 ( 
.A1(n_3548),
.A2(n_3348),
.B1(n_3424),
.B2(n_3408),
.Y(n_3657)
);

BUFx2_ASAP7_75t_L g3658 ( 
.A(n_3554),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3591),
.B(n_3264),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3566),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3540),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3597),
.B(n_3211),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3608),
.B(n_3353),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3547),
.Y(n_3664)
);

OR2x2_ASAP7_75t_L g3665 ( 
.A(n_3605),
.B(n_3264),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3557),
.Y(n_3666)
);

NAND3xp33_ASAP7_75t_SL g3667 ( 
.A(n_3637),
.B(n_3430),
.C(n_3416),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3590),
.B(n_3369),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3536),
.Y(n_3669)
);

OAI322xp33_ASAP7_75t_L g3670 ( 
.A1(n_3632),
.A2(n_3477),
.A3(n_3479),
.B1(n_3516),
.B2(n_3513),
.C1(n_3489),
.C2(n_3464),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3562),
.B(n_3242),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3537),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3552),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3596),
.B(n_3623),
.Y(n_3674)
);

OAI321xp33_ASAP7_75t_L g3675 ( 
.A1(n_3622),
.A2(n_3364),
.A3(n_3533),
.B1(n_3415),
.B2(n_3424),
.C(n_3408),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3543),
.Y(n_3676)
);

HB1xp67_ASAP7_75t_L g3677 ( 
.A(n_3550),
.Y(n_3677)
);

AOI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3569),
.A2(n_3461),
.B1(n_3454),
.B2(n_3339),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3551),
.B(n_3342),
.Y(n_3679)
);

OR2x2_ASAP7_75t_L g3680 ( 
.A(n_3570),
.B(n_3592),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3638),
.B(n_3171),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3552),
.Y(n_3682)
);

AOI211xp5_ASAP7_75t_L g3683 ( 
.A1(n_3637),
.A2(n_3412),
.B(n_3388),
.C(n_3440),
.Y(n_3683)
);

NAND3xp33_ASAP7_75t_L g3684 ( 
.A(n_3632),
.B(n_3428),
.C(n_3432),
.Y(n_3684)
);

BUFx6f_ASAP7_75t_L g3685 ( 
.A(n_3602),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3589),
.B(n_3524),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3570),
.B(n_3242),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3572),
.B(n_3214),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3609),
.B(n_3524),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3579),
.B(n_3302),
.Y(n_3690)
);

AOI33xp33_ASAP7_75t_L g3691 ( 
.A1(n_3622),
.A2(n_3371),
.A3(n_3357),
.B1(n_3286),
.B2(n_3296),
.B3(n_3067),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3578),
.B(n_3303),
.Y(n_3692)
);

INVx2_ASAP7_75t_SL g3693 ( 
.A(n_3626),
.Y(n_3693)
);

AND2x4_ASAP7_75t_SL g3694 ( 
.A(n_3626),
.B(n_3326),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3549),
.Y(n_3695)
);

AOI22xp33_ASAP7_75t_L g3696 ( 
.A1(n_3604),
.A2(n_3439),
.B1(n_3435),
.B2(n_3437),
.Y(n_3696)
);

AND2x2_ASAP7_75t_L g3697 ( 
.A(n_3576),
.B(n_3304),
.Y(n_3697)
);

INVxp67_ASAP7_75t_R g3698 ( 
.A(n_3610),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3577),
.B(n_3456),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3575),
.B(n_3216),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3606),
.Y(n_3701)
);

BUFx3_ASAP7_75t_L g3702 ( 
.A(n_3599),
.Y(n_3702)
);

HB1xp67_ASAP7_75t_L g3703 ( 
.A(n_3550),
.Y(n_3703)
);

NAND3xp33_ASAP7_75t_SL g3704 ( 
.A(n_3544),
.B(n_3385),
.C(n_3472),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3534),
.Y(n_3705)
);

NOR2x1_ASAP7_75t_L g3706 ( 
.A(n_3627),
.B(n_3396),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3581),
.B(n_3358),
.Y(n_3707)
);

OAI33xp33_ASAP7_75t_L g3708 ( 
.A1(n_3559),
.A2(n_3476),
.A3(n_3493),
.B1(n_3481),
.B2(n_3373),
.B3(n_3158),
.Y(n_3708)
);

AND2x4_ASAP7_75t_L g3709 ( 
.A(n_3629),
.B(n_3189),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3581),
.B(n_3338),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3586),
.B(n_3298),
.Y(n_3711)
);

OA21x2_ASAP7_75t_L g3712 ( 
.A1(n_3600),
.A2(n_3176),
.B(n_3173),
.Y(n_3712)
);

AOI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3569),
.A2(n_3419),
.B1(n_3433),
.B2(n_3425),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3534),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_3592),
.B(n_3189),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3628),
.B(n_3298),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3553),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3555),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3556),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3588),
.B(n_3350),
.Y(n_3720)
);

NAND3xp33_ASAP7_75t_L g3721 ( 
.A(n_3600),
.B(n_3473),
.C(n_3442),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3565),
.B(n_3270),
.Y(n_3722)
);

OAI21xp33_ASAP7_75t_L g3723 ( 
.A1(n_3629),
.A2(n_3459),
.B(n_3487),
.Y(n_3723)
);

OAI221xp5_ASAP7_75t_L g3724 ( 
.A1(n_3641),
.A2(n_3446),
.B1(n_3334),
.B2(n_3325),
.C(n_3352),
.Y(n_3724)
);

NOR2x1p5_ASAP7_75t_L g3725 ( 
.A(n_3667),
.B(n_3636),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3677),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3703),
.Y(n_3727)
);

INVxp67_ASAP7_75t_L g3728 ( 
.A(n_3658),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3652),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3645),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3653),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3647),
.Y(n_3732)
);

NAND2x1_ASAP7_75t_L g3733 ( 
.A(n_3706),
.B(n_3627),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3717),
.Y(n_3734)
);

BUFx2_ASAP7_75t_L g3735 ( 
.A(n_3642),
.Y(n_3735)
);

AND2x4_ASAP7_75t_L g3736 ( 
.A(n_3706),
.B(n_3636),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3663),
.B(n_3610),
.Y(n_3737)
);

NOR2x1p5_ASAP7_75t_L g3738 ( 
.A(n_3704),
.B(n_3603),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3718),
.Y(n_3739)
);

OR2x2_ASAP7_75t_L g3740 ( 
.A(n_3680),
.B(n_3568),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3705),
.B(n_3558),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3698),
.B(n_3674),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3714),
.B(n_3560),
.Y(n_3743)
);

OR2x2_ASAP7_75t_L g3744 ( 
.A(n_3643),
.B(n_3583),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3673),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3682),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3720),
.B(n_3615),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3661),
.Y(n_3748)
);

AND2x4_ASAP7_75t_L g3749 ( 
.A(n_3648),
.B(n_3641),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3664),
.Y(n_3750)
);

INVxp33_ASAP7_75t_L g3751 ( 
.A(n_3685),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3666),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3644),
.B(n_3583),
.Y(n_3753)
);

OR2x2_ASAP7_75t_L g3754 ( 
.A(n_3650),
.B(n_3580),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3710),
.B(n_3615),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3707),
.B(n_3544),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3659),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3649),
.B(n_3563),
.Y(n_3758)
);

BUFx2_ASAP7_75t_L g3759 ( 
.A(n_3685),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3719),
.B(n_3621),
.Y(n_3760)
);

OR2x2_ASAP7_75t_L g3761 ( 
.A(n_3671),
.B(n_3573),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3665),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3656),
.B(n_3621),
.Y(n_3763)
);

AND2x4_ASAP7_75t_L g3764 ( 
.A(n_3648),
.B(n_3620),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3655),
.B(n_3587),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3686),
.B(n_3689),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3690),
.B(n_3587),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3651),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3711),
.B(n_3613),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3715),
.Y(n_3770)
);

INVxp67_ASAP7_75t_L g3771 ( 
.A(n_3721),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3722),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3660),
.B(n_3582),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3662),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3687),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3668),
.B(n_3618),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3701),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3669),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3672),
.Y(n_3779)
);

NAND2x1_ASAP7_75t_SL g3780 ( 
.A(n_3713),
.B(n_3595),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3676),
.Y(n_3781)
);

INVxp33_ASAP7_75t_L g3782 ( 
.A(n_3685),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3695),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3679),
.B(n_3630),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3681),
.B(n_3614),
.Y(n_3785)
);

AND2x4_ASAP7_75t_L g3786 ( 
.A(n_3709),
.B(n_3616),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3697),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3693),
.B(n_3619),
.Y(n_3788)
);

AND2x4_ASAP7_75t_L g3789 ( 
.A(n_3709),
.B(n_3617),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3681),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3699),
.B(n_3633),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3712),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3712),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3646),
.B(n_3611),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3688),
.Y(n_3795)
);

NAND2xp33_ASAP7_75t_SL g3796 ( 
.A(n_3780),
.B(n_3657),
.Y(n_3796)
);

INVxp67_ASAP7_75t_L g3797 ( 
.A(n_3735),
.Y(n_3797)
);

OAI221xp5_ASAP7_75t_L g3798 ( 
.A1(n_3771),
.A2(n_3654),
.B1(n_3713),
.B2(n_3678),
.C(n_3724),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_3736),
.B(n_3657),
.Y(n_3799)
);

AO221x2_ASAP7_75t_L g3800 ( 
.A1(n_3792),
.A2(n_3721),
.B1(n_3335),
.B2(n_3684),
.C(n_3607),
.Y(n_3800)
);

NOR2xp33_ASAP7_75t_R g3801 ( 
.A(n_3742),
.B(n_3320),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3785),
.Y(n_3802)
);

OAI221xp5_ASAP7_75t_L g3803 ( 
.A1(n_3728),
.A2(n_3678),
.B1(n_3684),
.B2(n_3723),
.C(n_3683),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3790),
.B(n_3692),
.Y(n_3804)
);

NAND2xp33_ASAP7_75t_SL g3805 ( 
.A(n_3725),
.B(n_3634),
.Y(n_3805)
);

BUFx2_ASAP7_75t_L g3806 ( 
.A(n_3759),
.Y(n_3806)
);

NAND2xp33_ASAP7_75t_SL g3807 ( 
.A(n_3738),
.B(n_3546),
.Y(n_3807)
);

OAI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3736),
.A2(n_3675),
.B(n_3723),
.Y(n_3808)
);

OAI22xp33_ASAP7_75t_L g3809 ( 
.A1(n_3733),
.A2(n_3675),
.B1(n_3400),
.B2(n_3405),
.Y(n_3809)
);

OAI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3751),
.A2(n_3359),
.B1(n_3702),
.B2(n_3367),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3795),
.B(n_3716),
.Y(n_3811)
);

NAND2xp33_ASAP7_75t_SL g3812 ( 
.A(n_3749),
.B(n_3390),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3795),
.B(n_3700),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_3731),
.B(n_3708),
.Y(n_3814)
);

AO221x2_ASAP7_75t_L g3815 ( 
.A1(n_3792),
.A2(n_3585),
.B1(n_3584),
.B2(n_3670),
.C(n_3452),
.Y(n_3815)
);

NAND2xp33_ASAP7_75t_SL g3816 ( 
.A(n_3749),
.B(n_3696),
.Y(n_3816)
);

INVxp67_ASAP7_75t_L g3817 ( 
.A(n_3729),
.Y(n_3817)
);

AO221x2_ASAP7_75t_L g3818 ( 
.A1(n_3793),
.A2(n_3670),
.B1(n_3683),
.B2(n_3316),
.C(n_3313),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3772),
.B(n_3614),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3774),
.B(n_3593),
.Y(n_3820)
);

NAND2xp33_ASAP7_75t_SL g3821 ( 
.A(n_3782),
.B(n_3370),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_3756),
.B(n_3694),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3763),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3726),
.B(n_3593),
.Y(n_3824)
);

INVx3_ASAP7_75t_L g3825 ( 
.A(n_3789),
.Y(n_3825)
);

AO221x2_ASAP7_75t_L g3826 ( 
.A1(n_3793),
.A2(n_3500),
.B1(n_3601),
.B2(n_3322),
.C(n_3324),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3760),
.B(n_3365),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_3794),
.Y(n_3828)
);

NOR2xp33_ASAP7_75t_L g3829 ( 
.A(n_3789),
.B(n_3349),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3726),
.B(n_3538),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_R g3831 ( 
.A(n_3788),
.B(n_3332),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3727),
.B(n_3775),
.Y(n_3832)
);

OAI221xp5_ASAP7_75t_L g3833 ( 
.A1(n_3765),
.A2(n_3331),
.B1(n_3377),
.B2(n_3438),
.C(n_3594),
.Y(n_3833)
);

AOI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_3770),
.A2(n_3757),
.B1(n_3762),
.B2(n_3737),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3727),
.B(n_3538),
.Y(n_3835)
);

AO221x2_ASAP7_75t_L g3836 ( 
.A1(n_3758),
.A2(n_3349),
.B1(n_3321),
.B2(n_3336),
.C(n_3404),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3745),
.B(n_3542),
.Y(n_3837)
);

HB1xp67_ASAP7_75t_L g3838 ( 
.A(n_3730),
.Y(n_3838)
);

OAI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3740),
.A2(n_3363),
.B1(n_3594),
.B2(n_3545),
.Y(n_3839)
);

OR2x2_ASAP7_75t_L g3840 ( 
.A(n_3744),
.B(n_3542),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3746),
.B(n_3598),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3797),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3823),
.Y(n_3843)
);

OA22x2_ASAP7_75t_L g3844 ( 
.A1(n_3808),
.A2(n_3786),
.B1(n_3764),
.B2(n_3434),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3836),
.B(n_3786),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3836),
.B(n_3766),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3826),
.B(n_3764),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3824),
.Y(n_3848)
);

OR2x2_ASAP7_75t_L g3849 ( 
.A(n_3802),
.B(n_3767),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3832),
.Y(n_3850)
);

AND2x4_ASAP7_75t_L g3851 ( 
.A(n_3825),
.B(n_3791),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3806),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3840),
.Y(n_3853)
);

INVx1_ASAP7_75t_SL g3854 ( 
.A(n_3801),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3830),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3826),
.B(n_3747),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3835),
.Y(n_3857)
);

INVxp67_ASAP7_75t_SL g3858 ( 
.A(n_3814),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3813),
.B(n_3753),
.Y(n_3859)
);

NOR2x1_ASAP7_75t_L g3860 ( 
.A(n_3803),
.B(n_3396),
.Y(n_3860)
);

HB1xp67_ASAP7_75t_L g3861 ( 
.A(n_3838),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3819),
.Y(n_3862)
);

AND2x4_ASAP7_75t_L g3863 ( 
.A(n_3822),
.B(n_3829),
.Y(n_3863)
);

HB1xp67_ASAP7_75t_L g3864 ( 
.A(n_3818),
.Y(n_3864)
);

HB1xp67_ASAP7_75t_L g3865 ( 
.A(n_3818),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3800),
.B(n_3755),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3817),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3800),
.B(n_3815),
.Y(n_3868)
);

INVx1_ASAP7_75t_SL g3869 ( 
.A(n_3831),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3820),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3815),
.B(n_3776),
.Y(n_3871)
);

AOI22xp33_ASAP7_75t_L g3872 ( 
.A1(n_3798),
.A2(n_3375),
.B1(n_3449),
.B2(n_3517),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3837),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3834),
.B(n_3730),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3811),
.B(n_3748),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3804),
.B(n_3750),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3841),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3799),
.B(n_3787),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3816),
.B(n_3761),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3809),
.B(n_3752),
.Y(n_3880)
);

CKINVDCx16_ASAP7_75t_R g3881 ( 
.A(n_3821),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3828),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3827),
.Y(n_3883)
);

CKINVDCx16_ASAP7_75t_R g3884 ( 
.A(n_3807),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3796),
.B(n_3734),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3805),
.B(n_3773),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3812),
.B(n_3777),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3833),
.B(n_3739),
.Y(n_3888)
);

AND2x2_ASAP7_75t_L g3889 ( 
.A(n_3810),
.B(n_3784),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3839),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3836),
.B(n_3741),
.Y(n_3891)
);

INVx1_ASAP7_75t_SL g3892 ( 
.A(n_3801),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3847),
.B(n_3743),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3842),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3844),
.A2(n_3444),
.B(n_3769),
.Y(n_3895)
);

OAI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3844),
.A2(n_3754),
.B1(n_3526),
.B2(n_3528),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3884),
.B(n_3768),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3858),
.B(n_3778),
.Y(n_3898)
);

AOI22xp33_ASAP7_75t_L g3899 ( 
.A1(n_3868),
.A2(n_3410),
.B1(n_3598),
.B2(n_3340),
.Y(n_3899)
);

OAI22xp33_ASAP7_75t_L g3900 ( 
.A1(n_3879),
.A2(n_3518),
.B1(n_3545),
.B2(n_3508),
.Y(n_3900)
);

AOI22xp33_ASAP7_75t_L g3901 ( 
.A1(n_3864),
.A2(n_3865),
.B1(n_3860),
.B2(n_3891),
.Y(n_3901)
);

CKINVDCx16_ASAP7_75t_R g3902 ( 
.A(n_3854),
.Y(n_3902)
);

OAI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3864),
.A2(n_3410),
.B(n_3145),
.Y(n_3903)
);

INVxp67_ASAP7_75t_SL g3904 ( 
.A(n_3842),
.Y(n_3904)
);

INVxp67_ASAP7_75t_L g3905 ( 
.A(n_3882),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3892),
.B(n_3732),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3861),
.Y(n_3907)
);

OAI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3865),
.A2(n_3783),
.B1(n_3781),
.B2(n_3779),
.Y(n_3908)
);

OAI32xp33_ASAP7_75t_L g3909 ( 
.A1(n_3881),
.A2(n_3361),
.A3(n_3625),
.B1(n_3635),
.B2(n_3624),
.Y(n_3909)
);

NOR3xp33_ASAP7_75t_L g3910 ( 
.A(n_3858),
.B(n_3276),
.C(n_2999),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3845),
.B(n_3561),
.Y(n_3911)
);

OAI221xp5_ASAP7_75t_L g3912 ( 
.A1(n_3885),
.A2(n_3145),
.B1(n_3286),
.B2(n_3508),
.C(n_3257),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3861),
.Y(n_3913)
);

NOR2xp33_ASAP7_75t_L g3914 ( 
.A(n_3869),
.B(n_3527),
.Y(n_3914)
);

AOI21xp33_ASAP7_75t_L g3915 ( 
.A1(n_3890),
.A2(n_2841),
.B(n_3494),
.Y(n_3915)
);

INVx1_ASAP7_75t_SL g3916 ( 
.A(n_3852),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3876),
.Y(n_3917)
);

OAI21xp5_ASAP7_75t_SL g3918 ( 
.A1(n_3872),
.A2(n_2937),
.B(n_2988),
.Y(n_3918)
);

INVx3_ASAP7_75t_L g3919 ( 
.A(n_3863),
.Y(n_3919)
);

INVx1_ASAP7_75t_SL g3920 ( 
.A(n_3867),
.Y(n_3920)
);

AOI322xp5_ASAP7_75t_L g3921 ( 
.A1(n_3872),
.A2(n_3561),
.A3(n_3503),
.B1(n_3276),
.B2(n_3273),
.C1(n_3274),
.C2(n_3184),
.Y(n_3921)
);

OAI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3885),
.A2(n_2994),
.B(n_2765),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3876),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3853),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3849),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_3902),
.B(n_3919),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3920),
.B(n_3850),
.Y(n_3927)
);

NOR2x1_ASAP7_75t_L g3928 ( 
.A(n_3896),
.B(n_3856),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_3919),
.B(n_3863),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3920),
.B(n_3862),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3916),
.B(n_3904),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3894),
.Y(n_3932)
);

NOR2x1_ASAP7_75t_L g3933 ( 
.A(n_3907),
.B(n_3846),
.Y(n_3933)
);

NAND2x1_ASAP7_75t_SL g3934 ( 
.A(n_3913),
.B(n_3866),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3916),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3905),
.B(n_3870),
.Y(n_3936)
);

OAI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3895),
.A2(n_3880),
.B1(n_3888),
.B2(n_3871),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3897),
.B(n_3886),
.Y(n_3938)
);

AND2x2_ASAP7_75t_L g3939 ( 
.A(n_3911),
.B(n_3878),
.Y(n_3939)
);

NAND3xp33_ASAP7_75t_L g3940 ( 
.A(n_3901),
.B(n_3880),
.C(n_3888),
.Y(n_3940)
);

INVxp67_ASAP7_75t_SL g3941 ( 
.A(n_3906),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3921),
.B(n_3917),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3923),
.B(n_3873),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3898),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3914),
.B(n_3883),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3924),
.Y(n_3946)
);

NAND2xp33_ASAP7_75t_SL g3947 ( 
.A(n_3899),
.B(n_3488),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3925),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3910),
.B(n_3855),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3893),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3935),
.Y(n_3951)
);

HB1xp67_ASAP7_75t_L g3952 ( 
.A(n_3931),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3946),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3930),
.Y(n_3954)
);

CKINVDCx5p33_ASAP7_75t_R g3955 ( 
.A(n_3926),
.Y(n_3955)
);

INVxp33_ASAP7_75t_SL g3956 ( 
.A(n_3929),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3927),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3936),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3950),
.Y(n_3959)
);

CKINVDCx5p33_ASAP7_75t_R g3960 ( 
.A(n_3941),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3945),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3932),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3948),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3943),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3944),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3945),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3938),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3949),
.Y(n_3968)
);

INVxp33_ASAP7_75t_SL g3969 ( 
.A(n_3928),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3939),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3933),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3940),
.Y(n_3972)
);

INVx1_ASAP7_75t_SL g3973 ( 
.A(n_3947),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3960),
.B(n_3940),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3969),
.B(n_3937),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3955),
.B(n_3900),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3972),
.B(n_3951),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3956),
.A2(n_3942),
.B(n_3909),
.Y(n_3978)
);

NOR3x1_ASAP7_75t_L g3979 ( 
.A(n_3966),
.B(n_3903),
.C(n_3918),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3951),
.B(n_3934),
.Y(n_3980)
);

AOI222xp33_ASAP7_75t_L g3981 ( 
.A1(n_3952),
.A2(n_3912),
.B1(n_3908),
.B2(n_3922),
.C1(n_3874),
.C2(n_3889),
.Y(n_3981)
);

NAND3xp33_ASAP7_75t_L g3982 ( 
.A(n_3952),
.B(n_3915),
.C(n_3887),
.Y(n_3982)
);

AOI221xp5_ASAP7_75t_L g3983 ( 
.A1(n_3970),
.A2(n_3874),
.B1(n_3857),
.B2(n_3848),
.C(n_3877),
.Y(n_3983)
);

OAI211xp5_ASAP7_75t_SL g3984 ( 
.A1(n_3973),
.A2(n_3843),
.B(n_3875),
.C(n_2974),
.Y(n_3984)
);

OAI221xp5_ASAP7_75t_L g3985 ( 
.A1(n_3971),
.A2(n_3875),
.B1(n_3859),
.B2(n_2869),
.C(n_3042),
.Y(n_3985)
);

NAND3xp33_ASAP7_75t_SL g3986 ( 
.A(n_3953),
.B(n_3510),
.C(n_3498),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3967),
.Y(n_3987)
);

NAND3xp33_ASAP7_75t_L g3988 ( 
.A(n_3968),
.B(n_2979),
.C(n_3851),
.Y(n_3988)
);

NAND3xp33_ASAP7_75t_L g3989 ( 
.A(n_3953),
.B(n_2979),
.C(n_3851),
.Y(n_3989)
);

OAI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_3978),
.A2(n_3957),
.B(n_3954),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3975),
.A2(n_3961),
.B(n_3958),
.Y(n_3991)
);

HB1xp67_ASAP7_75t_L g3992 ( 
.A(n_3987),
.Y(n_3992)
);

OAI211xp5_ASAP7_75t_SL g3993 ( 
.A1(n_3974),
.A2(n_3965),
.B(n_3964),
.C(n_3959),
.Y(n_3993)
);

AOI22xp5_ASAP7_75t_L g3994 ( 
.A1(n_3986),
.A2(n_3967),
.B1(n_3963),
.B2(n_3962),
.Y(n_3994)
);

AOI211xp5_ASAP7_75t_SL g3995 ( 
.A1(n_3977),
.A2(n_2892),
.B(n_3048),
.C(n_3018),
.Y(n_3995)
);

OAI211xp5_ASAP7_75t_SL g3996 ( 
.A1(n_3976),
.A2(n_3980),
.B(n_3981),
.C(n_3982),
.Y(n_3996)
);

OAI322xp33_ASAP7_75t_L g3997 ( 
.A1(n_3988),
.A2(n_2948),
.A3(n_2963),
.B1(n_2939),
.B2(n_3070),
.C1(n_2805),
.C2(n_2845),
.Y(n_3997)
);

OAI211xp5_ASAP7_75t_SL g3998 ( 
.A1(n_3983),
.A2(n_3989),
.B(n_3979),
.C(n_3985),
.Y(n_3998)
);

O2A1O1Ixp33_ASAP7_75t_L g3999 ( 
.A1(n_3984),
.A2(n_2902),
.B(n_2917),
.C(n_2870),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3977),
.Y(n_4000)
);

AOI221xp5_ASAP7_75t_L g4001 ( 
.A1(n_3978),
.A2(n_3512),
.B1(n_3523),
.B2(n_2989),
.C(n_3411),
.Y(n_4001)
);

OAI221xp5_ASAP7_75t_L g4002 ( 
.A1(n_3978),
.A2(n_3022),
.B1(n_2945),
.B2(n_2960),
.C(n_2943),
.Y(n_4002)
);

OAI211xp5_ASAP7_75t_SL g4003 ( 
.A1(n_3974),
.A2(n_3068),
.B(n_3691),
.C(n_3071),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3992),
.Y(n_4004)
);

AOI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_3996),
.A2(n_3525),
.B1(n_3221),
.B2(n_3300),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_4000),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3991),
.B(n_813),
.Y(n_4007)
);

CKINVDCx16_ASAP7_75t_R g4008 ( 
.A(n_3990),
.Y(n_4008)
);

AND2x4_ASAP7_75t_L g4009 ( 
.A(n_3994),
.B(n_3480),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3993),
.Y(n_4010)
);

NAND2xp33_ASAP7_75t_R g4011 ( 
.A(n_4007),
.B(n_3998),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_4008),
.B(n_4001),
.Y(n_4012)
);

XNOR2xp5_ASAP7_75t_L g4013 ( 
.A(n_4009),
.B(n_4004),
.Y(n_4013)
);

XNOR2xp5_ASAP7_75t_L g4014 ( 
.A(n_4006),
.B(n_4002),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_R g4015 ( 
.A(n_4010),
.B(n_814),
.Y(n_4015)
);

NAND2x1_ASAP7_75t_L g4016 ( 
.A(n_4012),
.B(n_4013),
.Y(n_4016)
);

AOI22xp5_ASAP7_75t_SL g4017 ( 
.A1(n_4014),
.A2(n_4003),
.B1(n_3995),
.B2(n_4005),
.Y(n_4017)
);

NOR3xp33_ASAP7_75t_L g4018 ( 
.A(n_4016),
.B(n_4015),
.C(n_4011),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_4017),
.A2(n_3999),
.B(n_3997),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_SL g4020 ( 
.A(n_4018),
.B(n_3394),
.Y(n_4020)
);

NOR2xp33_ASAP7_75t_L g4021 ( 
.A(n_4019),
.B(n_814),
.Y(n_4021)
);

AOI31xp33_ASAP7_75t_L g4022 ( 
.A1(n_4021),
.A2(n_2864),
.A3(n_818),
.B(n_815),
.Y(n_4022)
);

AOI31xp33_ASAP7_75t_L g4023 ( 
.A1(n_4020),
.A2(n_818),
.A3(n_815),
.B(n_816),
.Y(n_4023)
);

OAI322xp33_ASAP7_75t_L g4024 ( 
.A1(n_4023),
.A2(n_3265),
.A3(n_3154),
.B1(n_3520),
.B2(n_3180),
.C1(n_3177),
.C2(n_3399),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_4024),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_4025),
.Y(n_4026)
);

AOI221xp5_ASAP7_75t_L g4027 ( 
.A1(n_4026),
.A2(n_4022),
.B1(n_3049),
.B2(n_2832),
.C(n_3221),
.Y(n_4027)
);

AOI211xp5_ASAP7_75t_L g4028 ( 
.A1(n_4027),
.A2(n_821),
.B(n_816),
.C(n_820),
.Y(n_4028)
);


endmodule