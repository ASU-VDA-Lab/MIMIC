module fake_netlist_5_1697_n_1826 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1826);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1826;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_SL g194 ( 
.A(n_38),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_123),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_31),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_42),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_18),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_101),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_65),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_88),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_94),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_125),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_77),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_151),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_92),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_159),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_54),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_139),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_38),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_164),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_63),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_47),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_17),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_56),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_115),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_98),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_76),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_114),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_131),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_14),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_5),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_122),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_28),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_121),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_90),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_130),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_18),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_136),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_66),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_96),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_158),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_116),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_23),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_32),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_162),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_105),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_150),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_11),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_4),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_144),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_48),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_58),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_124),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_42),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_87),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_183),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_128),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_75),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_129),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_182),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_5),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_107),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_157),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_135),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_29),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_188),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_0),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_110),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_152),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_8),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_4),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_52),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_142),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_17),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_108),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_181),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_12),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_172),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_177),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_45),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_184),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_36),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_137),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_81),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_106),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_84),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_154),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_73),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_138),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_179),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_132),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_80),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_167),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_3),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_166),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_119),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_78),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_48),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_2),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_59),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_40),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_143),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_6),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_153),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_103),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_16),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_120),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_91),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_165),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_155),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_13),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_111),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_12),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_23),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_34),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_72),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_145),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_163),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_71),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_10),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_99),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_36),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_58),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_74),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_160),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_60),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_25),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_187),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_68),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_50),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_146),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_51),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_51),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_176),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_186),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_82),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_15),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_64),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_45),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_15),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_53),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_6),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_173),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_41),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_10),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_30),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_140),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_33),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_102),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_52),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_79),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_26),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_83),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_126),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_190),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_67),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_28),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_70),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_156),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_62),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_174),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_35),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_19),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_3),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_34),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_1),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_20),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_22),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_27),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_85),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_291),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_388),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_228),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_228),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_212),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_228),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_228),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_228),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_224),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_228),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_228),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_376),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_228),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_393),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_391),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_196),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_229),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_271),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_243),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_249),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_212),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_197),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_198),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_257),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_267),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_292),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_248),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_293),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_271),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_327),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_236),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_368),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_220),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_386),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_211),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_208),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_208),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_308),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_225),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_308),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_313),
.Y(n_450)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_386),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_313),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_226),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_271),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_201),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_227),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_204),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_230),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_238),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_218),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_235),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_247),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_337),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_254),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_258),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_351),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_282),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_283),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_295),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_294),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_387),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_302),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_331),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_294),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_340),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_239),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_387),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_244),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_350),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_352),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_389),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_251),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_371),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_263),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_367),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_219),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_219),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_223),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_223),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_338),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_237),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_294),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_237),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_471),
.A2(n_389),
.B1(n_390),
.B2(n_217),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_417),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_417),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_437),
.B(n_241),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g509 ( 
.A(n_398),
.B(n_319),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_424),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_403),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_400),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_406),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_207),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_404),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_407),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_409),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_395),
.B(n_272),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_406),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_487),
.B(n_367),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_334),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_424),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_418),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_420),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_471),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_445),
.B(n_446),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_477),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_425),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_395),
.B(n_200),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_396),
.B(n_200),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_447),
.B(n_270),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

NOR2x1_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_367),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_450),
.B(n_270),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_425),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_474),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_467),
.B(n_273),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_452),
.B(n_194),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_427),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_467),
.B(n_273),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_495),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_434),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_455),
.B(n_259),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_435),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_495),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_439),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_427),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_431),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_408),
.A2(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_490),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_416),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_438),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_457),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_538),
.B(n_460),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_538),
.B(n_259),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_396),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_509),
.B(n_439),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_500),
.B(n_416),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_530),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_501),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_532),
.B(n_440),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_557),
.B(n_461),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_530),
.B(n_462),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_514),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_514),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_555),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_502),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_530),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_511),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_517),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_522),
.B(n_448),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_514),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_440),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_520),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_543),
.B(n_451),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_523),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_509),
.A2(n_465),
.B1(n_468),
.B2(n_464),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_520),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_557),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_399),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_520),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_523),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_525),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_521),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_525),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_557),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_526),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_526),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_557),
.B(n_469),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_521),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_521),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_561),
.B(n_472),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_529),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_561),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_SL g628 ( 
.A(n_513),
.B(n_448),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_509),
.A2(n_451),
.B1(n_456),
.B2(n_453),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_529),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_529),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_564),
.A2(n_552),
.B(n_544),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_506),
.B(n_453),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_545),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_506),
.B(n_456),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_545),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_508),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_512),
.A2(n_347),
.B1(n_322),
.B2(n_285),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_545),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_556),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_561),
.B(n_533),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_558),
.A2(n_475),
.B1(n_479),
.B2(n_473),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_506),
.B(n_458),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_558),
.B(n_480),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_533),
.B(n_481),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_556),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_534),
.B(n_458),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_555),
.B(n_484),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_515),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_541),
.B(n_459),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_497),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_555),
.B(n_486),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_554),
.B(n_459),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_562),
.Y(n_655)
);

AND3x2_ASAP7_75t_L g656 ( 
.A(n_550),
.B(n_278),
.C(n_276),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_524),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_562),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_555),
.B(n_488),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_573),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_546),
.B(n_276),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_497),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_497),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_567),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_566),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_555),
.B(n_476),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_531),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_566),
.Y(n_669)
);

NOR2x1p5_ASAP7_75t_L g670 ( 
.A(n_535),
.B(n_338),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_566),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_559),
.B(n_431),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_547),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_547),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_498),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_498),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_547),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_547),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_531),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_531),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_508),
.B(n_476),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_499),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_531),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_531),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_578),
.B(n_478),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_499),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_531),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_504),
.B(n_478),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_510),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_503),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_546),
.B(n_278),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_568),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_504),
.B(n_483),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_503),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_510),
.Y(n_695)
);

INVxp33_ASAP7_75t_SL g696 ( 
.A(n_537),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_505),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_504),
.B(n_483),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_510),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_505),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_507),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_535),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_536),
.Y(n_703)
);

INVxp33_ASAP7_75t_L g704 ( 
.A(n_537),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_524),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_507),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_578),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_578),
.B(n_493),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_575),
.Y(n_709)
);

CKINVDCx6p67_ASAP7_75t_R g710 ( 
.A(n_569),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_536),
.B(n_485),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_508),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_575),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_575),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_575),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_540),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_524),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_510),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_R g720 ( 
.A(n_508),
.B(n_485),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_540),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_539),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_548),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_548),
.A2(n_262),
.B1(n_306),
.B2(n_194),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_549),
.B(n_422),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_549),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_551),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_551),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_553),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_710),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_710),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_609),
.B(n_572),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_609),
.B(n_617),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_729),
.B(n_419),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_585),
.B(n_553),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_617),
.B(n_572),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_582),
.A2(n_261),
.B1(n_245),
.B2(n_240),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_588),
.A2(n_214),
.B1(n_203),
.B2(n_195),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_590),
.A2(n_560),
.B(n_563),
.C(n_574),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_729),
.B(n_432),
.Y(n_741)
);

OAI22x1_ASAP7_75t_SL g742 ( 
.A1(n_696),
.A2(n_466),
.B1(n_463),
.B2(n_436),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_596),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_596),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_627),
.A2(n_262),
.B1(n_306),
.B2(n_374),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_627),
.B(n_572),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_673),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_606),
.B(n_572),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_716),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_602),
.A2(n_311),
.B1(n_332),
.B2(n_377),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_605),
.B(n_477),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_606),
.B(n_584),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_716),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_726),
.B(n_482),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_591),
.A2(n_518),
.B(n_516),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_728),
.B(n_482),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_725),
.A2(n_374),
.B(n_405),
.C(n_574),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_591),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_673),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_674),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_723),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_584),
.B(n_572),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_597),
.B(n_572),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_591),
.B(n_336),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_723),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_597),
.B(n_577),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_600),
.A2(n_298),
.B1(n_316),
.B2(n_305),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_728),
.B(n_711),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_674),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_629),
.B(n_635),
.C(n_633),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_667),
.B(n_294),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_702),
.B(n_336),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_702),
.B(n_336),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_644),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_598),
.B(n_577),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_644),
.B(n_454),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_598),
.B(n_577),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_677),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_675),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_563),
.C(n_560),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_685),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_577),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_702),
.B(n_375),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_643),
.A2(n_280),
.B1(n_233),
.B2(n_394),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_603),
.B(n_577),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_675),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_649),
.B(n_430),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_610),
.B(n_430),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_676),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_676),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_612),
.B(n_577),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_589),
.A2(n_279),
.B1(n_222),
.B2(n_221),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_612),
.B(n_518),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_613),
.B(n_518),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_690),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_589),
.A2(n_315),
.B1(n_260),
.B2(n_255),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_697),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_677),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_660),
.B(n_430),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_579),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_678),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_621),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_678),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_616),
.B(n_504),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_616),
.B(n_516),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_688),
.B(n_294),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_632),
.A2(n_307),
.B1(n_355),
.B2(n_375),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_625),
.A2(n_277),
.B1(n_231),
.B2(n_232),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_625),
.A2(n_284),
.B1(n_234),
.B2(n_242),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_638),
.B(n_565),
.C(n_443),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_618),
.B(n_375),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_670),
.Y(n_813)
);

NOR2xp67_ASAP7_75t_L g814 ( 
.A(n_581),
.B(n_565),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_632),
.A2(n_321),
.B1(n_246),
.B2(n_250),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_592),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_632),
.A2(n_580),
.B1(n_698),
.B2(n_693),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_592),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_618),
.B(n_516),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_593),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_610),
.B(n_287),
.C(n_281),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_703),
.B(n_199),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_697),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_620),
.B(n_375),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_593),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_620),
.B(n_294),
.Y(n_826)
);

BUFx5_ASAP7_75t_L g827 ( 
.A(n_709),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_703),
.B(n_442),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_622),
.A2(n_444),
.B(n_307),
.C(n_355),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_706),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_580),
.A2(n_268),
.B1(n_252),
.B2(n_253),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_587),
.B(n_595),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_721),
.B(n_516),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_579),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_708),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_601),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_670),
.A2(n_360),
.B1(n_294),
.B2(n_289),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_601),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_641),
.A2(n_576),
.B(n_571),
.C(n_274),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_721),
.B(n_519),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_708),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_727),
.B(n_199),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_727),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_647),
.B(n_202),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_682),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_580),
.A2(n_264),
.B1(n_275),
.B2(n_286),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_682),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_587),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_689),
.B(n_519),
.Y(n_849)
);

NOR2x1p5_ASAP7_75t_L g850 ( 
.A(n_595),
.B(n_296),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_604),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_604),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_689),
.B(n_519),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_719),
.B(n_519),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_695),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_709),
.B(n_294),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_719),
.B(n_527),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_664),
.B(n_436),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_719),
.B(n_527),
.Y(n_859)
);

AND2x2_ASAP7_75t_SL g860 ( 
.A(n_637),
.B(n_576),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_580),
.B(n_202),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_713),
.B(n_715),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_650),
.B(n_205),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_713),
.B(n_715),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_686),
.B(n_694),
.Y(n_865)
);

OR2x6_ASAP7_75t_L g866 ( 
.A(n_637),
.B(n_463),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_656),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_621),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_583),
.B(n_210),
.C(n_385),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_686),
.B(n_527),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_694),
.B(n_527),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_714),
.B(n_360),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_608),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_700),
.B(n_288),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_700),
.B(n_290),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_608),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_611),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_701),
.B(n_299),
.Y(n_878)
);

AND2x2_ASAP7_75t_SL g879 ( 
.A(n_712),
.B(n_360),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_701),
.Y(n_880)
);

INVxp33_ASAP7_75t_L g881 ( 
.A(n_672),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_714),
.B(n_360),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_707),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_695),
.B(n_301),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_L g885 ( 
.A(n_654),
.B(n_205),
.C(n_209),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_611),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_664),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_718),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_722),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_648),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_699),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_887),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_781),
.B(n_653),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_889),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_883),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_781),
.B(n_659),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_776),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_768),
.B(n_645),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_865),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_845),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_L g901 ( 
.A(n_758),
.B(n_720),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_768),
.B(n_623),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_841),
.B(n_801),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_752),
.B(n_749),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_742),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_753),
.B(n_761),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_758),
.B(n_657),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_SL g908 ( 
.A1(n_757),
.A2(n_724),
.B1(n_642),
.B2(n_681),
.C(n_655),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_751),
.A2(n_834),
.B(n_808),
.C(n_770),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_787),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_847),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_880),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_770),
.A2(n_628),
.B1(n_661),
.B2(n_691),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_889),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_758),
.B(n_657),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_800),
.B(n_704),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_808),
.A2(n_661),
.B1(n_691),
.B2(n_360),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_834),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_758),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_814),
.A2(n_691),
.B1(n_661),
.B2(n_696),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_730),
.B(n_692),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_765),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_817),
.B(n_594),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_754),
.B(n_661),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_879),
.B(n_594),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_779),
.B(n_623),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_754),
.B(n_594),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_816),
.Y(n_928)
);

BUFx6f_ASAP7_75t_SL g929 ( 
.A(n_731),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_736),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_786),
.B(n_624),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_735),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_837),
.A2(n_661),
.B1(n_691),
.B2(n_360),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_818),
.Y(n_934)
);

OR2x2_ASAP7_75t_SL g935 ( 
.A(n_821),
.B(n_297),
.Y(n_935)
);

AND2x6_ASAP7_75t_L g936 ( 
.A(n_732),
.B(n_624),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_820),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_825),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_803),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_837),
.A2(n_691),
.B1(n_360),
.B2(n_634),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_736),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_SL g942 ( 
.A1(n_788),
.A2(n_318),
.B1(n_300),
.B2(n_303),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_855),
.B(n_705),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_789),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_890),
.A2(n_360),
.B1(n_639),
.B2(n_634),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_855),
.B(n_705),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_790),
.B(n_631),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_750),
.B(n_615),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_774),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_836),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_793),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_838),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_835),
.A2(n_639),
.B1(n_640),
.B2(n_646),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_796),
.B(n_631),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_739),
.A2(n_615),
.B1(n_216),
.B2(n_215),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_827),
.B(n_652),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_866),
.B(n_717),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_741),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_SL g959 ( 
.A(n_738),
.B(n_357),
.C(n_356),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_756),
.B(n_304),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_798),
.B(n_655),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_823),
.B(n_658),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_851),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_852),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_743),
.A2(n_744),
.B1(n_815),
.B2(n_734),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_830),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_843),
.B(n_658),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_862),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_885),
.A2(n_671),
.B1(n_614),
.B2(n_626),
.Y(n_969)
);

NAND2xp33_ASAP7_75t_SL g970 ( 
.A(n_813),
.B(n_206),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_858),
.B(n_206),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_873),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_844),
.A2(n_671),
.B1(n_599),
.B2(n_683),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_827),
.B(n_652),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_827),
.B(n_652),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_864),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_866),
.B(n_717),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_803),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_822),
.B(n_614),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_805),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_822),
.B(n_626),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_806),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_827),
.B(n_652),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_L g984 ( 
.A(n_827),
.B(n_717),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_885),
.A2(n_651),
.B1(n_630),
.B2(n_636),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_819),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_844),
.A2(n_586),
.B1(n_599),
.B2(n_683),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_867),
.B(n_717),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_868),
.B(n_828),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_881),
.A2(n_323),
.B1(n_330),
.B2(n_335),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_876),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_868),
.B(n_717),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_877),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_842),
.B(n_630),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_747),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_863),
.A2(n_586),
.B1(n_599),
.B2(n_683),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_828),
.B(n_619),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_886),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_863),
.A2(n_619),
.B1(n_662),
.B2(n_679),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_756),
.B(n_788),
.Y(n_1000)
);

NOR2x1p5_ASAP7_75t_L g1001 ( 
.A(n_780),
.B(n_339),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_860),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_745),
.A2(n_636),
.B1(n_651),
.B2(n_665),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_842),
.B(n_665),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_L g1005 ( 
.A(n_811),
.B(n_354),
.C(n_344),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_759),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_361),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_866),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_767),
.B(n_684),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_888),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_811),
.B(n_364),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_861),
.B(n_370),
.Y(n_1012)
);

OR2x2_ASAP7_75t_SL g1013 ( 
.A(n_869),
.B(n_372),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_827),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_861),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_748),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_874),
.B(n_684),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_760),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_891),
.B(n_652),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_769),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_875),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_778),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_762),
.B(n_668),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_833),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_757),
.B(n_869),
.Y(n_1025)
);

OR2x2_ASAP7_75t_SL g1026 ( 
.A(n_884),
.B(n_0),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_799),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_878),
.B(n_684),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_802),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_784),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_826),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_772),
.B(n_666),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_740),
.B(n_666),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_772),
.B(n_669),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_840),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_804),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_792),
.B(n_619),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_826),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_773),
.B(n_669),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_745),
.A2(n_213),
.B1(n_215),
.B2(n_373),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_763),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_797),
.B(n_662),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_733),
.A2(n_746),
.B(n_737),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_783),
.B(n_663),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_771),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_766),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_783),
.B(n_663),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_775),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_809),
.B(n_216),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_870),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_810),
.B(n_309),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_871),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_777),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_849),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_782),
.B(n_668),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_794),
.B(n_679),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_R g1057 ( 
.A(n_807),
.B(n_309),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_785),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_853),
.A2(n_687),
.B(n_680),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_791),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_854),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_795),
.B(n_687),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_872),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_831),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_764),
.B(n_668),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_968),
.B(n_899),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_922),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_SL g1069 ( 
.A1(n_925),
.A2(n_764),
.B(n_856),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1014),
.A2(n_859),
.B(n_857),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_898),
.B(n_839),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_895),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1000),
.B(n_846),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1014),
.A2(n_755),
.B(n_680),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_893),
.B(n_872),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_984),
.A2(n_687),
.B(n_680),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_892),
.B(n_882),
.Y(n_1077)
);

BUFx2_ASAP7_75t_SL g1078 ( 
.A(n_892),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_894),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_896),
.B(n_812),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_942),
.B(n_829),
.C(n_379),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_914),
.B(n_379),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_960),
.B(n_824),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_932),
.B(n_382),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_909),
.A2(n_1),
.B(n_2),
.C(n_7),
.Y(n_1085)
);

BUFx2_ASAP7_75t_SL g1086 ( 
.A(n_929),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_951),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_902),
.B(n_383),
.Y(n_1088)
);

AOI22x1_ASAP7_75t_L g1089 ( 
.A1(n_1025),
.A2(n_343),
.B1(n_312),
.B2(n_314),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_959),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_897),
.B(n_310),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_927),
.B(n_317),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_927),
.B(n_320),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_924),
.B(n_324),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_916),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_930),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_966),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_942),
.A2(n_345),
.B(n_328),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_948),
.A2(n_349),
.B1(n_329),
.B2(n_333),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_930),
.B(n_353),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_923),
.A2(n_687),
.B(n_668),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_904),
.B(n_1021),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1059),
.A2(n_93),
.B(n_185),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1011),
.A2(n_359),
.B1(n_358),
.B2(n_348),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_903),
.B(n_342),
.Y(n_1105)
);

BUFx8_ASAP7_75t_L g1106 ( 
.A(n_929),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_905),
.B(n_341),
.C(n_326),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_906),
.B(n_8),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_941),
.B(n_171),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_918),
.A2(n_14),
.B(n_19),
.C(n_20),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_917),
.A2(n_524),
.B1(n_22),
.B2(n_24),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_895),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1043),
.A2(n_161),
.B(n_148),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_SL g1114 ( 
.A(n_919),
.B(n_147),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1058),
.B(n_21),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_919),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1058),
.B(n_26),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_917),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1041),
.B(n_33),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_L g1120 ( 
.A(n_901),
.B(n_1005),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_SL g1121 ( 
.A(n_1030),
.B(n_37),
.C(n_39),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_958),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_903),
.B(n_920),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_910),
.B(n_118),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1020),
.Y(n_1125)
);

BUFx4f_ASAP7_75t_L g1126 ( 
.A(n_957),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1046),
.B(n_37),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_913),
.A2(n_39),
.B(n_41),
.C(n_43),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1053),
.B(n_44),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1017),
.A2(n_113),
.B(n_109),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1017),
.A2(n_104),
.B(n_100),
.Y(n_1131)
);

AND2x6_ASAP7_75t_SL g1132 ( 
.A(n_957),
.B(n_977),
.Y(n_1132)
);

BUFx5_ASAP7_75t_L g1133 ( 
.A(n_936),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_971),
.B(n_949),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1028),
.A2(n_97),
.B(n_95),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_949),
.B(n_44),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1028),
.A2(n_56),
.B(n_47),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1064),
.B(n_46),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_939),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1062),
.A2(n_55),
.B(n_49),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_948),
.A2(n_46),
.B(n_49),
.C(n_50),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_956),
.A2(n_53),
.B(n_55),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1010),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_1001),
.A2(n_1015),
.B1(n_965),
.B2(n_1051),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1054),
.A2(n_1055),
.B(n_1023),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1010),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_1007),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_997),
.B(n_989),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_956),
.A2(n_983),
.B(n_975),
.Y(n_1150)
);

INVx5_ASAP7_75t_L g1151 ( 
.A(n_936),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1036),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_997),
.B(n_989),
.Y(n_1153)
);

BUFx4f_ASAP7_75t_L g1154 ( 
.A(n_977),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1060),
.B(n_976),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1037),
.A2(n_1042),
.B(n_1009),
.C(n_1031),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_980),
.B(n_982),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_921),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_939),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_955),
.A2(n_1002),
.B(n_967),
.C(n_900),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1061),
.A2(n_940),
.B(n_945),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_911),
.A2(n_912),
.B(n_1049),
.C(n_1040),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_933),
.A2(n_1040),
.B1(n_940),
.B2(n_945),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_L g1164 ( 
.A(n_988),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_974),
.A2(n_983),
.B(n_975),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_978),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_986),
.B(n_1048),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_921),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_974),
.A2(n_1019),
.B(n_1056),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_926),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_SL g1171 ( 
.A1(n_1038),
.A2(n_1019),
.B(n_1063),
.C(n_1065),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_931),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1037),
.A2(n_1042),
.B1(n_1009),
.B2(n_908),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_933),
.A2(n_1038),
.B1(n_1016),
.B2(n_1035),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_979),
.A2(n_994),
.B(n_1004),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1036),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_953),
.A2(n_981),
.B1(n_1026),
.B2(n_935),
.Y(n_1177)
);

OAI22x1_ASAP7_75t_L g1178 ( 
.A1(n_1013),
.A2(n_987),
.B1(n_999),
.B2(n_996),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1054),
.A2(n_1052),
.B(n_1050),
.C(n_1035),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1027),
.C(n_970),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_947),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1023),
.A2(n_1055),
.B(n_1044),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_954),
.A2(n_962),
.B(n_961),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1057),
.Y(n_1184)
);

OA22x2_ASAP7_75t_L g1185 ( 
.A1(n_990),
.A2(n_1033),
.B1(n_998),
.B2(n_964),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_928),
.Y(n_1187)
);

AND3x1_ASAP7_75t_SL g1188 ( 
.A(n_1057),
.B(n_969),
.C(n_995),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1024),
.A2(n_938),
.B(n_963),
.C(n_937),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_928),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_953),
.B(n_950),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_934),
.B(n_972),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1047),
.A2(n_1039),
.B(n_1034),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1032),
.A2(n_1045),
.B(n_992),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_995),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_SL g1196 ( 
.A1(n_907),
.A2(n_915),
.B1(n_969),
.B2(n_985),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_934),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1003),
.A2(n_985),
.B(n_973),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1146),
.A2(n_992),
.B(n_915),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1079),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1122),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1192),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1066),
.B(n_1102),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1138),
.A2(n_936),
.B1(n_1029),
.B2(n_1022),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1116),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1175),
.A2(n_1045),
.B(n_946),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1067),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1073),
.B(n_907),
.C(n_1003),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1156),
.A2(n_1169),
.B(n_1198),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1074),
.A2(n_1045),
.B(n_943),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1078),
.B(n_943),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_SL g1212 ( 
.A(n_1151),
.B(n_1018),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1101),
.A2(n_946),
.B(n_991),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1095),
.B(n_1018),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1066),
.B(n_991),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1161),
.A2(n_1045),
.B(n_1018),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1158),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1070),
.A2(n_950),
.B(n_952),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1094),
.B(n_1104),
.C(n_1090),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1173),
.A2(n_1069),
.B(n_1071),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_SL g1221 ( 
.A(n_1098),
.B(n_1085),
.C(n_1099),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1178),
.A2(n_993),
.A3(n_1033),
.B(n_936),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1163),
.A2(n_993),
.B(n_1018),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1182),
.A2(n_1165),
.B(n_1150),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_1198),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1170),
.B(n_1172),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1181),
.B(n_1157),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1144),
.B(n_1088),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1068),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1134),
.B(n_1168),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1183),
.A2(n_1196),
.B(n_1194),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1167),
.B(n_1155),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1126),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1163),
.A2(n_1160),
.B(n_1092),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1179),
.A2(n_1189),
.A3(n_1145),
.B(n_1180),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1177),
.A2(n_1111),
.A3(n_1128),
.B(n_1137),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1193),
.A2(n_1076),
.B(n_1103),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1126),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1177),
.B(n_1075),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1112),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1113),
.A2(n_1093),
.B(n_1131),
.C(n_1135),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1111),
.A2(n_1118),
.A3(n_1141),
.B(n_1191),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1118),
.A2(n_1130),
.A3(n_1117),
.B(n_1115),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1143),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1075),
.A2(n_1171),
.B(n_1151),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1120),
.A2(n_1123),
.B(n_1080),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1162),
.A2(n_1083),
.B(n_1108),
.C(n_1119),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1087),
.B(n_1097),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1140),
.A2(n_1142),
.A3(n_1129),
.B(n_1127),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1151),
.A2(n_1114),
.B(n_1174),
.Y(n_1250)
);

AO32x2_ASAP7_75t_L g1251 ( 
.A1(n_1185),
.A2(n_1096),
.A3(n_1188),
.B1(n_1132),
.B2(n_1110),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1147),
.A2(n_1190),
.B(n_1187),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1106),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1164),
.B(n_1082),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1195),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1121),
.A2(n_1148),
.B(n_1084),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1184),
.B(n_1091),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1107),
.B(n_1081),
.C(n_1136),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1109),
.A2(n_1151),
.B(n_1185),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1186),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1106),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1116),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1149),
.B(n_1153),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1154),
.A2(n_1166),
.B1(n_1077),
.B2(n_1159),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1176),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1100),
.A2(n_1124),
.B(n_1159),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1125),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1152),
.B(n_1077),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1077),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1139),
.A2(n_1105),
.B(n_1133),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1086),
.B(n_1133),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1133),
.A2(n_1014),
.B(n_591),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1089),
.A2(n_1156),
.B(n_1073),
.C(n_751),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1133),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1066),
.B(n_781),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1106),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1156),
.A2(n_1178),
.A3(n_1179),
.B(n_1169),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1066),
.B(n_781),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1116),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1067),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1073),
.A2(n_751),
.B1(n_739),
.B2(n_750),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1175),
.A2(n_1014),
.B(n_591),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1156),
.A2(n_1169),
.B(n_1198),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1156),
.A2(n_1178),
.A3(n_1179),
.B(n_1169),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1156),
.A2(n_1169),
.B(n_1198),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_SL g1288 ( 
.A(n_1073),
.B(n_751),
.C(n_739),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_1113),
.B(n_1163),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1066),
.B(n_781),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1066),
.B(n_781),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1106),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1066),
.B(n_781),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1116),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1079),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1066),
.B(n_781),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1073),
.A2(n_751),
.B1(n_739),
.B2(n_750),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1066),
.B(n_781),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1066),
.B(n_781),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1156),
.A2(n_909),
.B(n_1173),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1156),
.A2(n_1073),
.B(n_751),
.C(n_1173),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1066),
.B(n_781),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1156),
.A2(n_1178),
.A3(n_1179),
.B(n_1169),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_R g1304 ( 
.A(n_1158),
.B(n_848),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1067),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1102),
.B(n_1000),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1146),
.A2(n_1101),
.B(n_1070),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1106),
.Y(n_1308)
);

AOI221xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1177),
.A2(n_751),
.B1(n_638),
.B2(n_909),
.C(n_1011),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1073),
.B(n_751),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1072),
.Y(n_1311)
);

AOI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1169),
.A2(n_923),
.B(n_1182),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1102),
.B(n_729),
.Y(n_1313)
);

NOR2x1_ASAP7_75t_SL g1314 ( 
.A(n_1151),
.B(n_919),
.Y(n_1314)
);

O2A1O1Ixp5_ASAP7_75t_L g1315 ( 
.A1(n_1113),
.A2(n_1093),
.B(n_1092),
.C(n_927),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1192),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1073),
.B(n_751),
.C(n_605),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1102),
.B(n_729),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1177),
.A2(n_751),
.B(n_1000),
.C(n_909),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1066),
.B(n_781),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1177),
.A2(n_751),
.B(n_1000),
.C(n_909),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1066),
.B(n_781),
.Y(n_1322)
);

AO32x2_ASAP7_75t_L g1323 ( 
.A1(n_1177),
.A2(n_1118),
.A3(n_1111),
.B1(n_1163),
.B2(n_1196),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1106),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1156),
.A2(n_1169),
.B(n_1198),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1156),
.A2(n_909),
.B(n_1180),
.C(n_1163),
.Y(n_1326)
);

AND2x6_ASAP7_75t_SL g1327 ( 
.A(n_1138),
.B(n_858),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1067),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1079),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1106),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1067),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1156),
.A2(n_1178),
.A3(n_1179),
.B(n_1169),
.Y(n_1332)
);

AND3x4_ASAP7_75t_L g1333 ( 
.A(n_1107),
.B(n_832),
.C(n_887),
.Y(n_1333)
);

AO32x2_ASAP7_75t_L g1334 ( 
.A1(n_1177),
.A2(n_1118),
.A3(n_1111),
.B1(n_1163),
.B2(n_1196),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1237),
.A2(n_1218),
.B(n_1307),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1259),
.B(n_1250),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1319),
.A2(n_1321),
.B(n_1271),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1310),
.A2(n_1317),
.B(n_1301),
.Y(n_1338)
);

INVx3_ASAP7_75t_SL g1339 ( 
.A(n_1278),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1220),
.A2(n_1231),
.B(n_1225),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1264),
.B(n_1233),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1300),
.A2(n_1297),
.B(n_1283),
.C(n_1309),
.Y(n_1342)
);

BUFx8_ASAP7_75t_SL g1343 ( 
.A(n_1253),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1264),
.B(n_1233),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1246),
.A2(n_1267),
.B(n_1223),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1213),
.A2(n_1224),
.B(n_1210),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1312),
.A2(n_1199),
.B(n_1284),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1288),
.A2(n_1289),
.B1(n_1219),
.B2(n_1221),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1274),
.A2(n_1315),
.B(n_1247),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1207),
.Y(n_1350)
);

OAI222xp33_ASAP7_75t_L g1351 ( 
.A1(n_1239),
.A2(n_1298),
.B1(n_1277),
.B2(n_1280),
.C1(n_1296),
.C2(n_1293),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1227),
.A2(n_1258),
.B(n_1226),
.C(n_1203),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1201),
.Y(n_1353)
);

BUFx4f_ASAP7_75t_L g1354 ( 
.A(n_1233),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1217),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1329),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1326),
.A2(n_1256),
.B1(n_1290),
.B2(n_1291),
.C(n_1299),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1208),
.A2(n_1322),
.B1(n_1320),
.B2(n_1302),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1230),
.B(n_1313),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1238),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1273),
.A2(n_1252),
.B(n_1276),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1209),
.A2(n_1325),
.B(n_1287),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1232),
.B(n_1228),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1209),
.A2(n_1285),
.B(n_1287),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1202),
.B(n_1316),
.Y(n_1365)
);

AND2x6_ASAP7_75t_L g1366 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1318),
.A2(n_1285),
.B1(n_1325),
.B2(n_1254),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1257),
.A2(n_1265),
.B(n_1269),
.C(n_1270),
.Y(n_1368)
);

OAI222xp33_ASAP7_75t_L g1369 ( 
.A1(n_1323),
.A2(n_1334),
.B1(n_1204),
.B2(n_1215),
.C1(n_1202),
.C2(n_1316),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1238),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1262),
.B(n_1272),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1268),
.A2(n_1214),
.B(n_1266),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1275),
.A2(n_1305),
.B(n_1331),
.C(n_1328),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1229),
.A2(n_1282),
.B(n_1311),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1205),
.A2(n_1281),
.B(n_1294),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1205),
.A2(n_1281),
.B(n_1294),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1200),
.B(n_1255),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1295),
.Y(n_1378)
);

AOI21xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1333),
.A2(n_1330),
.B(n_1292),
.Y(n_1379)
);

BUFx12f_ASAP7_75t_L g1380 ( 
.A(n_1324),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1279),
.A2(n_1286),
.B(n_1332),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1286),
.A2(n_1332),
.B(n_1303),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1286),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1304),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1263),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1211),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1327),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1303),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1235),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1308),
.B(n_1261),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1251),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1251),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1222),
.A2(n_1243),
.B(n_1249),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1323),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1323),
.A2(n_1334),
.B(n_1243),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1334),
.A2(n_1236),
.B1(n_1242),
.B2(n_1249),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1249),
.A2(n_1314),
.B(n_1236),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1242),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1212),
.B(n_1151),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1248),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1237),
.A2(n_1218),
.B(n_1307),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1237),
.A2(n_1218),
.B(n_1307),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1233),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1310),
.A2(n_1317),
.B1(n_1297),
.B2(n_1283),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1203),
.B(n_1306),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1248),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1231),
.A2(n_1245),
.B(n_1234),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1310),
.A2(n_751),
.B(n_1288),
.C(n_1317),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1310),
.A2(n_1317),
.B(n_1301),
.Y(n_1409)
);

OAI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1317),
.A2(n_1310),
.B1(n_751),
.B2(n_1297),
.C(n_1283),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_SL g1411 ( 
.A(n_1253),
.B(n_848),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1253),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1317),
.B(n_751),
.C(n_1310),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1317),
.B(n_751),
.C(n_1310),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1248),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1248),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1201),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1310),
.A2(n_1288),
.B1(n_1317),
.B2(n_1297),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1237),
.A2(n_1218),
.B(n_1307),
.Y(n_1419)
);

AO31x2_ASAP7_75t_L g1420 ( 
.A1(n_1289),
.A2(n_1231),
.A3(n_1225),
.B(n_1245),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1206),
.A2(n_1241),
.B(n_1216),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1253),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1310),
.B(n_1317),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1200),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1310),
.A2(n_1317),
.B(n_1301),
.Y(n_1425)
);

BUFx4f_ASAP7_75t_SL g1426 ( 
.A(n_1253),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1248),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1233),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1259),
.B(n_1250),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1260),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1310),
.A2(n_1288),
.B1(n_1317),
.B2(n_1297),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1310),
.A2(n_1321),
.B(n_1319),
.C(n_1301),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1248),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1310),
.A2(n_1288),
.B1(n_1317),
.B2(n_1297),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1310),
.A2(n_751),
.B1(n_1317),
.B2(n_1288),
.C(n_1319),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1310),
.A2(n_1288),
.B1(n_1317),
.B2(n_1297),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1304),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1206),
.A2(n_1241),
.B(n_1216),
.Y(n_1438)
);

AO31x2_ASAP7_75t_L g1439 ( 
.A1(n_1289),
.A2(n_1231),
.A3(n_1225),
.B(n_1245),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1317),
.A2(n_1310),
.B1(n_751),
.B2(n_1297),
.C(n_1283),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1310),
.A2(n_1288),
.B1(n_1297),
.B2(n_1283),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1310),
.A2(n_1317),
.B(n_1301),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1201),
.Y(n_1443)
);

OR3x4_ASAP7_75t_SL g1444 ( 
.A(n_1310),
.B(n_441),
.C(n_1255),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1237),
.A2(n_1218),
.B(n_1307),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1233),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1248),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1233),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1410),
.A2(n_1440),
.B1(n_1414),
.B2(n_1413),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1404),
.A2(n_1408),
.B(n_1432),
.Y(n_1450)
);

NOR2xp67_ASAP7_75t_L g1451 ( 
.A(n_1384),
.B(n_1437),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1441),
.A2(n_1431),
.B1(n_1436),
.B2(n_1434),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1377),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1432),
.A2(n_1352),
.B(n_1435),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1423),
.A2(n_1425),
.B(n_1442),
.C(n_1409),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1338),
.A2(n_1423),
.B(n_1342),
.C(n_1352),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1349),
.A2(n_1407),
.B(n_1336),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1407),
.A2(n_1429),
.B(n_1336),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1362),
.A2(n_1364),
.B(n_1393),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1365),
.B(n_1378),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1397),
.A2(n_1401),
.B(n_1335),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1418),
.A2(n_1431),
.B(n_1436),
.C(n_1434),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1355),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1343),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1443),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1399),
.A2(n_1336),
.B(n_1429),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1418),
.A2(n_1348),
.B1(n_1358),
.B2(n_1357),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1348),
.A2(n_1358),
.B1(n_1359),
.B2(n_1400),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1402),
.A2(n_1419),
.B(n_1445),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1341),
.B(n_1344),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1368),
.A2(n_1359),
.B(n_1447),
.C(n_1416),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1417),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1406),
.A2(n_1427),
.B(n_1433),
.C(n_1415),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1387),
.A2(n_1395),
.B1(n_1396),
.B2(n_1392),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1351),
.A2(n_1386),
.B(n_1444),
.C(n_1337),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1394),
.B(n_1391),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1424),
.B(n_1371),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1386),
.A2(n_1411),
.B1(n_1367),
.B2(n_1444),
.C(n_1430),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1395),
.A2(n_1396),
.B1(n_1350),
.B2(n_1340),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1395),
.A2(n_1367),
.B1(n_1354),
.B2(n_1353),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1354),
.A2(n_1385),
.B(n_1446),
.C(n_1370),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1379),
.A2(n_1356),
.B(n_1373),
.C(n_1345),
.Y(n_1482)
);

O2A1O1Ixp5_ASAP7_75t_L g1483 ( 
.A1(n_1369),
.A2(n_1398),
.B(n_1389),
.C(n_1388),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1403),
.B(n_1448),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1360),
.A2(n_1428),
.B(n_1390),
.C(n_1339),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1448),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1360),
.B(n_1372),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1420),
.B(n_1439),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1390),
.A2(n_1339),
.B(n_1388),
.C(n_1383),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1375),
.B(n_1376),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1426),
.A2(n_1422),
.B1(n_1380),
.B2(n_1412),
.Y(n_1492)
);

OA22x2_ASAP7_75t_L g1493 ( 
.A1(n_1361),
.A2(n_1347),
.B1(n_1366),
.B2(n_1346),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1420),
.B(n_1439),
.Y(n_1494)
);

CKINVDCx16_ASAP7_75t_R g1495 ( 
.A(n_1422),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1380),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1374),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1421),
.A2(n_1315),
.B(n_1241),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1410),
.A2(n_1310),
.B1(n_1283),
.B2(n_1297),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1374),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1410),
.A2(n_1440),
.B(n_1310),
.C(n_1408),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1410),
.A2(n_1440),
.B(n_1310),
.C(n_1408),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1410),
.A2(n_1310),
.B1(n_1283),
.B2(n_1297),
.Y(n_1503)
);

AOI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1410),
.A2(n_1310),
.B(n_1317),
.C(n_751),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1408),
.A2(n_1310),
.B(n_1317),
.C(n_1410),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1410),
.A2(n_1317),
.B1(n_1310),
.B2(n_1440),
.C(n_751),
.Y(n_1506)
);

AND2x2_ASAP7_75t_SL g1507 ( 
.A(n_1348),
.B(n_1418),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1408),
.A2(n_1310),
.B(n_1317),
.C(n_1410),
.Y(n_1508)
);

CKINVDCx6p67_ASAP7_75t_R g1509 ( 
.A(n_1339),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1349),
.A2(n_1438),
.B(n_1421),
.Y(n_1510)
);

O2A1O1Ixp5_ASAP7_75t_L g1511 ( 
.A1(n_1349),
.A2(n_1310),
.B(n_1289),
.C(n_1338),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1404),
.A2(n_1310),
.B1(n_1288),
.B2(n_1410),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1404),
.A2(n_1156),
.B(n_1301),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1363),
.B(n_1405),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1410),
.A2(n_1310),
.B1(n_1283),
.B2(n_1297),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1410),
.A2(n_1310),
.B1(n_1283),
.B2(n_1297),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1404),
.A2(n_1156),
.B(n_1301),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1421),
.A2(n_1315),
.B(n_1241),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1421),
.A2(n_1315),
.B(n_1241),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1366),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1410),
.A2(n_1310),
.B1(n_1283),
.B2(n_1297),
.Y(n_1521)
);

BUFx8_ASAP7_75t_SL g1522 ( 
.A(n_1464),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1510),
.B(n_1494),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1479),
.B(n_1488),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1498),
.A2(n_1519),
.B(n_1518),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1500),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1453),
.B(n_1455),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1490),
.B(n_1491),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1458),
.B(n_1457),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1499),
.A2(n_1515),
.B1(n_1516),
.B2(n_1521),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1459),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1459),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1496),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1476),
.B(n_1483),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1476),
.B(n_1474),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1474),
.B(n_1480),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1461),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1461),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1460),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1480),
.A2(n_1454),
.B(n_1450),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1493),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1469),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1520),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_SL g1545 ( 
.A1(n_1456),
.A2(n_1482),
.B(n_1475),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1487),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1466),
.B(n_1513),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1511),
.Y(n_1548)
);

AO21x2_ASAP7_75t_L g1549 ( 
.A1(n_1517),
.A2(n_1512),
.B(n_1467),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1473),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1468),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1468),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1471),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1467),
.A2(n_1508),
.B(n_1505),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1452),
.A2(n_1449),
.B(n_1503),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1477),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1489),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1507),
.Y(n_1558)
);

AO21x2_ASAP7_75t_L g1559 ( 
.A1(n_1452),
.A2(n_1449),
.B(n_1521),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1462),
.B(n_1502),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1515),
.A2(n_1501),
.B(n_1478),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1532),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1544),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1527),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1514),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1560),
.A2(n_1504),
.B1(n_1495),
.B2(n_1492),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1560),
.A2(n_1506),
.B1(n_1504),
.B2(n_1463),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1524),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1472),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1544),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1533),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1546),
.B(n_1470),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1546),
.B(n_1525),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1533),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1525),
.B(n_1529),
.Y(n_1577)
);

NAND4xp25_ASAP7_75t_L g1578 ( 
.A(n_1531),
.B(n_1485),
.C(n_1451),
.D(n_1481),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1556),
.B(n_1465),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1524),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1535),
.B(n_1486),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1526),
.B(n_1543),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1577),
.B(n_1542),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_L g1586 ( 
.A(n_1567),
.B(n_1553),
.C(n_1528),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1567),
.A2(n_1559),
.B1(n_1555),
.B2(n_1549),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1577),
.B(n_1542),
.Y(n_1588)
);

OAI211xp5_ASAP7_75t_L g1589 ( 
.A1(n_1568),
.A2(n_1531),
.B(n_1553),
.C(n_1528),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1567),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1578),
.B(n_1540),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1568),
.A2(n_1545),
.B1(n_1554),
.B2(n_1559),
.C(n_1555),
.Y(n_1592)
);

NAND4xp25_ASAP7_75t_L g1593 ( 
.A(n_1578),
.B(n_1552),
.C(n_1551),
.D(n_1558),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1570),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1563),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1570),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1564),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1580),
.Y(n_1598)
);

AO21x1_ASAP7_75t_SL g1599 ( 
.A1(n_1582),
.A2(n_1537),
.B(n_1557),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1575),
.B(n_1537),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1571),
.B(n_1540),
.Y(n_1601)
);

AND4x1_ASAP7_75t_L g1602 ( 
.A(n_1581),
.B(n_1552),
.C(n_1551),
.D(n_1554),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1584),
.A2(n_1539),
.B(n_1538),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1578),
.A2(n_1559),
.B1(n_1555),
.B2(n_1549),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1563),
.Y(n_1605)
);

AND2x4_ASAP7_75t_SL g1606 ( 
.A(n_1572),
.B(n_1544),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1563),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1565),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1572),
.A2(n_1560),
.B1(n_1547),
.B2(n_1558),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1556),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1566),
.B(n_1560),
.C(n_1548),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1579),
.A2(n_1545),
.B1(n_1554),
.B2(n_1555),
.C(n_1559),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1575),
.B(n_1542),
.Y(n_1613)
);

BUFx10_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1583),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1579),
.A2(n_1555),
.B(n_1541),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1536),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1583),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1615),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1603),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1595),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1602),
.A2(n_1573),
.B(n_1562),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1614),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1614),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1594),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1602),
.A2(n_1573),
.B(n_1562),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1530),
.Y(n_1627)
);

OR2x6_ASAP7_75t_L g1628 ( 
.A(n_1611),
.B(n_1530),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1615),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1595),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1611),
.A2(n_1569),
.B(n_1576),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1596),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1605),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1618),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1591),
.B(n_1554),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1607),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1618),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1592),
.B(n_1544),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1608),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1608),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1612),
.B(n_1544),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1635),
.B(n_1604),
.C(n_1586),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1635),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1560),
.C(n_1587),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1634),
.B(n_1606),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1634),
.B(n_1599),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1625),
.B(n_1600),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1625),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1634),
.B(n_1599),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1641),
.Y(n_1651)
);

NAND4xp25_ASAP7_75t_L g1652 ( 
.A(n_1642),
.B(n_1593),
.C(n_1589),
.D(n_1548),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1632),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1585),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1622),
.B(n_1585),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1632),
.B(n_1600),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1641),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1622),
.B(n_1588),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1620),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1642),
.B(n_1617),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1622),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1622),
.B(n_1588),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1621),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1619),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1621),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1622),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1627),
.A2(n_1590),
.B(n_1593),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_SL g1670 ( 
.A1(n_1626),
.A2(n_1572),
.B(n_1601),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1620),
.Y(n_1671)
);

OAI31xp33_ASAP7_75t_L g1672 ( 
.A1(n_1619),
.A2(n_1609),
.A3(n_1550),
.B(n_1590),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1620),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1637),
.B(n_1617),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1626),
.B(n_1623),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1626),
.B(n_1597),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1626),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1628),
.A2(n_1541),
.B1(n_1549),
.B2(n_1561),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1631),
.Y(n_1680)
);

NAND2x1_ASAP7_75t_L g1681 ( 
.A(n_1623),
.B(n_1624),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1649),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1660),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1660),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1648),
.B(n_1629),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1643),
.B(n_1629),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1643),
.B(n_1638),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1666),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1666),
.Y(n_1690)
);

AOI311xp33_ASAP7_75t_L g1691 ( 
.A1(n_1669),
.A2(n_1636),
.A3(n_1630),
.B(n_1640),
.C(n_1633),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_1638),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1646),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1647),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1630),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1623),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1665),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1623),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1646),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1650),
.B(n_1623),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1646),
.B(n_1623),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1667),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1652),
.B(n_1613),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1651),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1651),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_SL g1709 ( 
.A(n_1672),
.B(n_1572),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1657),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1657),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1656),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1659),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1646),
.B(n_1624),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1654),
.B(n_1624),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1654),
.B(n_1624),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1685),
.B(n_1674),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1685),
.B(n_1661),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1692),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1688),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1683),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1713),
.B(n_1676),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1689),
.B(n_1677),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1688),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1699),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1709),
.A2(n_1645),
.B1(n_1687),
.B2(n_1686),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1693),
.B(n_1677),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1699),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1696),
.B(n_1655),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1698),
.A2(n_1645),
.B1(n_1679),
.B2(n_1668),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1690),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1690),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1696),
.B(n_1655),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1716),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1658),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1658),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_1682),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1683),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1697),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1694),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1715),
.B(n_1664),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1697),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1742),
.B(n_1713),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1733),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1728),
.A2(n_1541),
.B1(n_1549),
.B2(n_1627),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1724),
.B(n_1715),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1724),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1732),
.A2(n_1707),
.B1(n_1711),
.B2(n_1708),
.C(n_1712),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1732),
.A2(n_1720),
.B1(n_1742),
.B2(n_1724),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1739),
.A2(n_1691),
.B(n_1672),
.C(n_1662),
.Y(n_1752)
);

AOI32xp33_ASAP7_75t_L g1753 ( 
.A1(n_1721),
.A2(n_1726),
.A3(n_1739),
.B1(n_1725),
.B2(n_1727),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1722),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1705),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1730),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1719),
.A2(n_1541),
.B1(n_1627),
.B2(n_1628),
.Y(n_1757)
);

AOI222xp33_ASAP7_75t_L g1758 ( 
.A1(n_1721),
.A2(n_1726),
.B1(n_1662),
.B2(n_1668),
.C1(n_1725),
.C2(n_1734),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1734),
.A2(n_1744),
.B1(n_1722),
.B2(n_1741),
.C(n_1740),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1718),
.A2(n_1627),
.B1(n_1628),
.B2(n_1675),
.C(n_1681),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1718),
.B(n_1522),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1719),
.A2(n_1541),
.B1(n_1627),
.B2(n_1628),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1740),
.Y(n_1763)
);

OAI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1730),
.A2(n_1627),
.B1(n_1628),
.B2(n_1675),
.C(n_1681),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1729),
.B(n_1703),
.Y(n_1765)
);

NAND2x1_ASAP7_75t_L g1766 ( 
.A(n_1765),
.B(n_1703),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1753),
.B(n_1734),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1749),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1761),
.B(n_1522),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1756),
.B(n_1736),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1745),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1746),
.B(n_1736),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1748),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1755),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1751),
.B(n_1496),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1758),
.B(n_1736),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1754),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1775),
.A2(n_1747),
.B(n_1750),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1773),
.Y(n_1779)
);

OAI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1767),
.A2(n_1750),
.B1(n_1752),
.B2(n_1757),
.C(n_1762),
.Y(n_1780)
);

AOI321xp33_ASAP7_75t_L g1781 ( 
.A1(n_1776),
.A2(n_1759),
.A3(n_1760),
.B1(n_1764),
.B2(n_1763),
.C(n_1729),
.Y(n_1781)
);

AOI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1771),
.A2(n_1759),
.B(n_1741),
.C(n_1744),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1770),
.B(n_1703),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1770),
.A2(n_1496),
.B(n_1723),
.Y(n_1784)
);

OAI211xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1774),
.A2(n_1723),
.B(n_1678),
.C(n_1714),
.Y(n_1785)
);

AOI21xp33_ASAP7_75t_L g1786 ( 
.A1(n_1766),
.A2(n_1702),
.B(n_1684),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1772),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1777),
.A2(n_1670),
.B(n_1678),
.C(n_1627),
.Y(n_1788)
);

O2A1O1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1780),
.A2(n_1782),
.B(n_1778),
.C(n_1779),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1784),
.A2(n_1769),
.B(n_1768),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1783),
.Y(n_1791)
);

NOR2x1p5_ASAP7_75t_L g1792 ( 
.A(n_1787),
.B(n_1509),
.Y(n_1792)
);

AOI22x1_ASAP7_75t_L g1793 ( 
.A1(n_1781),
.A2(n_1670),
.B1(n_1534),
.B2(n_1678),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1786),
.B(n_1743),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1785),
.Y(n_1795)
);

AOI211x1_ASAP7_75t_L g1796 ( 
.A1(n_1788),
.A2(n_1704),
.B(n_1706),
.C(n_1737),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1791),
.B(n_1743),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1792),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1794),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_L g1800 ( 
.A(n_1793),
.B(n_1731),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1795),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1790),
.B(n_1731),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1796),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1789),
.B(n_1706),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1797),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1804),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1802),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1804),
.Y(n_1808)
);

OAI322xp33_ASAP7_75t_L g1809 ( 
.A1(n_1803),
.A2(n_1678),
.A3(n_1680),
.B1(n_1714),
.B2(n_1738),
.C1(n_1737),
.C2(n_1735),
.Y(n_1809)
);

INVx5_ASAP7_75t_L g1810 ( 
.A(n_1806),
.Y(n_1810)
);

INVx3_ASAP7_75t_SL g1811 ( 
.A(n_1805),
.Y(n_1811)
);

NOR3xp33_ASAP7_75t_L g1812 ( 
.A(n_1807),
.B(n_1799),
.C(n_1798),
.Y(n_1812)
);

NAND4xp75_ASAP7_75t_L g1813 ( 
.A(n_1811),
.B(n_1801),
.C(n_1808),
.D(n_1806),
.Y(n_1813)
);

AOI322xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1812),
.A3(n_1800),
.B1(n_1810),
.B2(n_1735),
.C1(n_1738),
.C2(n_1680),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1814),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1814),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1815),
.A2(n_1534),
.B1(n_1809),
.B2(n_1695),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1816),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1818),
.A2(n_1695),
.B1(n_1710),
.B2(n_1716),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1817),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1820),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1819),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1680),
.B1(n_1671),
.B2(n_1673),
.C1(n_1663),
.C2(n_1659),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1823),
.A2(n_1717),
.B1(n_1680),
.B2(n_1664),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1717),
.B1(n_1659),
.B2(n_1673),
.Y(n_1825)
);

AOI211xp5_ASAP7_75t_L g1826 ( 
.A1(n_1825),
.A2(n_1663),
.B(n_1671),
.C(n_1673),
.Y(n_1826)
);


endmodule