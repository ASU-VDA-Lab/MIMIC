module fake_jpeg_21495_n_297 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_121;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_50),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_19),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_22),
.B1(n_25),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_59),
.B1(n_66),
.B2(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_51),
.B1(n_32),
.B2(n_43),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_20),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_34),
.B1(n_38),
.B2(n_0),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_18),
.C(n_30),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_33),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_80),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_33),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_28),
.B(n_19),
.C(n_36),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_28),
.B1(n_36),
.B2(n_35),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_86),
.B1(n_0),
.B2(n_1),
.Y(n_88)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_6),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_87),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_31),
.B1(n_27),
.B2(n_38),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_34),
.B1(n_8),
.B2(n_2),
.Y(n_87)
);

AO21x1_ASAP7_75t_SL g149 ( 
.A1(n_88),
.A2(n_110),
.B(n_113),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_3),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_103),
.C(n_54),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_93),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_3),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_111),
.B1(n_122),
.B2(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_105),
.Y(n_142)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_6),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_73),
.Y(n_109)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_7),
.Y(n_111)
);

OR2x4_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_15),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_65),
.B(n_7),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_70),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_8),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_66),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_70),
.A2(n_66),
.B1(n_68),
.B2(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_92),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_76),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_145),
.B(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_53),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_150),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_103),
.C(n_90),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_153),
.C(n_103),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_53),
.B1(n_79),
.B2(n_78),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_114),
.B1(n_96),
.B2(n_92),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_147),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_74),
.B1(n_57),
.B2(n_52),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_148),
.B1(n_116),
.B2(n_110),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_68),
.B1(n_74),
.B2(n_57),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_70),
.B1(n_83),
.B2(n_11),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_9),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_9),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_10),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_9),
.C(n_10),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_161),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_167),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_109),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_162),
.B1(n_178),
.B2(n_179),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_120),
.B1(n_97),
.B2(n_113),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_149),
.B(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_95),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_168),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_94),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_105),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_117),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_129),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_171),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_104),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_117),
.B1(n_114),
.B2(n_99),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_115),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_183),
.B(n_184),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_126),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_124),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_190),
.B(n_203),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_148),
.B1(n_134),
.B2(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_193),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_134),
.B(n_127),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_210),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_145),
.B1(n_141),
.B2(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_146),
.B1(n_129),
.B2(n_124),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_194),
.A2(n_199),
.B1(n_173),
.B2(n_164),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_129),
.B1(n_152),
.B2(n_153),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_154),
.B(n_167),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_140),
.B(n_100),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_92),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_152),
.B1(n_12),
.B2(n_13),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_177),
.B(n_188),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_158),
.C(n_166),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_162),
.C(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_157),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_225),
.B1(n_189),
.B2(n_194),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_159),
.B1(n_164),
.B2(n_178),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_176),
.C(n_183),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_185),
.B(n_156),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_196),
.A3(n_190),
.B1(n_186),
.B2(n_210),
.C1(n_171),
.C2(n_197),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_179),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_182),
.Y(n_246)
);

BUFx12f_ASAP7_75t_SL g230 ( 
.A(n_203),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_202),
.B(n_187),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_207),
.B1(n_195),
.B2(n_196),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_247),
.B(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_235),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_200),
.B1(n_202),
.B2(n_208),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_244),
.B1(n_223),
.B2(n_215),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_193),
.B1(n_187),
.B2(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_192),
.B1(n_195),
.B2(n_185),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_226),
.B(n_214),
.C(n_230),
.D(n_227),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_197),
.B1(n_188),
.B2(n_186),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_229),
.Y(n_249)
);

AOI21x1_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_255),
.B(n_256),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_260),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_218),
.C(n_212),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_261),
.C(n_244),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_256),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_252),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_222),
.B(n_215),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_222),
.B(n_220),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_245),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_247),
.B1(n_216),
.B2(n_217),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_242),
.B1(n_235),
.B2(n_198),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_219),
.B1(n_214),
.B2(n_198),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_239),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_182),
.C(n_160),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_242),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_269),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_259),
.B1(n_254),
.B2(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_276),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_261),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_255),
.B(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_279),
.C(n_249),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.C(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_264),
.B(n_248),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_252),
.B(n_251),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_278),
.C(n_160),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_288),
.A3(n_125),
.B1(n_92),
.B2(n_121),
.C1(n_101),
.C2(n_15),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_278),
.B1(n_13),
.B2(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_121),
.C(n_125),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_121),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_293),
.B(n_121),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_10),
.Y(n_297)
);


endmodule