module fake_ibex_977_n_1683 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_314, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1683);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1683;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1614;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_655;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_650;
wire n_409;
wire n_1575;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_633;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_1657;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1460;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_339;
wire n_348;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1673;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1586;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_336;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_416;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

BUFx2_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_265),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_30),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_288),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_37),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_43),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_215),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_50),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_177),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_61),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_128),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_142),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_293),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_0),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_237),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_94),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_130),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_68),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_99),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_38),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_229),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_28),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_217),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_234),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_274),
.Y(n_358)
);

BUFx8_ASAP7_75t_SL g359 ( 
.A(n_8),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_135),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_230),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_232),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_65),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_227),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_186),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_55),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_259),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_283),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_147),
.B(n_225),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_163),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_136),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_277),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_187),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_79),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_160),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_158),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_49),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_270),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_204),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_2),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_134),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_49),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_11),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_320),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_257),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_128),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_241),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_143),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_285),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_102),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_243),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_89),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_198),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_250),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_79),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_180),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_151),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_275),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_50),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_84),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_55),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_284),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_171),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_16),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_261),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_143),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_195),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_239),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_58),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_252),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_210),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_255),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_242),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_228),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_221),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_268),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_149),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_59),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_130),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_182),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_297),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_256),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_14),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_299),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_87),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_200),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_193),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_38),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_88),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_148),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_207),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_40),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_86),
.Y(n_437)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_23),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_319),
.B(n_167),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_51),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_310),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_123),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_32),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_223),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_137),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_175),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_24),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_294),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_119),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_240),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_18),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_273),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_63),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_214),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_1),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_258),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_315),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_303),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_220),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_100),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_216),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_62),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_291),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_311),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_281),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_205),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_262),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_235),
.Y(n_468)
);

BUFx8_ASAP7_75t_SL g469 ( 
.A(n_326),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_153),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_88),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_112),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_172),
.B(n_149),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_323),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_321),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_26),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_146),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_158),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_142),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_280),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_164),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_224),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_45),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_226),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_12),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_178),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_140),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_251),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_9),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_129),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_107),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_95),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_131),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_67),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_278),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_68),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_271),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_30),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_213),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_18),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_48),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_231),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_173),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_181),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_22),
.Y(n_505)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_290),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_309),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_124),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_292),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_132),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_21),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_276),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_145),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_263),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_306),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_146),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_286),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_192),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_318),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_313),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_21),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_24),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_138),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_245),
.B(n_46),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_87),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_282),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_102),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_15),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_156),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_42),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_194),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_63),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_127),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_222),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_59),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_44),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_131),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_219),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_244),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_150),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_179),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_212),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_260),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_90),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_236),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_108),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g547 ( 
.A(n_308),
.B(n_116),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_96),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_170),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_279),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_165),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_287),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_209),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_266),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_156),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_189),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_134),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_111),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_155),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_46),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_13),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_314),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_317),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_6),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_415),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_415),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_510),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_327),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_469),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_339),
.B(n_1),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_438),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_438),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_406),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_438),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_415),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_331),
.B(n_166),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_437),
.B(n_3),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_415),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_438),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_339),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_354),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_586)
);

AOI22x1_ASAP7_75t_SL g587 ( 
.A1(n_451),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_354),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_588)
);

NOR2x1_ASAP7_75t_L g589 ( 
.A(n_360),
.B(n_168),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_331),
.B(n_358),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_379),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_360),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_469),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_417),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_332),
.B(n_7),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_381),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_359),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_381),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_417),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_417),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_351),
.B(n_10),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_417),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_407),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_426),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_379),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_440),
.B(n_11),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_494),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_426),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_564),
.B(n_12),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_358),
.Y(n_610)
);

OA21x2_ASAP7_75t_L g611 ( 
.A1(n_391),
.A2(n_176),
.B(n_174),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_426),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_426),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_564),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_391),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_338),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_371),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_338),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_522),
.B(n_13),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_396),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_329),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_396),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_397),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_328),
.B(n_183),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_517),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_531),
.Y(n_629)
);

OA21x2_ASAP7_75t_L g630 ( 
.A1(n_397),
.A2(n_185),
.B(n_184),
.Y(n_630)
);

OA21x2_ASAP7_75t_L g631 ( 
.A1(n_424),
.A2(n_190),
.B(n_188),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_368),
.B(n_14),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_491),
.B(n_15),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_340),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_359),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_353),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_487),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_341),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_368),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_347),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_505),
.B(n_17),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_345),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_372),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_347),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_372),
.B(n_19),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_377),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_349),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_531),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_531),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_424),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_431),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_350),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_352),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_400),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_373),
.B(n_20),
.Y(n_656)
);

CKINVDCx16_ASAP7_75t_R g657 ( 
.A(n_361),
.Y(n_657)
);

NOR2x1_ASAP7_75t_L g658 ( 
.A(n_363),
.B(n_191),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_566),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_566),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_569),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_609),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_609),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_569),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_571),
.B(n_343),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_640),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_574),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_568),
.B(n_619),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_609),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_644),
.B(n_654),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_575),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_575),
.Y(n_674)
);

NOR2x1p5_ASAP7_75t_L g675 ( 
.A(n_570),
.B(n_508),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_632),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_622),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_646),
.B(n_486),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_577),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_578),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_607),
.B(n_373),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_622),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_656),
.A2(n_366),
.B1(n_378),
.B2(n_370),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_583),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_572),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_584),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_604),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_604),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_604),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_646),
.B(n_488),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_604),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_567),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_632),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_645),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_657),
.B(n_506),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_645),
.B(n_446),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_572),
.B(n_399),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_610),
.B(n_541),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_585),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_585),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_655),
.B(n_502),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_570),
.A2(n_487),
.B1(n_513),
.B2(n_511),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_636),
.A2(n_419),
.B1(n_463),
.B2(n_399),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_610),
.B(n_513),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_639),
.Y(n_709)
);

NOR2x1p5_ASAP7_75t_L g710 ( 
.A(n_576),
.B(n_516),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_591),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_624),
.B(n_516),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_582),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_634),
.B(n_384),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_582),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_639),
.B(n_521),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_593),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_643),
.B(n_541),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_636),
.B(n_506),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_591),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_605),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_643),
.B(n_334),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_580),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_658),
.B(n_336),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_589),
.B(n_342),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_582),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_576),
.B(n_346),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_617),
.B(n_348),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_617),
.Y(n_730)
);

BUFx4f_ASAP7_75t_L g731 ( 
.A(n_580),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_623),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_595),
.B(n_523),
.C(n_521),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_580),
.B(n_563),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

AND2x2_ASAP7_75t_SL g736 ( 
.A(n_627),
.B(n_473),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_625),
.B(n_355),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

INVxp67_ASAP7_75t_SL g739 ( 
.A(n_601),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_638),
.B(n_530),
.C(n_523),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_594),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_581),
.B(n_385),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_594),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_586),
.A2(n_548),
.B1(n_530),
.B2(n_451),
.Y(n_745)
);

NOR2x1p5_ASAP7_75t_L g746 ( 
.A(n_593),
.B(n_548),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_625),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_626),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_581),
.B(n_533),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_626),
.B(n_356),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_650),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_599),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_642),
.B(n_357),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_647),
.B(n_337),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_650),
.B(n_365),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_599),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_599),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_651),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_652),
.B(n_337),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_651),
.B(n_367),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_653),
.B(n_382),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_592),
.B(n_344),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_565),
.B(n_389),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_606),
.B(n_641),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_633),
.A2(n_463),
.B1(n_464),
.B2(n_419),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_599),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_599),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_600),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_565),
.B(n_392),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_600),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_600),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_606),
.B(n_376),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_602),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_602),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_602),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_602),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_641),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_596),
.B(n_394),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_573),
.B(n_335),
.C(n_333),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_592),
.B(n_344),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_597),
.B(n_533),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_608),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_592),
.B(n_388),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_611),
.A2(n_408),
.B(n_405),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_603),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_590),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_598),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_597),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_615),
.B(n_362),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_615),
.B(n_362),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_608),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_565),
.B(n_410),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_573),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_618),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_612),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_612),
.Y(n_797)
);

NOR2x1p5_ASAP7_75t_L g798 ( 
.A(n_635),
.B(n_402),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_611),
.B(n_338),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_612),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_580),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_612),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_618),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_612),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_613),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_613),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_621),
.B(n_423),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_613),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_635),
.B(n_649),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_649),
.B(n_411),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_588),
.B(n_377),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_668),
.B(n_533),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_662),
.A2(n_412),
.B(n_420),
.C(n_403),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_739),
.B(n_515),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_811),
.A2(n_427),
.B1(n_429),
.B2(n_422),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_755),
.B(n_515),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_789),
.Y(n_817)
);

INVx8_ASAP7_75t_L g818 ( 
.A(n_742),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_784),
.Y(n_819)
);

BUFx5_ASAP7_75t_L g820 ( 
.A(n_801),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_SL g821 ( 
.A1(n_707),
.A2(n_500),
.B1(n_637),
.B2(n_550),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_676),
.B(n_678),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_683),
.B(n_518),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_766),
.B(n_433),
.C(n_421),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_811),
.A2(n_765),
.B1(n_736),
.B2(n_696),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_750),
.A2(n_550),
.B1(n_464),
.B2(n_375),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_714),
.B(n_794),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_773),
.B(n_672),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_697),
.B(n_677),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_784),
.Y(n_830)
);

BUFx8_ASAP7_75t_L g831 ( 
.A(n_698),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_705),
.B(n_534),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_745),
.B(n_383),
.C(n_374),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_760),
.B(n_538),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_784),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_788),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_679),
.B(n_538),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_L g838 ( 
.A(n_706),
.B(n_545),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_691),
.B(n_549),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_708),
.B(n_549),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_716),
.B(n_551),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_811),
.A2(n_434),
.B1(n_442),
.B2(n_432),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_724),
.B(n_551),
.Y(n_843)
);

AO22x2_ASAP7_75t_L g844 ( 
.A1(n_778),
.A2(n_587),
.B1(n_500),
.B2(n_449),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_732),
.Y(n_845)
);

BUFx6f_ASAP7_75t_SL g846 ( 
.A(n_811),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_330),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_L g848 ( 
.A(n_740),
.B(n_393),
.C(n_390),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_712),
.B(n_398),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_732),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_786),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_811),
.A2(n_409),
.B1(n_436),
.B2(n_404),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_733),
.B(n_22),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_763),
.B(n_364),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_687),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_445),
.C(n_443),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_732),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_781),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_663),
.B(n_611),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_736),
.A2(n_462),
.B1(n_470),
.B2(n_447),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_759),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_671),
.B(n_699),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_702),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_801),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_699),
.B(n_630),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_720),
.B(n_386),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_665),
.B(n_435),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_670),
.B(n_444),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_709),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_703),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_790),
.B(n_380),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_791),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_789),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_728),
.B(n_782),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_754),
.B(n_630),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_798),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_742),
.B(n_471),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_742),
.B(n_456),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_667),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_762),
.B(n_630),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_762),
.B(n_631),
.Y(n_881)
);

INVx8_ASAP7_75t_L g882 ( 
.A(n_742),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_659),
.B(n_660),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_746),
.B(n_717),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_711),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_721),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_722),
.Y(n_887)
);

BUFx8_ASAP7_75t_L g888 ( 
.A(n_811),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_730),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_780),
.A2(n_477),
.B1(n_479),
.B2(n_476),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_684),
.A2(n_483),
.B1(n_485),
.B2(n_481),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_675),
.Y(n_892)
);

O2A1O1Ixp5_ASAP7_75t_L g893 ( 
.A1(n_723),
.A2(n_725),
.B(n_726),
.C(n_785),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_747),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_725),
.B(n_539),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_749),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_752),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_700),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_667),
.B(n_413),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_723),
.B(n_428),
.Y(n_900)
);

CKINVDCx11_ASAP7_75t_R g901 ( 
.A(n_686),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_809),
.B(n_542),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_710),
.B(n_492),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_704),
.B(n_430),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_659),
.B(n_631),
.Y(n_905)
);

BUFx8_ASAP7_75t_L g906 ( 
.A(n_717),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_779),
.B(n_453),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_701),
.A2(n_460),
.B1(n_472),
.B2(n_455),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_729),
.A2(n_498),
.B1(n_525),
.B2(n_493),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_660),
.B(n_631),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_807),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_661),
.B(n_414),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_726),
.B(n_529),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_661),
.B(n_416),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_737),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_701),
.B(n_452),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_787),
.B(n_458),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_751),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_756),
.B(n_761),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_761),
.A2(n_536),
.B1(n_537),
.B2(n_532),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_719),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_734),
.A2(n_544),
.B(n_546),
.C(n_540),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_664),
.B(n_418),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_666),
.B(n_425),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_799),
.A2(n_561),
.B1(n_557),
.B2(n_478),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_764),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_669),
.B(n_466),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_L g928 ( 
.A(n_795),
.B(n_803),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_673),
.B(n_448),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_764),
.B(n_770),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_674),
.B(n_450),
.Y(n_931)
);

BUFx5_ASAP7_75t_L g932 ( 
.A(n_799),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_770),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_680),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_680),
.B(n_480),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_681),
.B(n_482),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_734),
.A2(n_490),
.B1(n_496),
.B2(n_489),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_793),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_685),
.B(n_454),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_810),
.A2(n_555),
.B1(n_558),
.B2(n_501),
.Y(n_940)
);

O2A1O1Ixp5_ASAP7_75t_L g941 ( 
.A1(n_693),
.A2(n_459),
.B(n_461),
.C(n_457),
.Y(n_941)
);

INVx8_ASAP7_75t_L g942 ( 
.A(n_743),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_SL g943 ( 
.A(n_743),
.B(n_560),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_688),
.B(n_524),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_743),
.B(n_553),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_688),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_689),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_690),
.A2(n_395),
.B1(n_527),
.B2(n_338),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_692),
.B(n_369),
.C(n_465),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_693),
.A2(n_395),
.B1(n_535),
.B2(n_527),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_743),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_694),
.Y(n_952)
);

NOR2x1p5_ASAP7_75t_L g953 ( 
.A(n_694),
.B(n_387),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_772),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_695),
.A2(n_395),
.B1(n_535),
.B2(n_527),
.Y(n_955)
);

AO22x2_ASAP7_75t_L g956 ( 
.A1(n_695),
.A2(n_468),
.B1(n_474),
.B2(n_467),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_783),
.B(n_475),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_713),
.Y(n_958)
);

O2A1O1Ixp5_ASAP7_75t_L g959 ( 
.A1(n_715),
.A2(n_497),
.B(n_499),
.C(n_495),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_808),
.B(n_503),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_718),
.B(n_395),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_783),
.B(n_507),
.Y(n_962)
);

AND2x6_ASAP7_75t_L g963 ( 
.A(n_718),
.B(n_387),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_727),
.B(n_509),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_727),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_735),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_783),
.B(n_512),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_738),
.A2(n_519),
.B1(n_520),
.B2(n_514),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_738),
.B(n_526),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_741),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_744),
.B(n_547),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_748),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_800),
.B(n_543),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_753),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_757),
.B(n_552),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_758),
.A2(n_535),
.B1(n_559),
.B2(n_527),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_L g977 ( 
.A(n_767),
.B(n_23),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_L g978 ( 
.A(n_767),
.B(n_556),
.C(n_554),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_768),
.Y(n_979)
);

AND2x6_ASAP7_75t_SL g980 ( 
.A(n_802),
.B(n_562),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_828),
.B(n_535),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_818),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_818),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_859),
.A2(n_865),
.B(n_875),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_814),
.B(n_439),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_818),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_819),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_860),
.A2(n_441),
.B1(n_504),
.B2(n_401),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_882),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_880),
.A2(n_771),
.B(n_769),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_874),
.B(n_25),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_870),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_812),
.B(n_25),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_906),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_905),
.A2(n_775),
.B(n_774),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_910),
.A2(n_776),
.B(n_775),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_910),
.A2(n_777),
.B(n_776),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_830),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_L g999 ( 
.A(n_824),
.B(n_563),
.C(n_649),
.Y(n_999)
);

OA22x2_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_881),
.A2(n_822),
.B(n_829),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_882),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_911),
.B(n_31),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_826),
.B(n_849),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_898),
.B(n_31),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_878),
.B(n_32),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_893),
.A2(n_796),
.B(n_792),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_822),
.A2(n_804),
.B(n_797),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_882),
.A2(n_579),
.B1(n_649),
.B2(n_616),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_827),
.A2(n_862),
.B(n_883),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_827),
.A2(n_806),
.B(n_805),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_925),
.A2(n_806),
.B(n_35),
.C(n_33),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_813),
.A2(n_616),
.B(n_620),
.C(n_614),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_858),
.B(n_34),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_L g1015 ( 
.A(n_833),
.B(n_34),
.C(n_35),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_872),
.B(n_36),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_877),
.B(n_36),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_823),
.B(n_37),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_835),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_869),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_855),
.A2(n_628),
.B(n_629),
.C(n_620),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_877),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_941),
.A2(n_629),
.B(n_628),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_817),
.B(n_873),
.Y(n_1024)
);

OAI22x1_ASAP7_75t_L g1025 ( 
.A1(n_852),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_868),
.B(n_913),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_913),
.B(n_39),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_851),
.B(n_42),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_832),
.B(n_43),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_879),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_876),
.B(n_45),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_922),
.A2(n_648),
.B(n_51),
.C(n_47),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_843),
.A2(n_834),
.B(n_816),
.Y(n_1033)
);

O2A1O1Ixp5_ASAP7_75t_L g1034 ( 
.A1(n_959),
.A2(n_197),
.B(n_199),
.C(n_196),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_837),
.A2(n_202),
.B(n_201),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_937),
.B(n_48),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_839),
.A2(n_841),
.B(n_840),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_847),
.B(n_52),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_907),
.B(n_52),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_934),
.A2(n_206),
.B(n_203),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_825),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_901),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_854),
.B(n_54),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_863),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_871),
.B(n_57),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_SL g1046 ( 
.A1(n_967),
.A2(n_218),
.B(n_325),
.C(n_324),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_927),
.A2(n_211),
.B(n_208),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_815),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_885),
.A2(n_60),
.B(n_64),
.C(n_65),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_838),
.B(n_866),
.Y(n_1050)
);

AOI33xp33_ASAP7_75t_L g1051 ( 
.A1(n_842),
.A2(n_66),
.A3(n_67),
.B1(n_69),
.B2(n_70),
.B3(n_71),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_867),
.B(n_66),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_846),
.A2(n_919),
.B1(n_956),
.B2(n_896),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_886),
.B(n_69),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_887),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_903),
.B(n_70),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_892),
.B(n_72),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_889),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_894),
.B(n_73),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_897),
.B(n_74),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_895),
.B(n_74),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_906),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_956),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_890),
.B(n_75),
.Y(n_1064)
);

OAI321xp33_ASAP7_75t_L g1065 ( 
.A1(n_909),
.A2(n_76),
.A3(n_77),
.B1(n_78),
.B2(n_80),
.C(n_81),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_921),
.B(n_78),
.Y(n_1066)
);

AOI33xp33_ASAP7_75t_L g1067 ( 
.A1(n_903),
.A2(n_971),
.A3(n_908),
.B1(n_968),
.B2(n_918),
.B3(n_915),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_930),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_864),
.B(n_82),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_980),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_909),
.B(n_83),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_L g1072 ( 
.A(n_856),
.B(n_83),
.C(n_84),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_920),
.B(n_85),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_864),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_864),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_942),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_942),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_971),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_836),
.Y(n_1079)
);

BUFx4f_ASAP7_75t_L g1080 ( 
.A(n_944),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_912),
.A2(n_914),
.B1(n_924),
.B2(n_923),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_912),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_SL g1083 ( 
.A(n_820),
.B(n_233),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_940),
.B(n_914),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_846),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_923),
.B(n_92),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_924),
.A2(n_93),
.B(n_94),
.C(n_95),
.Y(n_1087)
);

NOR2x1_ASAP7_75t_R g1088 ( 
.A(n_888),
.B(n_96),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_884),
.B(n_97),
.C(n_98),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_848),
.B(n_97),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_831),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_888),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_929),
.B(n_98),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_929),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_931),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_931),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_831),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_900),
.B(n_100),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_844),
.B(n_101),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_939),
.A2(n_853),
.B(n_850),
.C(n_845),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_939),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_902),
.B(n_101),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_932),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_935),
.B(n_936),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_916),
.B(n_103),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_942),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_857),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_933),
.B(n_106),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_932),
.B(n_108),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_861),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_1110)
);

CKINVDCx10_ASAP7_75t_R g1111 ( 
.A(n_844),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_932),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_820),
.B(n_238),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_949),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_938),
.B(n_113),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_926),
.B(n_114),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_928),
.A2(n_115),
.B(n_116),
.C(n_117),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_932),
.B(n_115),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_944),
.Y(n_1119)
);

AOI33xp33_ASAP7_75t_L g1120 ( 
.A1(n_948),
.A2(n_117),
.A3(n_118),
.B1(n_119),
.B2(n_120),
.B3(n_121),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_820),
.B(n_118),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_975),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_975),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_899),
.B(n_120),
.Y(n_1124)
);

CKINVDCx8_ASAP7_75t_R g1125 ( 
.A(n_963),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_953),
.B(n_121),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_944),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_978),
.B(n_122),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_L g1129 ( 
.A(n_963),
.B(n_970),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_904),
.B(n_122),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_917),
.B(n_125),
.Y(n_1131)
);

NOR2xp67_ASAP7_75t_L g1132 ( 
.A(n_977),
.B(n_126),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_943),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_961),
.B(n_137),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_960),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_957),
.B(n_138),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_964),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_962),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_973),
.B(n_139),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_954),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_951),
.B(n_144),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_969),
.B(n_144),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_946),
.B(n_145),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_950),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_947),
.B(n_151),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_952),
.B(n_152),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_945),
.B(n_152),
.Y(n_1147)
);

INVx11_ASAP7_75t_L g1148 ( 
.A(n_955),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_958),
.B(n_153),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_976),
.B(n_154),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_965),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_966),
.A2(n_272),
.B(n_307),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_972),
.A2(n_974),
.B(n_979),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1004),
.B(n_157),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_989),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1022),
.B(n_159),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1076),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1099),
.A2(n_159),
.B(n_161),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_983),
.B(n_1101),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_989),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1094),
.B(n_161),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1010),
.A2(n_162),
.B(n_163),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1076),
.B(n_162),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1002),
.B(n_164),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1070),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1053),
.A2(n_246),
.A3(n_247),
.B(n_248),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1095),
.B(n_249),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1135),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_SL g1169 ( 
.A1(n_1081),
.A2(n_1152),
.B(n_1040),
.Y(n_1169)
);

AND3x2_ASAP7_75t_L g1170 ( 
.A(n_1062),
.B(n_253),
.C(n_254),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1050),
.B(n_269),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_SL g1172 ( 
.A(n_1130),
.B(n_982),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_1017),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1084),
.A2(n_296),
.B(n_300),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1081),
.B(n_302),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_995),
.A2(n_997),
.B(n_996),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1044),
.B(n_1055),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1026),
.B(n_986),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_1076),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1024),
.B(n_1056),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1058),
.B(n_1122),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1123),
.A2(n_1023),
.B(n_1034),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1012),
.A2(n_1006),
.B(n_1118),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_SL g1184 ( 
.A(n_1125),
.B(n_994),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1038),
.A2(n_1098),
.B(n_1052),
.C(n_1018),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1042),
.Y(n_1186)
);

OA22x2_ASAP7_75t_L g1187 ( 
.A1(n_1063),
.A2(n_1070),
.B1(n_1025),
.B2(n_1130),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1008),
.A2(n_1011),
.B(n_1100),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1119),
.B(n_1092),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1063),
.A2(n_1032),
.A3(n_1021),
.B(n_1013),
.Y(n_1190)
);

AOI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_999),
.A2(n_1102),
.B(n_1029),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1137),
.B(n_993),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1039),
.B(n_987),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1005),
.A2(n_1015),
.B1(n_1108),
.B2(n_1036),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1091),
.B(n_1127),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_SL g1196 ( 
.A(n_1042),
.B(n_1089),
.C(n_1085),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1086),
.A2(n_1093),
.B(n_1061),
.C(n_1087),
.Y(n_1197)
);

NOR2x1_ASAP7_75t_L g1198 ( 
.A(n_1072),
.B(n_1130),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1035),
.A2(n_1047),
.B(n_1028),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_998),
.B(n_1019),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1054),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1068),
.A2(n_1117),
.A3(n_1082),
.B(n_1110),
.Y(n_1202)
);

CKINVDCx16_ASAP7_75t_R g1203 ( 
.A(n_1106),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1027),
.B(n_981),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_992),
.B(n_1003),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1054),
.A2(n_1041),
.B1(n_988),
.B2(n_1141),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1059),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1080),
.B(n_1000),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1078),
.B(n_1071),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1060),
.A2(n_1105),
.B(n_1048),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1073),
.B(n_1020),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1097),
.B(n_1014),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1064),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1136),
.A2(n_1126),
.B(n_1147),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1048),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1109),
.A2(n_1142),
.B(n_1116),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1121),
.A2(n_1128),
.B(n_1043),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1079),
.A2(n_1083),
.B(n_1113),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1139),
.A2(n_1115),
.B(n_1045),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1016),
.B(n_1104),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1149),
.A2(n_1124),
.B(n_1049),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_985),
.B(n_1031),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1088),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1083),
.A2(n_1113),
.B(n_1129),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1051),
.B(n_1066),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1134),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1112),
.B(n_1134),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1131),
.B(n_1114),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1000),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1143),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1074),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_1120),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1138),
.B(n_1103),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1107),
.A2(n_1151),
.A3(n_1144),
.B(n_1140),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1146),
.B(n_1090),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1145),
.B(n_1069),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1133),
.A2(n_1132),
.B1(n_1148),
.B2(n_1075),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1111),
.Y(n_1238)
);

AOI21xp33_ASAP7_75t_L g1239 ( 
.A1(n_1065),
.A2(n_1150),
.B(n_1009),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1065),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1046),
.A2(n_984),
.A3(n_1053),
.B(n_1081),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1030),
.A2(n_984),
.B(n_1001),
.Y(n_1242)
);

CKINVDCx8_ASAP7_75t_R g1243 ( 
.A(n_1030),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_984),
.A2(n_731),
.B(n_859),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1101),
.B(n_765),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1101),
.B(n_765),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1248)
);

NOR2x1_ASAP7_75t_R g1249 ( 
.A(n_994),
.B(n_901),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1101),
.B(n_765),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_984),
.A2(n_1007),
.B(n_990),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_984),
.A2(n_1053),
.A3(n_1081),
.B(n_1100),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1254)
);

NOR4xp25_ASAP7_75t_L g1255 ( 
.A(n_1065),
.B(n_1063),
.C(n_860),
.D(n_1082),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1042),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_982),
.B(n_986),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1101),
.B(n_765),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1101),
.B(n_765),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_984),
.A2(n_1053),
.A3(n_1081),
.B(n_1100),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1101),
.B(n_765),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1081),
.A2(n_1094),
.B1(n_1096),
.B2(n_1095),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1004),
.B(n_828),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1101),
.B(n_765),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1081),
.A2(n_1094),
.B1(n_1096),
.B2(n_1095),
.Y(n_1267)
);

AO21x1_ASAP7_75t_L g1268 ( 
.A1(n_1053),
.A2(n_1063),
.B(n_1083),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1004),
.B(n_828),
.Y(n_1269)
);

NOR2x1_ASAP7_75t_L g1270 ( 
.A(n_994),
.B(n_1070),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1022),
.Y(n_1271)
);

AO21x2_ASAP7_75t_L g1272 ( 
.A1(n_1023),
.A2(n_984),
.B(n_1100),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_984),
.A2(n_731),
.B(n_859),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1081),
.A2(n_1094),
.B1(n_1096),
.B2(n_1095),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1081),
.A2(n_1094),
.B1(n_1096),
.B2(n_1095),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1004),
.B(n_828),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1099),
.A2(n_707),
.B(n_766),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1004),
.B(n_828),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1037),
.A2(n_1033),
.B(n_991),
.C(n_1067),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_982),
.B(n_986),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1037),
.A2(n_1033),
.B(n_991),
.C(n_1067),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_984),
.A2(n_1053),
.A3(n_1081),
.B(n_1100),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1023),
.A2(n_984),
.B(n_1100),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1097),
.B(n_707),
.Y(n_1284)
);

CKINVDCx8_ASAP7_75t_R g1285 ( 
.A(n_1111),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1081),
.A2(n_1094),
.B1(n_1096),
.B2(n_1095),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_L g1287 ( 
.A(n_1097),
.B(n_707),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1004),
.A2(n_891),
.B1(n_745),
.B2(n_821),
.C(n_860),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1053),
.A2(n_1063),
.B(n_1083),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1070),
.A2(n_707),
.B1(n_766),
.B2(n_818),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1292)
);

NOR2x1_ASAP7_75t_SL g1293 ( 
.A(n_1053),
.B(n_1130),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_989),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1101),
.B(n_765),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_983),
.Y(n_1296)
);

NOR2x1_ASAP7_75t_SL g1297 ( 
.A(n_1053),
.B(n_1130),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_984),
.A2(n_731),
.B(n_859),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1004),
.B(n_828),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1101),
.B(n_765),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_994),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1101),
.B(n_765),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_982),
.B(n_986),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1004),
.B(n_828),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1004),
.B(n_828),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1004),
.B(n_828),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1004),
.B(n_828),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1097),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1153),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_989),
.B(n_1076),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_984),
.A2(n_1001),
.B(n_1010),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1081),
.A2(n_1094),
.B1(n_1096),
.B2(n_1095),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1101),
.B(n_765),
.Y(n_1315)
);

NOR2xp67_ASAP7_75t_L g1316 ( 
.A(n_1097),
.B(n_707),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1317)
);

NAND2x1_ASAP7_75t_L g1318 ( 
.A(n_1076),
.B(n_1077),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1076),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_L g1320 ( 
.A(n_1074),
.B(n_818),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_SL g1321 ( 
.A(n_1053),
.B(n_1130),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1004),
.B(n_828),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1099),
.A2(n_707),
.B(n_766),
.Y(n_1324)
);

AO21x1_ASAP7_75t_L g1325 ( 
.A1(n_1053),
.A2(n_1063),
.B(n_1083),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_994),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1256),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1224),
.A2(n_1169),
.B(n_1262),
.Y(n_1328)
);

OAI222xp33_ASAP7_75t_L g1329 ( 
.A1(n_1187),
.A2(n_1215),
.B1(n_1262),
.B2(n_1267),
.C1(n_1314),
.C2(n_1274),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1187),
.A2(n_1172),
.B1(n_1274),
.B2(n_1267),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1229),
.A2(n_1288),
.B1(n_1233),
.B2(n_1278),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1197),
.A2(n_1281),
.B(n_1279),
.Y(n_1332)
);

CKINVDCx12_ASAP7_75t_R g1333 ( 
.A(n_1249),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1265),
.B(n_1276),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1243),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1275),
.A2(n_1286),
.B1(n_1314),
.B2(n_1297),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1269),
.A2(n_1309),
.B1(n_1305),
.B2(n_1275),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1242),
.A2(n_1176),
.B(n_1244),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1307),
.B(n_1322),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1203),
.Y(n_1341)
);

AO21x1_ASAP7_75t_L g1342 ( 
.A1(n_1237),
.A2(n_1206),
.B(n_1286),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1292),
.B(n_1304),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1186),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1158),
.A2(n_1308),
.B1(n_1317),
.B2(n_1304),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1168),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_1248),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1157),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1218),
.A2(n_1175),
.B(n_1188),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1263),
.A2(n_1291),
.B(n_1264),
.Y(n_1350)
);

AO221x2_ASAP7_75t_L g1351 ( 
.A1(n_1290),
.A2(n_1324),
.B1(n_1277),
.B2(n_1162),
.C(n_1206),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1264),
.A2(n_1313),
.B(n_1291),
.Y(n_1352)
);

AOI21xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1238),
.A2(n_1310),
.B(n_1208),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1323),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1180),
.B(n_1246),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1285),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1168),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1268),
.B(n_1289),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1326),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1185),
.A2(n_1183),
.B(n_1245),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1160),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1293),
.A2(n_1321),
.B1(n_1210),
.B2(n_1226),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1296),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1181),
.B(n_1201),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1223),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1159),
.B(n_1227),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1192),
.A2(n_1227),
.B1(n_1193),
.B2(n_1177),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1247),
.B(n_1250),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1155),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1179),
.B(n_1319),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1177),
.A2(n_1228),
.B1(n_1154),
.B2(n_1161),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1311),
.A2(n_1182),
.B(n_1199),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1325),
.A2(n_1182),
.B(n_1199),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1258),
.B(n_1259),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1261),
.B(n_1266),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_SL g1376 ( 
.A1(n_1174),
.A2(n_1237),
.B(n_1211),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1251),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1295),
.B(n_1300),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1240),
.A2(n_1228),
.B1(n_1163),
.B2(n_1225),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1302),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1294),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1183),
.A2(n_1298),
.B(n_1273),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1294),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1225),
.A2(n_1221),
.B(n_1214),
.C(n_1204),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1315),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1200),
.Y(n_1386)
);

OAI222xp33_ASAP7_75t_L g1387 ( 
.A1(n_1198),
.A2(n_1163),
.B1(n_1194),
.B2(n_1232),
.C1(n_1211),
.C2(n_1213),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1271),
.B(n_1178),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1230),
.A2(n_1207),
.B1(n_1220),
.B2(n_1204),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1196),
.A2(n_1219),
.B1(n_1221),
.B2(n_1209),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1219),
.A2(n_1209),
.B1(n_1220),
.B2(n_1214),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1270),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1164),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1156),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1301),
.B(n_1165),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1173),
.B(n_1212),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1255),
.A2(n_1222),
.B1(n_1217),
.B2(n_1320),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1257),
.B(n_1280),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1167),
.A2(n_1205),
.B1(n_1236),
.B2(n_1235),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1272),
.A2(n_1283),
.B(n_1216),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_L g1401 ( 
.A(n_1284),
.B(n_1316),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1184),
.B(n_1318),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1303),
.Y(n_1403)
);

BUFx12f_ASAP7_75t_L g1404 ( 
.A(n_1231),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1195),
.B(n_1287),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1189),
.A2(n_1171),
.B1(n_1235),
.B2(n_1205),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1239),
.A2(n_1191),
.B(n_1312),
.Y(n_1407)
);

NOR2xp67_ASAP7_75t_SL g1408 ( 
.A(n_1170),
.B(n_1166),
.Y(n_1408)
);

AOI222xp33_ASAP7_75t_L g1409 ( 
.A1(n_1202),
.A2(n_1234),
.B1(n_1253),
.B2(n_1260),
.C1(n_1282),
.C2(n_1166),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1190),
.B(n_1241),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1190),
.B(n_1252),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1256),
.Y(n_1412)
);

AO32x2_ASAP7_75t_L g1413 ( 
.A1(n_1237),
.A2(n_1063),
.A3(n_1267),
.B1(n_1274),
.B2(n_1262),
.Y(n_1413)
);

INVxp33_ASAP7_75t_L g1414 ( 
.A(n_1159),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1265),
.B(n_1276),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1256),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1262),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1215),
.A2(n_1262),
.B1(n_1274),
.B2(n_1267),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1187),
.A2(n_1215),
.B1(n_1000),
.B2(n_1229),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1252),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1265),
.B(n_1276),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1197),
.A2(n_1026),
.B(n_1101),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1187),
.A2(n_1215),
.B1(n_1000),
.B2(n_1229),
.Y(n_1423)
);

AOI21xp33_ASAP7_75t_L g1424 ( 
.A1(n_1210),
.A2(n_1050),
.B(n_1237),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1340),
.B(n_1337),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1351),
.A2(n_1345),
.B1(n_1338),
.B2(n_1418),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1404),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1340),
.B(n_1421),
.Y(n_1428)
);

BUFx8_ASAP7_75t_L g1429 ( 
.A(n_1343),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1343),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1354),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_L g1432 ( 
.A(n_1354),
.Y(n_1432)
);

CKINVDCx6p67_ASAP7_75t_R g1433 ( 
.A(n_1333),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1420),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1422),
.A2(n_1371),
.B(n_1338),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1341),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1363),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1349),
.A2(n_1332),
.B(n_1382),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1364),
.B(n_1351),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1370),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_SL g1441 ( 
.A1(n_1345),
.A2(n_1418),
.B(n_1329),
.C(n_1379),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1351),
.B(n_1386),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_R g1443 ( 
.A(n_1412),
.B(n_1416),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1367),
.B(n_1417),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1391),
.B(n_1331),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1411),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1391),
.B(n_1331),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1348),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1399),
.A2(n_1384),
.B(n_1389),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1415),
.B(n_1334),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1390),
.B(n_1330),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1417),
.B(n_1369),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1390),
.B(n_1330),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1406),
.A2(n_1376),
.B1(n_1327),
.B2(n_1344),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1395),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1342),
.B(n_1328),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1374),
.B(n_1380),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1381),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1413),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1385),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1383),
.B(n_1368),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1375),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1395),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1384),
.A2(n_1407),
.B(n_1360),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_SL g1466 ( 
.A(n_1359),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1355),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1377),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1341),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1327),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1347),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1388),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1378),
.B(n_1355),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1395),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1335),
.Y(n_1475)
);

CKINVDCx6p67_ASAP7_75t_R g1476 ( 
.A(n_1359),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1405),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1414),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1452),
.B(n_1350),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_1410),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1456),
.B(n_1352),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1434),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1442),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1456),
.B(n_1409),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1445),
.B(n_1336),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1434),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1429),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1456),
.B(n_1442),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1445),
.B(n_1336),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1429),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1429),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1472),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1373),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1440),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1465),
.B(n_1478),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1432),
.B(n_1329),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1426),
.A2(n_1424),
.B1(n_1397),
.B2(n_1394),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1431),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1461),
.B(n_1358),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1471),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1440),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1440),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1447),
.B(n_1397),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1461),
.B(n_1400),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_L g1507 ( 
.A(n_1448),
.B(n_1387),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1482),
.B(n_1494),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1506),
.B(n_1459),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1500),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1502),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1493),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1482),
.B(n_1438),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1482),
.B(n_1339),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1500),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1488),
.B(n_1470),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1505),
.B(n_1449),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1496),
.B(n_1432),
.Y(n_1518)
);

NOR2x1_ASAP7_75t_SL g1519 ( 
.A(n_1488),
.B(n_1455),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1487),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1505),
.B(n_1451),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1497),
.B(n_1451),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1496),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1501),
.B(n_1458),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1483),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1499),
.A2(n_1435),
.B1(n_1430),
.B2(n_1454),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1497),
.B(n_1372),
.Y(n_1527)
);

AND2x2_ASAP7_75t_SL g1528 ( 
.A(n_1481),
.B(n_1432),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1484),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1486),
.B(n_1453),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1510),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1512),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1523),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1511),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1510),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1515),
.Y(n_1539)
);

NOR2xp67_ASAP7_75t_L g1540 ( 
.A(n_1525),
.B(n_1488),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1517),
.B(n_1486),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1517),
.B(n_1490),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1523),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1520),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1508),
.B(n_1489),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1513),
.B(n_1527),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1546),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1536),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1534),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1548),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1537),
.B(n_1547),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1542),
.B(n_1522),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1538),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1540),
.B(n_1514),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1536),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1546),
.Y(n_1567)
);

NAND4xp25_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1526),
.C(n_1498),
.D(n_1490),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1534),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1533),
.B(n_1527),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1537),
.B(n_1491),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1538),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1533),
.B(n_1535),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1532),
.Y(n_1574)
);

INVx5_ASAP7_75t_L g1575 ( 
.A(n_1541),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1539),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1557),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1560),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1556),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1560),
.Y(n_1580)
);

AOI222xp33_ASAP7_75t_L g1581 ( 
.A1(n_1574),
.A2(n_1526),
.B1(n_1543),
.B2(n_1542),
.C1(n_1521),
.C2(n_1530),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1535),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1562),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1556),
.Y(n_1584)
);

OAI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1568),
.A2(n_1561),
.B(n_1559),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1555),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1555),
.A2(n_1544),
.B(n_1545),
.Y(n_1587)
);

AOI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1571),
.A2(n_1516),
.B(n_1528),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1559),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1563),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1571),
.A2(n_1528),
.B1(n_1492),
.B2(n_1491),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1566),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1571),
.A2(n_1507),
.B(n_1344),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1563),
.Y(n_1595)
);

OAI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1557),
.A2(n_1353),
.B(n_1492),
.C(n_1491),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1564),
.Y(n_1597)
);

AOI21xp33_ASAP7_75t_L g1598 ( 
.A1(n_1569),
.A2(n_1543),
.B(n_1392),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1557),
.A2(n_1507),
.B(n_1492),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1565),
.A2(n_1528),
.B1(n_1518),
.B2(n_1476),
.Y(n_1600)
);

AOI21xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1592),
.A2(n_1577),
.B(n_1600),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1578),
.B(n_1547),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1570),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1577),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1577),
.Y(n_1605)
);

OAI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1585),
.A2(n_1569),
.B1(n_1567),
.B2(n_1554),
.C(n_1521),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1586),
.B(n_1570),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1595),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1597),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1581),
.A2(n_1530),
.B1(n_1498),
.B2(n_1522),
.C(n_1436),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1583),
.Y(n_1611)
);

AND3x2_ASAP7_75t_L g1612 ( 
.A(n_1599),
.B(n_1437),
.C(n_1433),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1598),
.A2(n_1453),
.B1(n_1439),
.B2(n_1514),
.Y(n_1613)
);

AOI322xp5_ASAP7_75t_L g1614 ( 
.A1(n_1587),
.A2(n_1544),
.A3(n_1573),
.B1(n_1549),
.B2(n_1545),
.C1(n_1550),
.C2(n_1551),
.Y(n_1614)
);

OAI322xp33_ASAP7_75t_L g1615 ( 
.A1(n_1590),
.A2(n_1582),
.A3(n_1588),
.B1(n_1591),
.B2(n_1589),
.C1(n_1583),
.C2(n_1495),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1605),
.B(n_1596),
.C(n_1594),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1615),
.A2(n_1591),
.B1(n_1589),
.B2(n_1441),
.C(n_1584),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1601),
.A2(n_1519),
.B(n_1565),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1614),
.B(n_1573),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_SL g1620 ( 
.A(n_1604),
.B(n_1470),
.C(n_1356),
.Y(n_1620)
);

AOI211xp5_ASAP7_75t_L g1621 ( 
.A1(n_1610),
.A2(n_1441),
.B(n_1443),
.C(n_1401),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1605),
.A2(n_1518),
.B(n_1362),
.Y(n_1622)
);

OAI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1606),
.A2(n_1565),
.B(n_1469),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1613),
.A2(n_1519),
.B(n_1608),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1612),
.A2(n_1427),
.B(n_1518),
.Y(n_1625)
);

AOI221x1_ASAP7_75t_L g1626 ( 
.A1(n_1609),
.A2(n_1477),
.B1(n_1584),
.B2(n_1593),
.C(n_1579),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1613),
.B(n_1408),
.C(n_1579),
.Y(n_1627)
);

OAI31xp33_ASAP7_75t_L g1628 ( 
.A1(n_1602),
.A2(n_1523),
.A3(n_1518),
.B(n_1503),
.Y(n_1628)
);

OAI211xp5_ASAP7_75t_L g1629 ( 
.A1(n_1612),
.A2(n_1365),
.B(n_1469),
.C(n_1436),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1603),
.A2(n_1503),
.B(n_1504),
.C(n_1496),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1607),
.B(n_1551),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1611),
.A2(n_1467),
.B1(n_1439),
.B2(n_1514),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1617),
.A2(n_1593),
.B1(n_1572),
.B2(n_1576),
.C(n_1564),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1362),
.B(n_1387),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1619),
.B(n_1549),
.Y(n_1635)
);

NAND4xp75_ASAP7_75t_L g1636 ( 
.A(n_1624),
.B(n_1433),
.C(n_1476),
.D(n_1475),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_SL g1637 ( 
.A(n_1629),
.B(n_1495),
.C(n_1550),
.D(n_1466),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1623),
.B(n_1552),
.Y(n_1638)
);

NOR2xp67_ASAP7_75t_L g1639 ( 
.A(n_1618),
.B(n_1575),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1628),
.B(n_1427),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1626),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1620),
.A2(n_1428),
.B(n_1425),
.Y(n_1642)
);

NOR3x1_ASAP7_75t_L g1643 ( 
.A(n_1625),
.B(n_1475),
.C(n_1463),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1622),
.B(n_1632),
.Y(n_1644)
);

NOR3x1_ASAP7_75t_L g1645 ( 
.A(n_1636),
.B(n_1627),
.C(n_1621),
.Y(n_1645)
);

NOR4xp25_ASAP7_75t_L g1646 ( 
.A(n_1641),
.B(n_1633),
.C(n_1637),
.D(n_1640),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1644),
.A2(n_1632),
.B1(n_1630),
.B2(n_1631),
.C(n_1464),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1638),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1640),
.B(n_1365),
.C(n_1335),
.Y(n_1649)
);

NOR3xp33_ASAP7_75t_L g1650 ( 
.A(n_1634),
.B(n_1396),
.C(n_1357),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1635),
.B(n_1552),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1642),
.Y(n_1652)
);

NOR3xp33_ASAP7_75t_L g1653 ( 
.A(n_1639),
.B(n_1396),
.C(n_1346),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1361),
.C(n_1403),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1633),
.B(n_1427),
.C(n_1479),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1633),
.A2(n_1427),
.B(n_1450),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1652),
.B(n_1427),
.Y(n_1657)
);

NAND4xp75_ASAP7_75t_L g1658 ( 
.A(n_1645),
.B(n_1473),
.C(n_1455),
.D(n_1463),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1647),
.B(n_1503),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1572),
.Y(n_1660)
);

XNOR2xp5_ASAP7_75t_L g1661 ( 
.A(n_1650),
.B(n_1462),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1648),
.Y(n_1662)
);

XNOR2xp5_ASAP7_75t_L g1663 ( 
.A(n_1646),
.B(n_1457),
.Y(n_1663)
);

AND3x1_ASAP7_75t_L g1664 ( 
.A(n_1653),
.B(n_1474),
.C(n_1460),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1656),
.B(n_1504),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1657),
.Y(n_1666)
);

XNOR2xp5_ASAP7_75t_L g1667 ( 
.A(n_1663),
.B(n_1654),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1661),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1662),
.B(n_1655),
.Y(n_1669)
);

NAND4xp75_ASAP7_75t_L g1670 ( 
.A(n_1659),
.B(n_1651),
.C(n_1474),
.D(n_1393),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1660),
.B(n_1576),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1668),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_1670),
.B(n_1658),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_L g1674 ( 
.A(n_1669),
.B(n_1665),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1664),
.Y(n_1675)
);

AO22x2_ASAP7_75t_L g1676 ( 
.A1(n_1672),
.A2(n_1666),
.B1(n_1669),
.B2(n_1667),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1674),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1676),
.A2(n_1673),
.B1(n_1675),
.B2(n_1666),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1678),
.B(n_1677),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1679),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1680),
.B(n_1671),
.Y(n_1681)
);

NAND2x2_ASAP7_75t_L g1682 ( 
.A(n_1681),
.B(n_1504),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1398),
.B1(n_1402),
.B2(n_1366),
.Y(n_1683)
);


endmodule