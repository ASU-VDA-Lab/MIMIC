module fake_jpeg_3269_n_542 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g125 ( 
.A(n_47),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_56),
.Y(n_98)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_54),
.Y(n_116)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_63),
.Y(n_112)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_59),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_77),
.Y(n_119)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_9),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_69),
.B(n_32),
.C(n_31),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_16),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_18),
.Y(n_131)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_79),
.B1(n_46),
.B2(n_38),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_99),
.A2(n_44),
.B1(n_92),
.B2(n_89),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_104),
.B(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_110),
.B(n_117),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_41),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_62),
.A2(n_19),
.B(n_41),
.Y(n_123)
);

OR2x4_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_48),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_13),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_45),
.A2(n_17),
.B1(n_28),
.B2(n_39),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_133),
.A2(n_153),
.B1(n_49),
.B2(n_60),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_32),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_53),
.B(n_17),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_157),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_54),
.A2(n_39),
.B1(n_28),
.B2(n_40),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_152),
.A2(n_96),
.B1(n_72),
.B2(n_48),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_38),
.B1(n_44),
.B2(n_40),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_81),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_65),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_167),
.Y(n_229)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g169 ( 
.A(n_125),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_169),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_178),
.Y(n_215)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_198),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_202),
.B(n_203),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_208)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_59),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_187),
.Y(n_225)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_66),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_71),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_192),
.Y(n_238)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_147),
.B1(n_148),
.B2(n_108),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_197),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_61),
.B1(n_64),
.B2(n_74),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_108),
.B1(n_118),
.B2(n_105),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_97),
.A2(n_73),
.A3(n_84),
.B1(n_70),
.B2(n_86),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_136),
.A2(n_44),
.B1(n_85),
.B2(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_95),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_99),
.B(n_158),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_209),
.A2(n_224),
.B(n_188),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_210),
.A2(n_217),
.B1(n_232),
.B2(n_233),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_169),
.A2(n_155),
.B(n_114),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_193),
.A2(n_137),
.B1(n_122),
.B2(n_135),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_198),
.A2(n_137),
.B1(n_122),
.B2(n_135),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_184),
.B(n_207),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_184),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_163),
.B(n_161),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_225),
.Y(n_257)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_246),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_189),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_249),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_251),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_165),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_252),
.B(n_257),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_254),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_243),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_240),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_266),
.B(n_267),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_195),
.B1(n_204),
.B2(n_118),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_273),
.B1(n_105),
.B2(n_235),
.Y(n_298)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_216),
.B(n_173),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_271),
.Y(n_297)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_263),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_238),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_179),
.Y(n_302)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_225),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_219),
.A2(n_194),
.B(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_211),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_209),
.A2(n_173),
.B(n_160),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_272),
.B(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_142),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_186),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_217),
.A2(n_113),
.B1(n_181),
.B2(n_176),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_212),
.A2(n_155),
.B1(n_168),
.B2(n_164),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_145),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_226),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_218),
.A2(n_206),
.B(n_156),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_276),
.A2(n_238),
.B(n_215),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_250),
.A2(n_234),
.B1(n_208),
.B2(n_232),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_300),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_233),
.B1(n_218),
.B2(n_237),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_279),
.A2(n_261),
.B1(n_249),
.B2(n_247),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_223),
.B1(n_215),
.B2(n_230),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_294),
.B1(n_274),
.B2(n_250),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_308),
.B(n_276),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_255),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_251),
.A2(n_223),
.B1(n_230),
.B2(n_235),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_240),
.C(n_231),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_269),
.C(n_264),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

AO21x1_ASAP7_75t_SL g305 ( 
.A1(n_267),
.A2(n_120),
.B(n_127),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_256),
.B(n_222),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_267),
.A2(n_222),
.B(n_220),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_263),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_281),
.B(n_287),
.C(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_320),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_257),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_311),
.B(n_323),
.Y(n_375)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_253),
.Y(n_316)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_316),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_317),
.A2(n_342),
.B(n_241),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_292),
.C(n_288),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_249),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_252),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_254),
.Y(n_325)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_255),
.B(n_275),
.C(n_271),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_328),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_293),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_302),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_340),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_266),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_332),
.B(n_170),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_333),
.A2(n_222),
.B(n_106),
.Y(n_374)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_334),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_278),
.B(n_272),
.Y(n_335)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_245),
.Y(n_338)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_279),
.A2(n_283),
.B1(n_277),
.B2(n_305),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_339),
.A2(n_260),
.B1(n_262),
.B2(n_246),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_263),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_341),
.A2(n_297),
.B1(n_308),
.B2(n_288),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_241),
.B(n_226),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_221),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_345),
.B(n_364),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_348),
.B(n_314),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_351),
.A2(n_359),
.B1(n_372),
.B2(n_315),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_329),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_308),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_376),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_317),
.A2(n_301),
.B(n_299),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_357),
.A2(n_358),
.B(n_363),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_307),
.B(n_304),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_336),
.A2(n_295),
.B1(n_290),
.B2(n_280),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_295),
.C(n_290),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_324),
.C(n_340),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_314),
.A2(n_280),
.B1(n_282),
.B2(n_303),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_361),
.A2(n_368),
.B1(n_313),
.B2(n_319),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_333),
.A2(n_303),
.B(n_282),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_221),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_220),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_369),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_SL g406 ( 
.A(n_370),
.B(n_315),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_260),
.B1(n_262),
.B2(n_244),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_374),
.A2(n_315),
.B(n_326),
.C(n_340),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_93),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_399),
.Y(n_412)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_379),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_328),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_380),
.B(n_382),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_392),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_343),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_384),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_310),
.C(n_324),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_389),
.C(n_408),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_365),
.A2(n_339),
.B1(n_331),
.B2(n_313),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_387),
.A2(n_400),
.B1(n_401),
.B2(n_372),
.Y(n_411)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_342),
.C(n_322),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_321),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_391),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_320),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_393),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_321),
.Y(n_394)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_394),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_350),
.B(n_319),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_356),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_346),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_402),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_362),
.B(n_334),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_398),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_347),
.A2(n_313),
.B1(n_329),
.B2(n_322),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_338),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_374),
.B1(n_354),
.B2(n_312),
.Y(n_428)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_315),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_361),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_406),
.A2(n_106),
.B(n_150),
.Y(n_436)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_213),
.C(n_199),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_414),
.B1(n_422),
.B2(n_383),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_387),
.A2(n_366),
.B1(n_371),
.B2(n_356),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_392),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_399),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_183),
.Y(n_454)
);

AOI21xp33_ASAP7_75t_L g419 ( 
.A1(n_395),
.A2(n_366),
.B(n_357),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_419),
.A2(n_109),
.B(n_138),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_373),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_436),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_384),
.A2(n_363),
.B1(n_373),
.B2(n_358),
.Y(n_422)
);

FAx1_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_374),
.CI(n_359),
.CON(n_423),
.SN(n_423)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_423),
.A2(n_146),
.B(n_101),
.C(n_179),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_424),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_428),
.A2(n_431),
.B1(n_407),
.B2(n_378),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_389),
.A2(n_213),
.B1(n_159),
.B2(n_191),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_377),
.C(n_381),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_434),
.C(n_408),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_213),
.C(n_128),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_446),
.Y(n_469)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_455),
.B1(n_461),
.B2(n_436),
.Y(n_467)
);

BUFx12_ASAP7_75t_L g440 ( 
.A(n_423),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_442),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_441),
.B(n_431),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_383),
.C(n_385),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_413),
.A2(n_205),
.B(n_162),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_443),
.B(n_445),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_138),
.C(n_128),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_177),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_447),
.B(n_429),
.Y(n_475)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_450),
.Y(n_472)
);

XOR2x2_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_447),
.Y(n_473)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_425),
.B(n_171),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_451),
.B(n_453),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_422),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_458),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_190),
.B1(n_146),
.B2(n_143),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_457),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_134),
.C(n_179),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_412),
.B(n_433),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_412),
.B(n_140),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_460),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_109),
.B1(n_127),
.B2(n_101),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_434),
.C(n_414),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_464),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_458),
.B(n_421),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_477),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_446),
.C(n_444),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_428),
.B1(n_423),
.B2(n_435),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_474),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_473),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_429),
.C(n_410),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_480),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_410),
.C(n_416),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_478),
.B(n_440),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_409),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_470),
.A2(n_452),
.B(n_445),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_482),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_460),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_487),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_409),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_440),
.C(n_101),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_489),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_476),
.B(n_468),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_493),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_466),
.A2(n_53),
.B(n_82),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_492),
.A2(n_473),
.B(n_475),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_84),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_11),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_497),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_472),
.A2(n_82),
.B1(n_11),
.B2(n_12),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_10),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_498),
.B(n_9),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_474),
.A2(n_73),
.B1(n_10),
.B2(n_11),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_493),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_462),
.C(n_480),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_505),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_502),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_490),
.A2(n_477),
.B(n_10),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_507),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_9),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_6),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_490),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_486),
.A2(n_488),
.B(n_485),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_512),
.Y(n_517)
);

INVx11_ASAP7_75t_L g514 ( 
.A(n_486),
.Y(n_514)
);

AOI31xp67_ASAP7_75t_L g522 ( 
.A1(n_514),
.A2(n_6),
.A3(n_14),
.B(n_12),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_508),
.B(n_499),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_519),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_491),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_500),
.B(n_6),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_523),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_522),
.A2(n_509),
.B1(n_502),
.B2(n_511),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_14),
.Y(n_523)
);

AOI322xp5_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_24),
.A3(n_37),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g525 ( 
.A1(n_510),
.A2(n_24),
.A3(n_37),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_516),
.Y(n_526)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_526),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_529),
.B(n_524),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_506),
.C(n_512),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_531),
.B1(n_532),
.B2(n_525),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_506),
.B(n_37),
.Y(n_531)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_520),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_533),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_536),
.B(n_528),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_1),
.B(n_5),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_534),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_530),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_537),
.Y(n_542)
);


endmodule