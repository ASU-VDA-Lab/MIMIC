module real_jpeg_13115_n_12 (n_5, n_4, n_8, n_0, n_278, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_278;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_2),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_3),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_43),
.B1(n_46),
.B2(n_154),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_100),
.B1(n_101),
.B2(n_154),
.Y(n_253)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_6),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_6),
.A2(n_45),
.B1(n_148),
.B2(n_149),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_7),
.B(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_27),
.C(n_48),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_30),
.B1(n_43),
.B2(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_7),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_7),
.B(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_7),
.A2(n_30),
.B1(n_100),
.B2(n_101),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_57),
.B(n_101),
.C(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_7),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_7),
.A2(n_30),
.B1(n_148),
.B2(n_149),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_10),
.A2(n_37),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_37),
.B1(n_148),
.B2(n_149),
.Y(n_161)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_256),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_237),
.B(n_255),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_216),
.B(n_236),
.Y(n_14)
);

AOI321xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_177),
.A3(n_209),
.B1(n_214),
.B2(n_215),
.C(n_278),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_138),
.B(n_176),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_116),
.B(n_137),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_93),
.B(n_115),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_71),
.B(n_92),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_23),
.B(n_89),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_35),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_30),
.A2(n_46),
.B(n_58),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_30),
.B(n_101),
.C(n_134),
.Y(n_147)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_32),
.A2(n_89),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_35),
.A2(n_153),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_41),
.B(n_68),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_41),
.A2(n_174),
.B(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_42),
.B(n_51),
.Y(n_108)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_47),
.Y(n_175)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_51),
.Y(n_174)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_59),
.C(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_99),
.Y(n_98)
);

NAND2x1_ASAP7_75t_SL g185 ( 
.A(n_55),
.B(n_106),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_55),
.A2(n_103),
.B(n_106),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_55),
.A2(n_170),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_56),
.B(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_70),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_85),
.B(n_91),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_79),
.B(n_84),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_81),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_107),
.C(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_101),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_102),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_104),
.B(n_127),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_104),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_108),
.A2(n_175),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_108),
.B(n_120),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_110),
.A2(n_111),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_110),
.A2(n_111),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_111),
.B(n_233),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_111),
.A2(n_244),
.B(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_136),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_136),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_131),
.C(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_126),
.B(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_126),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_133),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_133),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_135),
.B1(n_148),
.B2(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_140),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_156),
.B2(n_157),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_144),
.C(n_156),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_155),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_167),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_169),
.C(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_164),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_162),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_163),
.A2(n_166),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_182),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_172),
.A2(n_173),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_204),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_204),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_189),
.C(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_187),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_184),
.CI(n_187),
.CON(n_206),
.SN(n_206)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_181),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_200),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_197),
.C(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_193),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_206),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_206),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_213),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_235),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_231),
.B2(n_232),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_232),
.C(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.C(n_229),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_233),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_239),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_242),
.C(n_250),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_249),
.B2(n_250),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_263),
.B1(n_264),
.B2(n_274),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_254),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_275),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);


endmodule