module fake_jpeg_2035_n_51 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_51);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_51;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_20),
.B(n_18),
.Y(n_27)
);

CKINVDCx12_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

OAI22x1_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AND2x6_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_9),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_21),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_31),
.C(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_26),
.B1(n_24),
.B2(n_2),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_1),
.B(n_3),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

OA21x2_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_1),
.B(n_4),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_37),
.B1(n_39),
.B2(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_47),
.C(n_7),
.Y(n_50)
);

NOR3x1_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_5),
.C(n_8),
.Y(n_51)
);


endmodule