module real_aes_7721_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_753;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_88), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g461 ( .A(n_0), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_1), .A2(n_105), .B1(n_114), .B2(n_768), .Y(n_104) );
INVx1_ASAP7_75t_L g511 ( .A(n_2), .Y(n_511) );
INVx1_ASAP7_75t_L g208 ( .A(n_3), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_4), .A2(n_81), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_4), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_5), .A2(n_38), .B1(n_164), .B2(n_527), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g188 ( .A1(n_6), .A2(n_145), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_7), .B(n_138), .Y(n_502) );
AND2x6_ASAP7_75t_L g150 ( .A(n_8), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_9), .A2(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_10), .B(n_39), .Y(n_108) );
INVx1_ASAP7_75t_L g195 ( .A(n_11), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_12), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g143 ( .A(n_13), .Y(n_143) );
INVx1_ASAP7_75t_L g506 ( .A(n_14), .Y(n_506) );
INVx1_ASAP7_75t_L g253 ( .A(n_15), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_16), .B(n_176), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_17), .B(n_139), .Y(n_483) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_18), .A2(n_138), .A3(n_173), .B1(n_489), .B2(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_19), .B(n_164), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_20), .B(n_159), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_21), .B(n_139), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_22), .A2(n_52), .B1(n_164), .B2(n_527), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_23), .B(n_145), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g533 ( .A1(n_24), .A2(n_77), .B1(n_164), .B2(n_176), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_25), .B(n_164), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_26), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_27), .A2(n_251), .B(n_252), .C(n_254), .Y(n_250) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_29), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_29), .B(n_197), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_30), .B(n_193), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_31), .A2(n_42), .B1(n_759), .B2(n_760), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_31), .Y(n_759) );
INVx1_ASAP7_75t_L g182 ( .A(n_32), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_33), .B(n_197), .Y(n_550) );
INVx2_ASAP7_75t_L g148 ( .A(n_34), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_35), .B(n_164), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_36), .B(n_197), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_37), .A2(n_150), .B(n_154), .C(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g180 ( .A(n_40), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_41), .B(n_193), .Y(n_263) );
CKINVDCx14_ASAP7_75t_R g760 ( .A(n_42), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_43), .B(n_164), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_44), .A2(n_467), .B1(n_753), .B2(n_754), .C1(n_763), .C2(n_765), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_45), .A2(n_758), .B1(n_761), .B2(n_762), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_45), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_46), .A2(n_89), .B1(n_226), .B2(n_527), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_47), .B(n_164), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_48), .B(n_164), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_49), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_50), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_51), .B(n_145), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_53), .A2(n_62), .B1(n_164), .B2(n_176), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_54), .A2(n_154), .B1(n_176), .B2(n_178), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_55), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_56), .B(n_164), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_57), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_58), .B(n_164), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_59), .A2(n_163), .B(n_192), .C(n_194), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_60), .Y(n_267) );
INVx1_ASAP7_75t_L g190 ( .A(n_61), .Y(n_190) );
INVx1_ASAP7_75t_L g151 ( .A(n_63), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_64), .B(n_164), .Y(n_512) );
INVx1_ASAP7_75t_L g142 ( .A(n_65), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
AO32x2_ASAP7_75t_L g530 ( .A1(n_67), .A2(n_138), .A3(n_233), .B1(n_489), .B2(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g569 ( .A(n_68), .Y(n_569) );
INVx1_ASAP7_75t_L g545 ( .A(n_69), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_70), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_70), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_SL g158 ( .A1(n_71), .A2(n_159), .B(n_160), .C(n_163), .Y(n_158) );
INVxp67_ASAP7_75t_L g161 ( .A(n_72), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_73), .B(n_176), .Y(n_546) );
INVx1_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_75), .Y(n_186) );
INVx1_ASAP7_75t_L g260 ( .A(n_76), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_78), .B(n_463), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_79), .A2(n_150), .B(n_154), .C(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_80), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_81), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_82), .B(n_176), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_83), .B(n_209), .Y(n_222) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_85), .B(n_159), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_86), .B(n_176), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_87), .A2(n_150), .B(n_154), .C(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g458 ( .A(n_88), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g470 ( .A(n_88), .B(n_460), .Y(n_470) );
INVx2_ASAP7_75t_L g474 ( .A(n_88), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_90), .A2(n_103), .B1(n_176), .B2(n_177), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_91), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_92), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_93), .A2(n_150), .B(n_154), .C(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_94), .Y(n_243) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_96), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_97), .B(n_209), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_98), .B(n_176), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_99), .B(n_138), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_101), .A2(n_145), .B(n_152), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_102), .A2(n_124), .B1(n_125), .B2(n_128), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_102), .Y(n_128) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g768 ( .A(n_107), .Y(n_768) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g460 ( .A(n_108), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_465), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_115), .B(n_462), .C(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_455), .B(n_462), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_129), .B2(n_130), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22x1_ASAP7_75t_SL g763 ( .A1(n_129), .A2(n_473), .B1(n_476), .B2(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_130), .A2(n_468), .B1(n_471), .B2(n_475), .Y(n_467) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_392), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_322), .C(n_353), .D(n_372), .Y(n_131) );
NAND4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_280), .C(n_295), .D(n_313), .Y(n_132) );
AOI222xp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_215), .B1(n_256), .B2(n_268), .C1(n_273), .C2(n_275), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_198), .Y(n_134) );
INVx1_ASAP7_75t_L g336 ( .A(n_135), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
AND2x2_ASAP7_75t_L g199 ( .A(n_136), .B(n_187), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_136), .B(n_202), .Y(n_365) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g272 ( .A(n_137), .B(n_171), .Y(n_272) );
AND2x2_ASAP7_75t_L g281 ( .A(n_137), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g307 ( .A(n_137), .Y(n_307) );
AND2x2_ASAP7_75t_L g328 ( .A(n_137), .B(n_171), .Y(n_328) );
BUFx2_ASAP7_75t_L g351 ( .A(n_137), .Y(n_351) );
AND2x2_ASAP7_75t_L g375 ( .A(n_137), .B(n_172), .Y(n_375) );
AND2x2_ASAP7_75t_L g439 ( .A(n_137), .B(n_187), .Y(n_439) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_166), .Y(n_137) );
INVx4_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_138), .A2(n_494), .B(n_502), .Y(n_493) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_140), .B(n_141), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g247 ( .A(n_145), .Y(n_247) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_146), .B(n_150), .Y(n_184) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g501 ( .A(n_147), .Y(n_501) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
INVx4_ASAP7_75t_SL g165 ( .A(n_150), .Y(n_165) );
BUFx3_ASAP7_75t_L g489 ( .A(n_150), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_150), .A2(n_495), .B(n_498), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_150), .A2(n_505), .B(n_509), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_150), .A2(n_520), .B(n_524), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_150), .A2(n_544), .B(n_547), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_158), .C(n_165), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_153), .A2(n_165), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_153), .A2(n_165), .B(n_249), .C(n_250), .Y(n_248) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
BUFx3_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
INVx1_ASAP7_75t_L g527 ( .A(n_155), .Y(n_527) );
INVx1_ASAP7_75t_L g523 ( .A(n_159), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_162), .B(n_195), .Y(n_194) );
INVx5_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g531 ( .A1(n_162), .A2(n_193), .B1(n_532), .B2(n_533), .Y(n_531) );
O2A1O1Ixp5_ASAP7_75t_SL g544 ( .A1(n_163), .A2(n_209), .B(n_545), .C(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_164), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_165), .A2(n_175), .B1(n_183), .B2(n_184), .Y(n_174) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_167), .A2(n_188), .B(n_196), .Y(n_187) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g228 ( .A(n_168), .B(n_229), .Y(n_228) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_168), .B(n_485), .C(n_489), .Y(n_484) );
AO21x1_ASAP7_75t_L g577 ( .A1(n_168), .A2(n_485), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g340 ( .A(n_169), .B(n_271), .Y(n_340) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_170), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_187), .Y(n_170) );
OR2x2_ASAP7_75t_L g300 ( .A(n_171), .B(n_203), .Y(n_300) );
AND2x2_ASAP7_75t_L g312 ( .A(n_171), .B(n_271), .Y(n_312) );
BUFx2_ASAP7_75t_L g444 ( .A(n_171), .Y(n_444) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OR2x2_ASAP7_75t_L g201 ( .A(n_172), .B(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g294 ( .A(n_172), .B(n_203), .Y(n_294) );
AND2x2_ASAP7_75t_L g347 ( .A(n_172), .B(n_187), .Y(n_347) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_172), .Y(n_383) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_185), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_173), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_204), .B(n_212), .Y(n_203) );
INVx2_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
INVx2_ASAP7_75t_L g211 ( .A(n_176), .Y(n_211) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_178) );
INVx2_ASAP7_75t_L g181 ( .A(n_179), .Y(n_181) );
INVx4_ASAP7_75t_L g251 ( .A(n_179), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_184), .A2(n_205), .B(n_206), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_184), .A2(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g270 ( .A(n_187), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g282 ( .A(n_187), .Y(n_282) );
INVx2_ASAP7_75t_L g293 ( .A(n_187), .Y(n_293) );
BUFx2_ASAP7_75t_L g317 ( .A(n_187), .Y(n_317) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_187), .B(n_375), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_192), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp5_ASAP7_75t_L g568 ( .A1(n_192), .A2(n_510), .B(n_569), .C(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx4_ASAP7_75t_L g239 ( .A(n_193), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_193), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_193), .A2(n_487), .B1(n_537), .B2(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g214 ( .A(n_197), .Y(n_214) );
INVx2_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_197), .A2(n_246), .B(n_255), .Y(n_245) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_197), .A2(n_519), .B(n_528), .Y(n_518) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_197), .A2(n_543), .B(n_550), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AOI332xp33_ASAP7_75t_L g295 ( .A1(n_199), .A2(n_296), .A3(n_300), .B1(n_301), .B2(n_305), .B3(n_308), .C1(n_309), .C2(n_311), .Y(n_295) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_199), .B(n_271), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_199), .B(n_285), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_SL g313 ( .A1(n_200), .A2(n_314), .B(n_317), .C(n_318), .Y(n_313) );
AND2x2_ASAP7_75t_L g452 ( .A(n_200), .B(n_293), .Y(n_452) );
INVx3_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g349 ( .A(n_201), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g354 ( .A(n_201), .B(n_351), .Y(n_354) );
INVx1_ASAP7_75t_L g285 ( .A(n_202), .Y(n_285) );
AND2x2_ASAP7_75t_L g388 ( .A(n_202), .B(n_347), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_202), .B(n_328), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_202), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_202), .B(n_306), .Y(n_414) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g271 ( .A(n_203), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .C(n_211), .Y(n_207) );
INVx2_ASAP7_75t_L g487 ( .A(n_209), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_209), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_209), .A2(n_566), .B(n_567), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_211), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_214), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_214), .B(n_267), .Y(n_266) );
OAI31xp33_ASAP7_75t_L g453 ( .A1(n_215), .A2(n_374), .A3(n_381), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_230), .Y(n_215) );
AND2x2_ASAP7_75t_L g256 ( .A(n_216), .B(n_257), .Y(n_256) );
NAND2x1_ASAP7_75t_SL g276 ( .A(n_216), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_216), .Y(n_363) );
AND2x2_ASAP7_75t_L g368 ( .A(n_216), .B(n_279), .Y(n_368) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_217), .A2(n_281), .B(n_283), .C(n_286), .Y(n_280) );
OR2x2_ASAP7_75t_L g297 ( .A(n_217), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g310 ( .A(n_217), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_217), .B(n_258), .Y(n_316) );
INVx2_ASAP7_75t_L g334 ( .A(n_217), .Y(n_334) );
AND2x2_ASAP7_75t_L g345 ( .A(n_217), .B(n_299), .Y(n_345) );
AND2x2_ASAP7_75t_L g377 ( .A(n_217), .B(n_335), .Y(n_377) );
AND2x2_ASAP7_75t_L g381 ( .A(n_217), .B(n_304), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_217), .B(n_230), .Y(n_386) );
AND2x2_ASAP7_75t_L g420 ( .A(n_217), .B(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_217), .B(n_323), .Y(n_454) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_228), .Y(n_217) );
AOI21xp5_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_220), .B(n_227), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_224), .A2(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g254 ( .A(n_226), .Y(n_254) );
INVx1_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_227), .A2(n_504), .B(n_513), .Y(n_503) );
OA21x2_ASAP7_75t_L g563 ( .A1(n_227), .A2(n_564), .B(n_571), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_230), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g362 ( .A(n_230), .Y(n_362) );
AND2x2_ASAP7_75t_L g424 ( .A(n_230), .B(n_345), .Y(n_424) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_244), .Y(n_230) );
OR2x2_ASAP7_75t_L g278 ( .A(n_231), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g288 ( .A(n_231), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_231), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g396 ( .A(n_231), .Y(n_396) );
AND2x2_ASAP7_75t_L g413 ( .A(n_231), .B(n_258), .Y(n_413) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g304 ( .A(n_232), .B(n_244), .Y(n_304) );
AND2x2_ASAP7_75t_L g333 ( .A(n_232), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g344 ( .A(n_232), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_232), .B(n_299), .Y(n_435) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_242), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g257 ( .A(n_245), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g279 ( .A(n_245), .Y(n_279) );
AND2x2_ASAP7_75t_L g335 ( .A(n_245), .B(n_299), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_251), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g508 ( .A(n_251), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_251), .A2(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g437 ( .A(n_256), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_257), .Y(n_441) );
INVx2_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_265), .B(n_266), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_270), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_270), .B(n_375), .Y(n_433) );
OR2x2_ASAP7_75t_L g274 ( .A(n_271), .B(n_272), .Y(n_274) );
INVx1_ASAP7_75t_SL g326 ( .A(n_271), .Y(n_326) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_277), .A2(n_330), .B1(n_332), .B2(n_336), .C(n_337), .Y(n_329) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g357 ( .A(n_278), .B(n_321), .Y(n_357) );
INVx2_ASAP7_75t_L g289 ( .A(n_279), .Y(n_289) );
INVx1_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_279), .B(n_299), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_279), .B(n_302), .Y(n_409) );
INVx1_ASAP7_75t_L g417 ( .A(n_279), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_281), .B(n_285), .Y(n_331) );
AND2x4_ASAP7_75t_L g306 ( .A(n_282), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g419 ( .A(n_285), .B(n_375), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_288), .B(n_320), .Y(n_319) );
INVxp67_ASAP7_75t_L g427 ( .A(n_289), .Y(n_427) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_293), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g399 ( .A(n_293), .B(n_375), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_293), .B(n_312), .Y(n_405) );
AOI322xp5_ASAP7_75t_L g359 ( .A1(n_294), .A2(n_328), .A3(n_335), .B1(n_360), .B2(n_363), .C1(n_364), .C2(n_366), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_294), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g425 ( .A(n_297), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g371 ( .A(n_298), .Y(n_371) );
INVx2_ASAP7_75t_L g302 ( .A(n_299), .Y(n_302) );
INVx1_ASAP7_75t_L g361 ( .A(n_299), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_300), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g397 ( .A(n_302), .B(n_310), .Y(n_397) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_304), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g352 ( .A(n_304), .B(n_345), .Y(n_352) );
AND2x2_ASAP7_75t_L g356 ( .A(n_304), .B(n_316), .Y(n_356) );
OAI21xp33_ASAP7_75t_SL g366 ( .A1(n_305), .A2(n_367), .B(n_369), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_305), .A2(n_437), .B1(n_438), .B2(n_440), .Y(n_436) );
INVx3_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_306), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_306), .B(n_326), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_308), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g448 ( .A(n_315), .Y(n_448) );
INVx4_ASAP7_75t_L g321 ( .A(n_316), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_316), .B(n_343), .Y(n_391) );
INVx1_ASAP7_75t_SL g403 ( .A(n_317), .Y(n_403) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_321), .B(n_417), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_324), .B(n_329), .C(n_346), .Y(n_322) );
OAI221xp5_ASAP7_75t_SL g442 ( .A1(n_324), .A2(n_362), .B1(n_441), .B2(n_443), .C(n_445), .Y(n_442) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_326), .B(n_439), .Y(n_438) );
OAI31xp33_ASAP7_75t_L g418 ( .A1(n_327), .A2(n_404), .A3(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g408 ( .A(n_333), .Y(n_408) );
AND2x2_ASAP7_75t_L g421 ( .A(n_335), .B(n_344), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B(n_341), .Y(n_337) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_345), .B(n_448), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_355), .B1(n_357), .B2(n_358), .C(n_359), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_354), .A2(n_423), .B(n_425), .C(n_428), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_357), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g384 ( .A(n_365), .Y(n_384) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g370 ( .A(n_368), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_368), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B(n_378), .C(n_387), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_376), .A2(n_386), .B1(n_450), .B2(n_451), .C(n_453), .Y(n_449) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_382), .B2(n_385), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_SL g450 ( .A(n_389), .Y(n_450) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_422), .C(n_442), .D(n_449), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_398), .B(n_400), .C(n_418), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B(n_406), .C(n_410), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g429 ( .A(n_407), .Y(n_429) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
OR2x2_ASAP7_75t_L g440 ( .A(n_408), .B(n_441), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_432), .B2(n_434), .C(n_436), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_439), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g464 ( .A(n_458), .Y(n_464) );
NOR2x2_ASAP7_75t_L g767 ( .A(n_459), .B(n_474), .Y(n_767) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g473 ( .A(n_460), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g764 ( .A(n_469), .Y(n_764) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_478), .B(n_687), .Y(n_477) );
NOR5xp2_ASAP7_75t_L g478 ( .A(n_479), .B(n_600), .C(n_646), .D(n_659), .E(n_671), .Y(n_478) );
OAI211xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_514), .B(n_554), .C(n_581), .Y(n_479) );
INVx1_ASAP7_75t_SL g682 ( .A(n_480), .Y(n_682) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
AND2x2_ASAP7_75t_L g606 ( .A(n_481), .B(n_491), .Y(n_606) );
AND2x2_ASAP7_75t_L g634 ( .A(n_481), .B(n_580), .Y(n_634) );
AND2x2_ASAP7_75t_L g642 ( .A(n_481), .B(n_585), .Y(n_642) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g572 ( .A(n_482), .B(n_492), .Y(n_572) );
INVx2_ASAP7_75t_L g584 ( .A(n_482), .Y(n_584) );
AND2x2_ASAP7_75t_L g709 ( .A(n_482), .B(n_651), .Y(n_709) );
OR2x2_ASAP7_75t_L g711 ( .A(n_482), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g578 ( .A(n_483), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_487), .A2(n_499), .B(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_487), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_489), .A2(n_565), .B(n_568), .Y(n_564) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g622 ( .A(n_491), .B(n_594), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_491), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g736 ( .A(n_491), .B(n_576), .Y(n_736) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g626 ( .A(n_492), .Y(n_626) );
AND2x2_ASAP7_75t_L g651 ( .A(n_492), .B(n_563), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_492), .B(n_684), .Y(n_721) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g585 ( .A(n_493), .B(n_563), .Y(n_585) );
AND2x2_ASAP7_75t_L g599 ( .A(n_493), .B(n_562), .Y(n_599) );
AND2x2_ASAP7_75t_L g616 ( .A(n_493), .B(n_503), .Y(n_616) );
AND2x2_ASAP7_75t_L g673 ( .A(n_493), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_493), .B(n_580), .Y(n_686) );
AND2x2_ASAP7_75t_L g738 ( .A(n_493), .B(n_663), .Y(n_738) );
INVx2_ASAP7_75t_L g510 ( .A(n_501), .Y(n_510) );
AND2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g580 ( .A(n_503), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_503), .B(n_563), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_539), .B(n_551), .Y(n_514) );
INVx1_ASAP7_75t_SL g670 ( .A(n_515), .Y(n_670) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_529), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_517), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g553 ( .A(n_518), .Y(n_553) );
INVx1_ASAP7_75t_L g590 ( .A(n_518), .Y(n_590) );
AND2x2_ASAP7_75t_L g611 ( .A(n_518), .B(n_534), .Y(n_611) );
AND2x2_ASAP7_75t_L g645 ( .A(n_518), .B(n_535), .Y(n_645) );
OR2x2_ASAP7_75t_L g664 ( .A(n_518), .B(n_541), .Y(n_664) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_518), .Y(n_678) );
AND2x2_ASAP7_75t_L g691 ( .A(n_518), .B(n_692), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_523), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_529), .A2(n_613), .B1(n_614), .B2(n_623), .Y(n_612) );
AND2x2_ASAP7_75t_L g696 ( .A(n_529), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
INVx1_ASAP7_75t_L g557 ( .A(n_530), .Y(n_557) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_530), .Y(n_594) );
INVx1_ASAP7_75t_L g605 ( .A(n_530), .Y(n_605) );
AND2x2_ASAP7_75t_L g620 ( .A(n_530), .B(n_535), .Y(n_620) );
OR2x2_ASAP7_75t_L g574 ( .A(n_534), .B(n_559), .Y(n_574) );
AND2x2_ASAP7_75t_L g604 ( .A(n_534), .B(n_605), .Y(n_604) );
NOR2xp67_ASAP7_75t_L g692 ( .A(n_534), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g552 ( .A(n_535), .B(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g661 ( .A(n_535), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_539), .B(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g639 ( .A(n_540), .B(n_605), .Y(n_639) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g551 ( .A(n_541), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g610 ( .A(n_541), .Y(n_610) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g559 ( .A(n_542), .Y(n_559) );
OR2x2_ASAP7_75t_L g589 ( .A(n_542), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_542), .Y(n_644) );
AOI32xp33_ASAP7_75t_L g681 ( .A1(n_551), .A2(n_611), .A3(n_682), .B1(n_683), .B2(n_685), .Y(n_681) );
AND2x2_ASAP7_75t_L g607 ( .A(n_552), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_552), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_552), .B(n_639), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_552), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_560), .B1(n_573), .B2(n_575), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g660 ( .A(n_556), .B(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_557), .B(n_559), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_558), .A2(n_582), .B1(n_586), .B2(n_596), .Y(n_581) );
AND2x2_ASAP7_75t_L g603 ( .A(n_558), .B(n_604), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_558), .A2(n_572), .B(n_620), .C(n_655), .Y(n_654) );
OAI332xp33_ASAP7_75t_L g659 ( .A1(n_558), .A2(n_660), .A3(n_662), .B1(n_664), .B2(n_665), .B3(n_667), .C1(n_668), .C2(n_670), .Y(n_659) );
INVx2_ASAP7_75t_L g700 ( .A(n_558), .Y(n_700) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_559), .Y(n_618) );
INVx1_ASAP7_75t_L g693 ( .A(n_559), .Y(n_693) );
AND2x2_ASAP7_75t_L g747 ( .A(n_559), .B(n_611), .Y(n_747) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_572), .Y(n_560) );
AND2x2_ASAP7_75t_L g627 ( .A(n_562), .B(n_577), .Y(n_627) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g576 ( .A(n_563), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g675 ( .A(n_563), .B(n_577), .Y(n_675) );
INVx1_ASAP7_75t_L g684 ( .A(n_563), .Y(n_684) );
INVx1_ASAP7_75t_L g658 ( .A(n_572), .Y(n_658) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g742 ( .A(n_574), .B(n_594), .Y(n_742) );
INVx1_ASAP7_75t_SL g653 ( .A(n_575), .Y(n_653) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
AND2x2_ASAP7_75t_L g680 ( .A(n_576), .B(n_638), .Y(n_680) );
INVx1_ASAP7_75t_L g699 ( .A(n_576), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_576), .B(n_666), .Y(n_701) );
INVx1_ASAP7_75t_L g598 ( .A(n_577), .Y(n_598) );
AND2x2_ASAP7_75t_L g602 ( .A(n_579), .B(n_583), .Y(n_602) );
AND2x2_ASAP7_75t_L g669 ( .A(n_579), .B(n_627), .Y(n_669) );
INVx2_ASAP7_75t_L g712 ( .A(n_579), .Y(n_712) );
INVx2_ASAP7_75t_L g595 ( .A(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g597 ( .A(n_580), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g613 ( .A(n_583), .Y(n_613) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_584), .B(n_657), .Y(n_663) );
OR2x2_ASAP7_75t_L g727 ( .A(n_584), .B(n_686), .Y(n_727) );
INVx1_ASAP7_75t_L g751 ( .A(n_584), .Y(n_751) );
INVx1_ASAP7_75t_L g707 ( .A(n_585), .Y(n_707) );
AND2x2_ASAP7_75t_L g752 ( .A(n_585), .B(n_595), .Y(n_752) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_589), .A2(n_615), .B1(n_617), .B2(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI322xp33_ASAP7_75t_SL g698 ( .A1(n_592), .A2(n_699), .A3(n_700), .B1(n_701), .B2(n_702), .C1(n_705), .C2(n_707), .Y(n_698) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_L g695 ( .A(n_593), .B(n_611), .Y(n_695) );
OR2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g732 ( .A(n_593), .B(n_664), .Y(n_732) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g677 ( .A(n_594), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g733 ( .A(n_594), .B(n_664), .Y(n_733) );
INVx3_ASAP7_75t_L g666 ( .A(n_595), .Y(n_666) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g722 ( .A(n_597), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_599), .A2(n_602), .B1(n_603), .B2(n_606), .C1(n_607), .C2(n_609), .Y(n_601) );
INVx1_ASAP7_75t_L g632 ( .A(n_599), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_601), .B(n_612), .C(n_629), .Y(n_600) );
AND2x2_ASAP7_75t_L g717 ( .A(n_604), .B(n_618), .Y(n_717) );
BUFx2_ASAP7_75t_L g608 ( .A(n_605), .Y(n_608) );
INVx1_ASAP7_75t_L g649 ( .A(n_605), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_606), .A2(n_642), .B1(n_695), .B2(n_696), .C(n_698), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_608), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_611), .Y(n_635) );
AND2x2_ASAP7_75t_L g648 ( .A(n_611), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_616), .B(n_627), .Y(n_628) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_618), .A2(n_624), .B(n_628), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_618), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g715 ( .A(n_620), .B(n_697), .Y(n_715) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g638 ( .A(n_626), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_627), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g744 ( .A(n_627), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_635), .B1(n_636), .B2(n_639), .C(n_640), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_631), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g740 ( .A(n_639), .B(n_645), .Y(n_740) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OAI31xp33_ASAP7_75t_SL g708 ( .A1(n_643), .A2(n_682), .A3(n_709), .B(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g697 ( .A(n_644), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_645), .B(n_649), .Y(n_748) );
OAI221xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_650), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_646) );
INVx1_ASAP7_75t_L g652 ( .A(n_648), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_651), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g667 ( .A(n_660), .Y(n_667) );
INVx2_ASAP7_75t_L g703 ( .A(n_661), .Y(n_703) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g689 ( .A(n_666), .B(n_675), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_666), .A2(n_683), .B(n_740), .C(n_741), .Y(n_739) );
OAI221xp5_ASAP7_75t_SL g671 ( .A1(n_667), .A2(n_672), .B1(n_676), .B2(n_679), .C(n_681), .Y(n_671) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_670), .A2(n_735), .B(n_737), .C(n_739), .Y(n_734) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_673), .A2(n_724), .B1(n_726), .B2(n_728), .C(n_731), .Y(n_723) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
NOR4xp25_ASAP7_75t_L g687 ( .A(n_688), .B(n_713), .C(n_734), .D(n_745), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_690), .B(n_694), .C(n_708), .Y(n_688) );
INVx1_ASAP7_75t_SL g743 ( .A(n_695), .Y(n_743) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_SL g706 ( .A(n_704), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_711), .A2(n_720), .B1(n_732), .B2(n_733), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B(n_718), .C(n_723), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI31xp33_ASAP7_75t_L g745 ( .A1(n_716), .A2(n_746), .A3(n_748), .B(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
CKINVDCx14_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g761 ( .A(n_758), .Y(n_761) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx3_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
endmodule