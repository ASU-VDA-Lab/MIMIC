module real_jpeg_6574_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_1),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_1),
.A2(n_47),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_1),
.A2(n_47),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_1),
.B(n_119),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_1),
.A2(n_153),
.B(n_252),
.C(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_277),
.C(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_1),
.B(n_77),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_1),
.B(n_141),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_1),
.B(n_64),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_104),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_2),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_127),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_127),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_2),
.A2(n_127),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_3),
.Y(n_174)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_5),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_26),
.B1(n_36),
.B2(n_39),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_39),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_39),
.B1(n_102),
.B2(n_105),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_39),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_7),
.Y(n_116)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_7),
.Y(n_124)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_9),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_21),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_11),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_219),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_217),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_188),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_16),
.B(n_188),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.C(n_167),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_17),
.B(n_167),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_75),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_18),
.B(n_99),
.C(n_132),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_40),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_19),
.B(n_40),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_33),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_20),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_28),
.B(n_35),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_28),
.A2(n_171),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_28),
.B(n_171),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_28),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_33),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_33),
.B(n_285),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_37),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_69),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_41),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_42),
.Y(n_244)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_46),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_47),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_47),
.A2(n_148),
.B(n_197),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_47),
.A2(n_254),
.B(n_257),
.Y(n_253)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_49),
.B(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_50),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_51),
.B(n_70),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_51),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_51),
.B(n_265),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_64),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AO22x1_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_78)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_62),
.Y(n_267)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_64),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_64),
.B(n_265),
.Y(n_281)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_69),
.A2(n_181),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_69),
.B(n_264),
.Y(n_291)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_74),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_99),
.B1(n_132),
.B2(n_133),
.Y(n_75)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_94),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_77),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_77),
.B(n_160),
.Y(n_241)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_78),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_80),
.Y(n_256)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_81),
.Y(n_252)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_86),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_86),
.B(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_87),
.B(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_94),
.Y(n_158)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_125),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_119),
.Y(n_136)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_107),
.B(n_196),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_119),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_117),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_119),
.B(n_196),
.Y(n_195)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_125),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_144),
.A3(n_146),
.B1(n_147),
.B2(n_151),
.Y(n_143)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_134),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_155),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_135),
.B(n_155),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_138),
.B(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_143),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_159),
.B(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_179),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_169),
.B(n_284),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_178),
.B(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B(n_187),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_180),
.A2(n_214),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_180),
.B(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_187),
.B(n_281),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_188),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_208),
.CI(n_216),
.CON(n_188),
.SN(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_207),
.B(n_241),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_209),
.A2(n_215),
.B1(n_251),
.B2(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_337),
.B(n_350),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_269),
.B(n_336),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_246),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_222),
.B(n_246),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_231),
.B2(n_232),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_225),
.B(n_231),
.C(n_233),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.C(n_229),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_301),
.Y(n_313)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_234),
.B(n_237),
.C(n_243),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_260),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_247),
.B(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_250),
.A2(n_260),
.B1(n_261),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_250),
.Y(n_333)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_251),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_330),
.B(n_335),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_320),
.B(n_329),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_295),
.B(n_319),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_282),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_275),
.B1(n_280),
.B2(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_293),
.C(n_322),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_306),
.B(n_318),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_299),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_314),
.B(n_317),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_316),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_323),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_326),
.C(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_334),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_343),
.C(n_344),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_346),
.A2(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_347),
.B(n_349),
.Y(n_352)
);


endmodule