module fake_jpeg_3075_n_44 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

BUFx24_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_3),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_20),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_22),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_16),
.B(n_1),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_23),
.C(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_5),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_4),
.B(n_6),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_18),
.C(n_15),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_15),
.B1(n_10),
.B2(n_14),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_14),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_26),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

OAI211xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_36),
.B(n_12),
.C(n_10),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_26),
.B1(n_21),
.B2(n_12),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.Y(n_42)
);

OA21x2_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_14),
.B(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_9),
.C(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_39),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_42),
.B(n_39),
.Y(n_44)
);


endmodule