module fake_ariane_698_n_1824 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1824);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1824;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_33),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_104),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_79),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_60),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_42),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_93),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_140),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_94),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_16),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_82),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_137),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_95),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_37),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_42),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_143),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_18),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_43),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_133),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_99),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_29),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_87),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_38),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_146),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_109),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_78),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_145),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_11),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_48),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_38),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_127),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_121),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_37),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_7),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_17),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_88),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_161),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_72),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_160),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_168),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_116),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_101),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_175),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_98),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_126),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_136),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_49),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_110),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_170),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_114),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_15),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_45),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_174),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_162),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_40),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_53),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_112),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_113),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_41),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_152),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_64),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_67),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_31),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_76),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_128),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_61),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_130),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_181),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_69),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_8),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_52),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_173),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_89),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_158),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_124),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_134),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_153),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_10),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_163),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_25),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_58),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_103),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_5),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_90),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_106),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_3),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_4),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_108),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_25),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_10),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_115),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_19),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_32),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_75),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_169),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_131),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_1),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_81),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_155),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_166),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_125),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_83),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_4),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_91),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_165),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_39),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_47),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_3),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_77),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_43),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_179),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_167),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_92),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_157),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_15),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_58),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_52),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_117),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_8),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_51),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_118),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_2),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_46),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_62),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_132),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_22),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_138),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_147),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_96),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_24),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_23),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_80),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_50),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_71),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_2),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_12),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_16),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_360),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_194),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_242),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_300),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_0),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_319),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_264),
.B(n_0),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_264),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_6),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_226),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_280),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_R g376 ( 
.A(n_334),
.B(n_172),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_264),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_249),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_264),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_264),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_253),
.Y(n_382)
);

BUFx2_ASAP7_75t_SL g383 ( 
.A(n_294),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_322),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_264),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_264),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_294),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_294),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_328),
.B(n_6),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_189),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_351),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_264),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_295),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_352),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_230),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_186),
.B(n_7),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_204),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_234),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_295),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_295),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_252),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_257),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_266),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_308),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_272),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_230),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_283),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_9),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_329),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_260),
.B(n_345),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_349),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_231),
.B(n_9),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_184),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_184),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_296),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_353),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_304),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_220),
.B(n_11),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_235),
.B(n_13),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_214),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_230),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_325),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_185),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_185),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_330),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_187),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_187),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_214),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_224),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_224),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_189),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_220),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_188),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_230),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_R g439 ( 
.A(n_188),
.B(n_164),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_255),
.B(n_14),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_190),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_292),
.B(n_14),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_292),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_190),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_230),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_236),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_191),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_236),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_191),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_236),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_358),
.B(n_19),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_363),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_396),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_361),
.B(n_267),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_364),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_445),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_405),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_259),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_410),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_412),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_370),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_365),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_379),
.B(n_267),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_384),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_371),
.A2(n_357),
.B(n_289),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_417),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_361),
.B(n_267),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_386),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_391),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_395),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_414),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_422),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_383),
.B(n_277),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_414),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_431),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_379),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_438),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_436),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_R g495 ( 
.A(n_415),
.B(n_183),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_413),
.B(n_213),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_415),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_R g505 ( 
.A(n_425),
.B(n_207),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_425),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_387),
.B(n_192),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_426),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_433),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_426),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_428),
.B(n_267),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_367),
.B(n_227),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_418),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_428),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_369),
.B(n_378),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_429),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_429),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_446),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_437),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_227),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_387),
.B(n_299),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_479),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_470),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_479),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_479),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_478),
.B(n_458),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_492),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_501),
.B(n_441),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_411),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_453),
.B(n_362),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_479),
.B(n_441),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_458),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_529),
.A2(n_382),
.B1(n_409),
.B2(n_450),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_491),
.B(n_444),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_464),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_362),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_491),
.B(n_444),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_493),
.B(n_388),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_488),
.B(n_388),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_374),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_484),
.B(n_449),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_481),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_521),
.B(n_366),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_455),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_L g556 ( 
.A(n_500),
.B(n_201),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_478),
.B(n_374),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_478),
.B(n_394),
.Y(n_558)
);

NAND2x1p5_ASAP7_75t_L g559 ( 
.A(n_478),
.B(n_368),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_491),
.B(n_448),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_480),
.B(n_394),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_521),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_481),
.B(n_213),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_491),
.B(n_448),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_495),
.B(n_450),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_498),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_481),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_482),
.B(n_400),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_499),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_503),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_518),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_373),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_518),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_510),
.B(n_392),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_510),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_518),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_525),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_489),
.B(n_375),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_487),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_482),
.B(n_401),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_451),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_508),
.B(n_382),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_500),
.A2(n_440),
.B1(n_420),
.B2(n_389),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_454),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_502),
.B(n_419),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_456),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_460),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_505),
.B(n_375),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_512),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_525),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_502),
.B(n_401),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_506),
.B(n_442),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_485),
.B(n_390),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_506),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_460),
.B(n_274),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_514),
.B(n_435),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_520),
.B(n_303),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_507),
.B(n_452),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_490),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_518),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_522),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_500),
.A2(n_439),
.B1(n_356),
.B2(n_212),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_473),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_509),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_466),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_523),
.B(n_306),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_473),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_526),
.B(n_315),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_485),
.B(n_333),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_454),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_466),
.A2(n_376),
.B(n_337),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_500),
.A2(n_297),
.B1(n_267),
.B2(n_250),
.Y(n_618)
);

CKINVDCx16_ASAP7_75t_R g619 ( 
.A(n_467),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_500),
.B(n_193),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_500),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_517),
.A2(n_200),
.B1(n_197),
.B2(n_343),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_465),
.B(n_336),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_516),
.B(n_350),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_518),
.B(n_350),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_459),
.B(n_197),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_517),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_500),
.B(n_195),
.Y(n_628)
);

INVx6_ASAP7_75t_L g629 ( 
.A(n_518),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_528),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_475),
.A2(n_278),
.B1(n_274),
.B2(n_326),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_528),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_519),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_519),
.B(n_278),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_472),
.B(n_192),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_519),
.B(n_198),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_463),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_475),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_475),
.A2(n_527),
.B1(n_519),
.B2(n_496),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_468),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_463),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_519),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_527),
.B(n_198),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_200),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_527),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_527),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_527),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_473),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_475),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_463),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_496),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_476),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_454),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_516),
.B(n_199),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_497),
.B(n_343),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_454),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_454),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_454),
.B(n_326),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_494),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_494),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_461),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_477),
.A2(n_240),
.B1(n_182),
.B2(n_342),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_477),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_461),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_461),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_457),
.B(n_354),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_461),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_471),
.B(n_354),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_471),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_461),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_461),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_462),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_462),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_474),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_515),
.B(n_199),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_538),
.B(n_202),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_532),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_537),
.A2(n_324),
.B(n_228),
.C(n_233),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

BUFx8_ASAP7_75t_L g681 ( 
.A(n_640),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_592),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_587),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_538),
.B(n_202),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_653),
.B(n_483),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_626),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_550),
.B(n_206),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_558),
.B(n_210),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_535),
.A2(n_537),
.B1(n_541),
.B2(n_602),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_531),
.A2(n_462),
.B(n_347),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_626),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_596),
.B(n_203),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_660),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_588),
.A2(n_245),
.B1(n_275),
.B2(n_281),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_652),
.B(n_203),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_347),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_541),
.B(n_348),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_546),
.B(n_348),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_660),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_587),
.Y(n_700)
);

AND2x6_ASAP7_75t_SL g701 ( 
.A(n_601),
.B(n_524),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_542),
.A2(n_263),
.B1(n_291),
.B2(n_261),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_531),
.B(n_533),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_596),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_661),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_540),
.B(n_211),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_535),
.B(n_355),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_606),
.B(n_554),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_546),
.B(n_355),
.Y(n_709)
);

NOR2x1p5_ASAP7_75t_L g710 ( 
.A(n_584),
.B(n_217),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_535),
.B(n_218),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_574),
.Y(n_712)
);

BUFx6f_ASAP7_75t_SL g713 ( 
.A(n_675),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_545),
.B(n_222),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_661),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_618),
.A2(n_556),
.B1(n_600),
.B2(n_631),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_599),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_540),
.B(n_229),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_623),
.B(n_238),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_611),
.A2(n_243),
.B1(n_262),
.B2(n_341),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_607),
.B(n_256),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_591),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_614),
.B(n_305),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_561),
.B(n_307),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_556),
.B(n_196),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_534),
.B(n_309),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_604),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_644),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_667),
.B(n_310),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_554),
.B(n_513),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_557),
.A2(n_225),
.B1(n_241),
.B2(n_239),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_543),
.B(n_547),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_531),
.B(n_201),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_669),
.B(n_312),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_669),
.B(n_317),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_591),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_562),
.A2(n_663),
.B1(n_548),
.B2(n_656),
.C(n_598),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_544),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_610),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_SL g741 ( 
.A(n_565),
.B(n_332),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_568),
.B(n_335),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_543),
.A2(n_216),
.B1(n_219),
.B2(n_215),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_579),
.B(n_462),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_547),
.B(n_339),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_609),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_583),
.B(n_340),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_613),
.B(n_208),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_560),
.B(n_20),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_627),
.B(n_630),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_632),
.B(n_562),
.Y(n_751)
);

NOR2x1p5_ASAP7_75t_L g752 ( 
.A(n_584),
.B(n_209),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_560),
.A2(n_276),
.B1(n_331),
.B2(n_327),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_644),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_539),
.B(n_221),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_564),
.B(n_20),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_600),
.A2(n_462),
.B1(n_205),
.B2(n_196),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_564),
.A2(n_279),
.B1(n_323),
.B2(n_321),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_597),
.B(n_603),
.Y(n_759)
);

NOR2x1p5_ASAP7_75t_L g760 ( 
.A(n_585),
.B(n_656),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_598),
.A2(n_270),
.B1(n_318),
.B2(n_316),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_622),
.A2(n_268),
.B1(n_314),
.B2(n_311),
.C(n_301),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_615),
.A2(n_258),
.B(n_298),
.C(n_293),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_610),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_637),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_565),
.B(n_254),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_597),
.B(n_265),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_574),
.A2(n_251),
.B1(n_290),
.B2(n_287),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_551),
.A2(n_247),
.B1(n_286),
.B2(n_285),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_559),
.B(n_21),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_544),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_566),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_570),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_555),
.B(n_196),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_603),
.B(n_284),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_571),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_559),
.B(n_21),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_636),
.A2(n_22),
.B(n_23),
.C(n_26),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_549),
.B(n_282),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_585),
.B(n_244),
.C(n_269),
.Y(n_780)
);

INVx8_ASAP7_75t_L g781 ( 
.A(n_574),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_641),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_549),
.B(n_232),
.Y(n_783)
);

BUFx5_ASAP7_75t_L g784 ( 
.A(n_621),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_549),
.B(n_26),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_SL g786 ( 
.A(n_675),
.B(n_237),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_619),
.B(n_27),
.Y(n_787)
);

BUFx2_ASAP7_75t_R g788 ( 
.A(n_593),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_533),
.A2(n_223),
.B1(n_246),
.B2(n_248),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_651),
.Y(n_790)
);

AO22x1_ASAP7_75t_L g791 ( 
.A1(n_536),
.A2(n_271),
.B1(n_196),
.B2(n_205),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_600),
.A2(n_620),
.B1(n_628),
.B2(n_567),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_676),
.A2(n_273),
.B1(n_201),
.B2(n_205),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_572),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_590),
.B(n_273),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_594),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_600),
.A2(n_205),
.B1(n_196),
.B2(n_201),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_594),
.B(n_635),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_578),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_577),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_651),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_553),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_594),
.B(n_205),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_590),
.B(n_27),
.Y(n_804)
);

NAND2x1_ASAP7_75t_L g805 ( 
.A(n_533),
.B(n_273),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_590),
.B(n_273),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_580),
.B(n_273),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_552),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_553),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_595),
.B(n_273),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_617),
.A2(n_273),
.B1(n_201),
.B2(n_34),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_567),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_577),
.B(n_273),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_574),
.B(n_201),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_617),
.B(n_664),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_593),
.B(n_617),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_664),
.B(n_201),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_579),
.B(n_30),
.Y(n_818)
);

AND2x6_ASAP7_75t_SL g819 ( 
.A(n_675),
.B(n_655),
.Y(n_819)
);

INVx8_ASAP7_75t_L g820 ( 
.A(n_600),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_534),
.B(n_201),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_534),
.B(n_30),
.Y(n_822)
);

BUFx6f_ASAP7_75t_SL g823 ( 
.A(n_624),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_643),
.B(n_32),
.C(n_34),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_621),
.B(n_35),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_534),
.B(n_621),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_534),
.B(n_35),
.C(n_36),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_670),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_638),
.B(n_36),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_633),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_600),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_638),
.B(n_650),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_639),
.A2(n_74),
.B(n_150),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_650),
.B(n_49),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_563),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_648),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_704),
.B(n_624),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_686),
.B(n_575),
.Y(n_838)
);

NOR2x1p5_ASAP7_75t_L g839 ( 
.A(n_796),
.B(n_575),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_708),
.B(n_569),
.Y(n_840)
);

OAI321xp33_ASAP7_75t_L g841 ( 
.A1(n_831),
.A2(n_625),
.A3(n_634),
.B1(n_659),
.B2(n_646),
.C(n_647),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_733),
.B(n_648),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_712),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_749),
.A2(n_569),
.B1(n_608),
.B2(n_586),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_765),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_734),
.A2(n_649),
.B(n_586),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_734),
.A2(n_649),
.B(n_586),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_760),
.A2(n_629),
.B1(n_625),
.B2(n_642),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_733),
.B(n_649),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_826),
.A2(n_575),
.B(n_608),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_691),
.B(n_608),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_678),
.B(n_612),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_800),
.B(n_612),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_826),
.A2(n_612),
.B(n_668),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_829),
.A2(n_645),
.B(n_634),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_749),
.A2(n_629),
.B1(n_658),
.B2(n_668),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_714),
.B(n_665),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_805),
.A2(n_666),
.B(n_658),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_717),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_689),
.B(n_573),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_832),
.A2(n_666),
.B(n_658),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_834),
.A2(n_659),
.B(n_674),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_756),
.A2(n_668),
.B(n_666),
.C(n_665),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_750),
.A2(n_665),
.B(n_654),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_725),
.A2(n_654),
.B(n_671),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_742),
.A2(n_654),
.B(n_671),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_756),
.A2(n_673),
.B(n_672),
.C(n_662),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_764),
.A2(n_672),
.B(n_673),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_688),
.B(n_573),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_770),
.B(n_573),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_688),
.B(n_573),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_702),
.A2(n_662),
.B(n_55),
.C(n_56),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_800),
.B(n_677),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_718),
.Y(n_874)
);

INVx11_ASAP7_75t_L g875 ( 
.A(n_681),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_684),
.B(n_605),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_706),
.A2(n_605),
.B(n_576),
.C(n_657),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_712),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_720),
.B(n_605),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_738),
.B(n_54),
.C(n_57),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_731),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_820),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_747),
.A2(n_605),
.B(n_576),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_759),
.B(n_576),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_706),
.A2(n_657),
.B(n_616),
.C(n_589),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_719),
.A2(n_657),
.B(n_616),
.C(n_589),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_719),
.B(n_563),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_695),
.A2(n_657),
.B(n_616),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_771),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_696),
.A2(n_657),
.B(n_616),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_745),
.B(n_563),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_739),
.B(n_729),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_745),
.A2(n_563),
.B1(n_616),
.B2(n_589),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_751),
.B(n_563),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_818),
.A2(n_589),
.B(n_63),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_712),
.B(n_59),
.Y(n_896)
);

INVx11_ASAP7_75t_L g897 ( 
.A(n_681),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_820),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_746),
.B(n_65),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_804),
.B(n_84),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_833),
.A2(n_85),
.B(n_86),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_770),
.A2(n_105),
.B(n_107),
.C(n_123),
.Y(n_902)
);

INVx3_ASAP7_75t_SL g903 ( 
.A(n_685),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_726),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_777),
.A2(n_726),
.B1(n_816),
.B2(n_754),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_R g907 ( 
.A(n_786),
.B(n_713),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_821),
.A2(n_815),
.B(n_817),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_718),
.B(n_728),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_830),
.A2(n_748),
.B(n_690),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_804),
.B(n_752),
.Y(n_911)
);

AOI33xp33_ASAP7_75t_L g912 ( 
.A1(n_835),
.A2(n_831),
.A3(n_785),
.B1(n_762),
.B2(n_679),
.B3(n_778),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_683),
.A2(n_737),
.B(n_700),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_723),
.A2(n_740),
.B(n_755),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_716),
.A2(n_680),
.B1(n_682),
.B2(n_835),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_768),
.B(n_777),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_692),
.B(n_707),
.C(n_780),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_730),
.B(n_735),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_698),
.A2(n_709),
.B(n_697),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_736),
.B(n_693),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_728),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_685),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_836),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_816),
.A2(n_768),
.B1(n_798),
.B2(n_721),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_744),
.A2(n_766),
.B(n_812),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_710),
.B(n_685),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_699),
.B(n_705),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_807),
.A2(n_810),
.B(n_795),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_769),
.B(n_694),
.C(n_732),
.Y(n_929)
);

BUFx4f_ASAP7_75t_L g930 ( 
.A(n_781),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_715),
.B(n_773),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_724),
.B(n_781),
.Y(n_932)
);

AO21x1_ASAP7_75t_L g933 ( 
.A1(n_811),
.A2(n_818),
.B(n_793),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_767),
.B(n_775),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_789),
.A2(n_722),
.B1(n_774),
.B2(n_741),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_744),
.A2(n_802),
.B(n_809),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_781),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_772),
.B(n_794),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_819),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_776),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_L g941 ( 
.A(n_779),
.B(n_783),
.C(n_711),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_808),
.B(n_774),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_716),
.A2(n_797),
.B1(n_827),
.B2(n_825),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_799),
.B(n_813),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_782),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_787),
.B(n_824),
.C(n_763),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_828),
.B(n_761),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_790),
.A2(n_801),
.B(n_822),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_743),
.B(n_753),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_L g950 ( 
.A(n_758),
.B(n_824),
.C(n_727),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_806),
.A2(n_792),
.B(n_803),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_823),
.B(n_788),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_784),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_814),
.A2(n_792),
.B(n_797),
.C(n_757),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_823),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_791),
.B(n_757),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_713),
.B(n_701),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_784),
.A2(n_749),
.B1(n_756),
.B2(n_726),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_784),
.B(n_708),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_784),
.B(n_708),
.Y(n_960)
);

OAI321xp33_ASAP7_75t_L g961 ( 
.A1(n_784),
.A2(n_831),
.A3(n_835),
.B1(n_811),
.B2(n_756),
.C(n_749),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_784),
.A2(n_704),
.B(n_537),
.C(n_749),
.Y(n_962)
);

CKINVDCx16_ASAP7_75t_R g963 ( 
.A(n_713),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_760),
.A2(n_756),
.B1(n_749),
.B2(n_704),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_733),
.A2(n_704),
.B1(n_714),
.B2(n_716),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_687),
.B(n_538),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_687),
.B(n_538),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_687),
.B(n_538),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_796),
.B(n_820),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_687),
.B(n_538),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_L g975 ( 
.A1(n_725),
.A2(n_747),
.B(n_742),
.C(n_540),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_765),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_733),
.A2(n_704),
.B1(n_714),
.B2(n_716),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_687),
.B(n_538),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_749),
.A2(n_756),
.B(n_733),
.C(n_706),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_678),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_749),
.A2(n_756),
.B(n_733),
.C(n_706),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_689),
.B(n_768),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_704),
.A2(n_537),
.B(n_756),
.C(n_749),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_689),
.B(n_768),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_678),
.B(n_453),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_713),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_678),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_687),
.B(n_538),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_717),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_765),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_717),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_765),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_804),
.B(n_680),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_687),
.B(n_538),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_678),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_765),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_704),
.A2(n_537),
.B(n_756),
.C(n_749),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_749),
.A2(n_756),
.B1(n_726),
.B2(n_733),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_712),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_749),
.A2(n_756),
.B1(n_726),
.B2(n_733),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_687),
.B(n_538),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_678),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_689),
.B(n_768),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_703),
.A2(n_734),
.B(n_826),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_704),
.A2(n_537),
.B(n_756),
.C(n_749),
.Y(n_1008)
);

BUFx8_ASAP7_75t_L g1009 ( 
.A(n_713),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_712),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_733),
.A2(n_834),
.B(n_829),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_968),
.B(n_969),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_859),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_889),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_948),
.A2(n_928),
.B(n_862),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_909),
.B(n_881),
.Y(n_1018)
);

OAI22x1_ASAP7_75t_L g1019 ( 
.A1(n_965),
.A2(n_916),
.B1(n_924),
.B2(n_985),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_862),
.A2(n_855),
.B(n_951),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_875),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_970),
.B(n_973),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_958),
.A2(n_856),
.B(n_1001),
.Y(n_1023)
);

AO31x2_ASAP7_75t_L g1024 ( 
.A1(n_933),
.A2(n_901),
.A3(n_1001),
.B(n_1003),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_980),
.A2(n_1008),
.B(n_984),
.C(n_1000),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_869),
.A2(n_871),
.B(n_919),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_978),
.B(n_989),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_921),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_996),
.B(n_1004),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_1009),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_868),
.A2(n_966),
.B(n_964),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_873),
.B(n_918),
.Y(n_1032)
);

CKINVDCx11_ASAP7_75t_R g1033 ( 
.A(n_903),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_897),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_971),
.A2(n_979),
.B(n_974),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_882),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_929),
.B(n_880),
.C(n_1003),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_849),
.A2(n_842),
.B(n_967),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_960),
.B(n_840),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_874),
.B(n_942),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_905),
.A2(n_977),
.B1(n_983),
.B2(n_1006),
.Y(n_1041)
);

AO31x2_ASAP7_75t_L g1042 ( 
.A1(n_958),
.A2(n_915),
.A3(n_943),
.B(n_954),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_868),
.A2(n_1007),
.B(n_997),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_992),
.A2(n_867),
.B(n_910),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_857),
.A2(n_879),
.B(n_962),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_990),
.B(n_993),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_1010),
.B(n_843),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_853),
.B(n_920),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_995),
.B(n_896),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_892),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_930),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_988),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_922),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_863),
.A2(n_953),
.B(n_861),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_998),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_853),
.B(n_938),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_953),
.A2(n_856),
.B(n_925),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_936),
.A2(n_888),
.B(n_890),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_914),
.A2(n_854),
.B(n_883),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_934),
.A2(n_944),
.B(n_876),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_911),
.B(n_926),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_940),
.B(n_838),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_851),
.B(n_837),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_913),
.A2(n_850),
.B(n_847),
.Y(n_1064)
);

OAI222xp33_ASAP7_75t_L g1065 ( 
.A1(n_943),
.A2(n_896),
.B1(n_904),
.B2(n_900),
.C1(n_935),
.C2(n_961),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_882),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_846),
.A2(n_899),
.B(n_891),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_961),
.A2(n_950),
.B(n_947),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_945),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_975),
.A2(n_886),
.B(n_885),
.C(n_877),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_1010),
.B(n_930),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_887),
.A2(n_860),
.B(n_844),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_844),
.A2(n_864),
.B(n_858),
.Y(n_1073)
);

AOI21x1_ASAP7_75t_L g1074 ( 
.A1(n_894),
.A2(n_884),
.B(n_866),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_976),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_907),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_898),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_865),
.A2(n_893),
.B(n_904),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_995),
.B(n_852),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_912),
.A2(n_872),
.B(n_946),
.C(n_902),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_852),
.B(n_870),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_931),
.A2(n_941),
.B(n_841),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_991),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_1009),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_870),
.B(n_1005),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_911),
.A2(n_932),
.B1(n_986),
.B2(n_917),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_981),
.A2(n_927),
.B(n_923),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_841),
.B(n_906),
.Y(n_1088)
);

BUFx12f_ASAP7_75t_L g1089 ( 
.A(n_987),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_994),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_937),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_956),
.A2(n_898),
.B(n_906),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_999),
.A2(n_955),
.A3(n_957),
.B(n_952),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_972),
.A2(n_848),
.B(n_923),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_937),
.A2(n_896),
.B(n_843),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_839),
.A2(n_843),
.B(n_878),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_939),
.A2(n_878),
.B(n_1002),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_878),
.A2(n_939),
.B(n_963),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_939),
.A2(n_908),
.B(n_1011),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_939),
.A2(n_908),
.B(n_1011),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_845),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_909),
.B(n_708),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_909),
.B(n_708),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_968),
.B(n_969),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_980),
.A2(n_982),
.B(n_1011),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_909),
.B(n_708),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_909),
.B(n_708),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_968),
.B(n_969),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_921),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_980),
.A2(n_982),
.B(n_1011),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_889),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_968),
.B(n_969),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_1009),
.Y(n_1124)
);

AOI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_949),
.A2(n_532),
.B(n_984),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_968),
.B(n_969),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_875),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_968),
.B(n_969),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_845),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_843),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_875),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_968),
.B(n_969),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_875),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_980),
.A2(n_982),
.B(n_1011),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_908),
.A2(n_958),
.B(n_856),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1140)
);

OAI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_968),
.A2(n_601),
.B(n_969),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_980),
.B(n_982),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_968),
.B(n_969),
.Y(n_1143)
);

BUFx8_ASAP7_75t_L g1144 ( 
.A(n_922),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_968),
.B(n_969),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_921),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_968),
.B(n_969),
.Y(n_1148)
);

BUFx4f_ASAP7_75t_L g1149 ( 
.A(n_903),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_SL g1150 ( 
.A1(n_965),
.A2(n_601),
.B(n_542),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_895),
.A2(n_1011),
.B(n_982),
.Y(n_1153)
);

AOI221x1_ASAP7_75t_L g1154 ( 
.A1(n_1001),
.A2(n_1003),
.B1(n_980),
.B2(n_982),
.C(n_880),
.Y(n_1154)
);

AOI21x1_ASAP7_75t_L g1155 ( 
.A1(n_908),
.A2(n_958),
.B(n_856),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_968),
.B(n_969),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_908),
.A2(n_1011),
.B(n_895),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_895),
.A2(n_1000),
.B(n_984),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1146),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1146),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1030),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1013),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1150),
.A2(n_1027),
.B1(n_1037),
.B2(n_1138),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1065),
.B(n_1041),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1027),
.A2(n_1119),
.B1(n_1111),
.B2(n_1108),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1016),
.A2(n_1126),
.B1(n_1102),
.B2(n_1153),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_1051),
.B(n_1091),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_L g1168 ( 
.A(n_1141),
.B(n_1012),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1107),
.B(n_1109),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_L g1170 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1014),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1110),
.B(n_1116),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1047),
.B(n_1097),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1030),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1113),
.B(n_1114),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1080),
.A2(n_1025),
.B(n_1142),
.C(n_1158),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1124),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1049),
.B(n_1095),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1104),
.A2(n_1137),
.B(n_1152),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1112),
.A2(n_1132),
.B(n_1151),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_1021),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1061),
.B(n_1097),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1125),
.A2(n_1068),
.B(n_1123),
.C(n_1147),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1021),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1140),
.A2(n_1142),
.B(n_1038),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1149),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1122),
.B(n_1127),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1071),
.Y(n_1188)
);

OAI21xp33_ASAP7_75t_L g1189 ( 
.A1(n_1080),
.A2(n_1145),
.B(n_1156),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1045),
.A2(n_1026),
.B(n_1025),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1071),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1133),
.B(n_1096),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1143),
.Y(n_1193)
);

CKINVDCx8_ASAP7_75t_R g1194 ( 
.A(n_1084),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1028),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1135),
.B(n_1032),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1133),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1018),
.B(n_1050),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1133),
.B(n_1076),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1040),
.B(n_1121),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1033),
.Y(n_1201)
);

AO32x1_ASAP7_75t_L g1202 ( 
.A1(n_1154),
.A2(n_1024),
.A3(n_1042),
.B1(n_1023),
.B2(n_1131),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1046),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1035),
.A2(n_1078),
.B(n_1157),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1133),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1036),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1078),
.A2(n_1015),
.B(n_1128),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_1034),
.B(n_1129),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1062),
.A2(n_1056),
.B1(n_1039),
.B2(n_1048),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1015),
.A2(n_1157),
.B(n_1101),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1082),
.B(n_1063),
.C(n_1086),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1019),
.A2(n_1069),
.B1(n_1090),
.B2(n_1131),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1042),
.B(n_1060),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1117),
.B(n_1052),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1075),
.Y(n_1215)
);

AOI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1088),
.A2(n_1118),
.B(n_1105),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1079),
.B(n_1098),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1085),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1105),
.A2(n_1106),
.B(n_1115),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_SL g1220 ( 
.A(n_1081),
.B(n_1088),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1115),
.A2(n_1118),
.B(n_1128),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1094),
.A2(n_1042),
.B1(n_1155),
.B2(n_1139),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1042),
.B(n_1024),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1036),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1024),
.B(n_1103),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1024),
.B(n_1103),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1074),
.A2(n_1072),
.B(n_1017),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1055),
.B(n_1087),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1083),
.B(n_1090),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1134),
.B(n_1136),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1033),
.B(n_1084),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1053),
.A2(n_1144),
.B1(n_1089),
.B2(n_1124),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1066),
.B(n_1077),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1066),
.B(n_1077),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1120),
.A2(n_1073),
.B(n_1057),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1093),
.B(n_1089),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1099),
.B(n_1100),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1053),
.A2(n_1144),
.B1(n_1100),
.B2(n_1099),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1073),
.A2(n_1057),
.B(n_1070),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1053),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1020),
.A2(n_1144),
.B1(n_1031),
.B2(n_1043),
.Y(n_1241)
);

CKINVDCx6p67_ASAP7_75t_R g1242 ( 
.A(n_1093),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1058),
.A2(n_1067),
.B(n_1044),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1093),
.B(n_1092),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1092),
.B(n_1031),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1054),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1064),
.B(n_1059),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1059),
.A2(n_363),
.B1(n_370),
.B2(n_364),
.Y(n_1248)
);

AND2x6_ASAP7_75t_L g1249 ( 
.A(n_1058),
.B(n_959),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1150),
.B(n_544),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1013),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1107),
.B(n_1109),
.Y(n_1252)
);

AOI222xp33_ASAP7_75t_L g1253 ( 
.A1(n_1150),
.A2(n_1065),
.B1(n_916),
.B2(n_970),
.C1(n_973),
.C2(n_969),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1111),
.A2(n_1138),
.B(n_1119),
.C(n_581),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1016),
.A2(n_982),
.B(n_980),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1047),
.B(n_1010),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1056),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1107),
.B(n_1109),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1146),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1146),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1071),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1047),
.B(n_1010),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1149),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1047),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1049),
.B(n_1095),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1269)
);

INVx3_ASAP7_75t_SL g1270 ( 
.A(n_1084),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1016),
.A2(n_1104),
.B(n_1102),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1027),
.A2(n_1000),
.B(n_1008),
.C(n_984),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1150),
.A2(n_982),
.B1(n_980),
.B2(n_965),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1013),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1027),
.A2(n_1000),
.B(n_1008),
.C(n_984),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1013),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1047),
.B(n_1010),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1071),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1021),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1283)
);

CKINVDCx11_ASAP7_75t_R g1284 ( 
.A(n_1030),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1013),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1047),
.B(n_1010),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1107),
.B(n_1109),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1027),
.A2(n_969),
.B1(n_973),
.B2(n_970),
.C(n_968),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1284),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1171),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1174),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1200),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1174),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1164),
.A2(n_1253),
.B1(n_1163),
.B2(n_1288),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1192),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1164),
.A2(n_1253),
.B1(n_1273),
.B2(n_1250),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1282),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1214),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1249),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1260),
.A2(n_1263),
.B1(n_1276),
.B2(n_1277),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1273),
.A2(n_1248),
.B1(n_1189),
.B2(n_1168),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1165),
.B(n_1255),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1267),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1251),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1267),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1216),
.A2(n_1183),
.B(n_1225),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1179),
.A2(n_1271),
.B(n_1180),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1159),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1160),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1261),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1176),
.A2(n_1209),
.B(n_1255),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1170),
.A2(n_1209),
.B1(n_1277),
.B2(n_1260),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_1205),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1274),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1195),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1263),
.A2(n_1280),
.B1(n_1269),
.B2(n_1265),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1278),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1227),
.A2(n_1190),
.B(n_1241),
.Y(n_1319)
);

BUFx4f_ASAP7_75t_SL g1320 ( 
.A(n_1161),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1194),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1285),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1211),
.A2(n_1280),
.B1(n_1269),
.B2(n_1265),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1216),
.A2(n_1226),
.B(n_1225),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1177),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1215),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1223),
.B(n_1169),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1223),
.B(n_1175),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1259),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1272),
.A2(n_1275),
.B(n_1193),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1276),
.A2(n_1283),
.B1(n_1287),
.B2(n_1258),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1283),
.A2(n_1196),
.B1(n_1187),
.B2(n_1198),
.Y(n_1332)
);

INVx8_ASAP7_75t_L g1333 ( 
.A(n_1178),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1256),
.B(n_1264),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1249),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1187),
.A2(n_1196),
.B1(n_1185),
.B2(n_1252),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1243),
.A2(n_1239),
.B(n_1204),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1270),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1267),
.Y(n_1339)
);

BUFx2_ASAP7_75t_R g1340 ( 
.A(n_1201),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1235),
.A2(n_1219),
.B(n_1221),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1172),
.A2(n_1236),
.B1(n_1203),
.B2(n_1257),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1228),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1231),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1229),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1249),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1233),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1182),
.A2(n_1199),
.B1(n_1186),
.B2(n_1266),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1229),
.Y(n_1349)
);

CKINVDCx11_ASAP7_75t_R g1350 ( 
.A(n_1181),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1240),
.A2(n_1268),
.B1(n_1178),
.B2(n_1238),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1226),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_SL g1353 ( 
.A(n_1181),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_1213),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1256),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1230),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1220),
.A2(n_1268),
.B1(n_1178),
.B2(n_1218),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1264),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1241),
.A2(n_1210),
.B(n_1247),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1233),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1184),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1234),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1244),
.Y(n_1363)
);

CKINVDCx14_ASAP7_75t_R g1364 ( 
.A(n_1184),
.Y(n_1364)
);

BUFx2_ASAP7_75t_R g1365 ( 
.A(n_1188),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1166),
.A2(n_1207),
.B(n_1222),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1268),
.A2(n_1188),
.B1(n_1191),
.B2(n_1262),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1279),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1234),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1218),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1206),
.A2(n_1224),
.B1(n_1254),
.B2(n_1208),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1212),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1213),
.B(n_1173),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1279),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1197),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1249),
.Y(n_1376)
);

BUFx5_ASAP7_75t_L g1377 ( 
.A(n_1246),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1167),
.A2(n_1206),
.B(n_1224),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1237),
.A2(n_1245),
.B(n_1217),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1202),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1286),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1217),
.Y(n_1382)
);

AND2x2_ASAP7_75t_SL g1383 ( 
.A(n_1232),
.B(n_1286),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1242),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1197),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1281),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1202),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1202),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1284),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1171),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1249),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1171),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1256),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1164),
.A2(n_1150),
.B1(n_965),
.B2(n_916),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1249),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1162),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1379),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1379),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1379),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1366),
.A2(n_1319),
.B(n_1341),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1352),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1303),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1303),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1354),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1324),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1387),
.A2(n_1388),
.B(n_1380),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1380),
.A2(n_1330),
.B(n_1359),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1326),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1345),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1301),
.B(n_1313),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1292),
.B(n_1391),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1349),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1373),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1373),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1292),
.B(n_1391),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1347),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1360),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1307),
.A2(n_1351),
.B(n_1395),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1362),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1369),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1333),
.B(n_1300),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1372),
.A2(n_1312),
.B(n_1397),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1342),
.A2(n_1295),
.B(n_1363),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1309),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_L g1428 ( 
.A(n_1336),
.B(n_1335),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1295),
.A2(n_1297),
.B1(n_1302),
.B2(n_1317),
.C(n_1323),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1343),
.B(n_1331),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1335),
.B(n_1346),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1305),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1315),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1316),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1318),
.B(n_1322),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1370),
.A2(n_1367),
.B(n_1384),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1382),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1323),
.B(n_1332),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1293),
.B(n_1310),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1342),
.A2(n_1297),
.B(n_1302),
.Y(n_1440)
);

AO21x1_ASAP7_75t_L g1441 ( 
.A1(n_1371),
.A2(n_1378),
.B(n_1348),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1376),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1290),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1337),
.A2(n_1308),
.B(n_1396),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1392),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1392),
.Y(n_1446)
);

BUFx4f_ASAP7_75t_SL g1447 ( 
.A(n_1289),
.Y(n_1447)
);

BUFx2_ASAP7_75t_SL g1448 ( 
.A(n_1361),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1311),
.B(n_1299),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1396),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1390),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1377),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1377),
.B(n_1296),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1296),
.A2(n_1375),
.B(n_1386),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1377),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1386),
.A2(n_1329),
.B(n_1393),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1383),
.A2(n_1314),
.B(n_1353),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1403),
.B(n_1356),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1413),
.B(n_1353),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1413),
.A2(n_1333),
.B(n_1357),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1405),
.B(n_1385),
.Y(n_1461)
);

BUFx4f_ASAP7_75t_SL g1462 ( 
.A(n_1443),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1406),
.B(n_1314),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1411),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1406),
.B(n_1314),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1454),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1429),
.A2(n_1334),
.B1(n_1368),
.B2(n_1358),
.C(n_1374),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1404),
.B(n_1333),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1411),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1454),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1414),
.B(n_1383),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1406),
.B(n_1364),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1404),
.B(n_1430),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1431),
.B(n_1368),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1414),
.B(n_1364),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1438),
.B(n_1361),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1414),
.B(n_1339),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1429),
.A2(n_1289),
.B1(n_1389),
.B2(n_1333),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1418),
.B(n_1306),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1398),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1418),
.B(n_1306),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1418),
.B(n_1306),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1440),
.A2(n_1389),
.B1(n_1394),
.B2(n_1381),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1398),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1454),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1419),
.B(n_1304),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1454),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1399),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1454),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1398),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1399),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1416),
.B(n_1417),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1430),
.B(n_1409),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1400),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1447),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1440),
.A2(n_1438),
.B1(n_1421),
.B2(n_1426),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1425),
.B(n_1355),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_SL g1498 ( 
.A(n_1441),
.B(n_1344),
.C(n_1294),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1400),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1478),
.A2(n_1440),
.B1(n_1428),
.B2(n_1434),
.Y(n_1500)
);

NAND4xp25_ASAP7_75t_L g1501 ( 
.A(n_1476),
.B(n_1443),
.C(n_1451),
.D(n_1427),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1496),
.B(n_1427),
.C(n_1440),
.Y(n_1502)
);

NAND4xp25_ASAP7_75t_L g1503 ( 
.A(n_1498),
.B(n_1476),
.C(n_1478),
.D(n_1459),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1434),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1459),
.A2(n_1440),
.B1(n_1428),
.B2(n_1448),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1475),
.B(n_1417),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1475),
.B(n_1453),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1462),
.B(n_1441),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1458),
.B(n_1449),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1462),
.B(n_1457),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1475),
.B(n_1453),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1467),
.A2(n_1471),
.B1(n_1483),
.B2(n_1460),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1496),
.B(n_1422),
.C(n_1420),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1495),
.B(n_1340),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1472),
.B(n_1453),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1467),
.A2(n_1448),
.B1(n_1344),
.B2(n_1442),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1498),
.A2(n_1472),
.B(n_1483),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1460),
.A2(n_1421),
.B1(n_1426),
.B2(n_1436),
.Y(n_1520)
);

NAND4xp25_ASAP7_75t_L g1521 ( 
.A(n_1472),
.B(n_1433),
.C(n_1432),
.D(n_1435),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1463),
.B(n_1409),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1463),
.B(n_1409),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1466),
.A2(n_1401),
.B(n_1444),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1493),
.B(n_1422),
.C(n_1420),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1471),
.A2(n_1457),
.B1(n_1426),
.B2(n_1424),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1493),
.A2(n_1442),
.B(n_1456),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1463),
.B(n_1409),
.Y(n_1528)
);

NAND4xp25_ASAP7_75t_L g1529 ( 
.A(n_1493),
.B(n_1433),
.C(n_1435),
.D(n_1423),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1492),
.B(n_1423),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1465),
.B(n_1410),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1465),
.B(n_1410),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1492),
.B(n_1465),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1477),
.B(n_1479),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1474),
.B(n_1456),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1477),
.B(n_1410),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1492),
.B(n_1425),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1477),
.B(n_1425),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1468),
.A2(n_1446),
.B1(n_1450),
.B2(n_1445),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1464),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1497),
.A2(n_1421),
.B1(n_1426),
.B2(n_1436),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1479),
.B(n_1410),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1479),
.B(n_1425),
.Y(n_1543)
);

NAND4xp25_ASAP7_75t_L g1544 ( 
.A(n_1461),
.B(n_1455),
.C(n_1452),
.D(n_1412),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1481),
.B(n_1407),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1481),
.B(n_1482),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1481),
.B(n_1407),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1482),
.B(n_1452),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1466),
.A2(n_1412),
.B1(n_1415),
.B2(n_1402),
.C(n_1408),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_1486),
.B(n_1408),
.C(n_1437),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1540),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1522),
.B(n_1490),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1537),
.B(n_1488),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1522),
.B(n_1490),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1470),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1524),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1524),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1524),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1549),
.B(n_1488),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1523),
.B(n_1470),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1531),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1540),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1538),
.B(n_1491),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1531),
.B(n_1480),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1532),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1509),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1536),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1532),
.B(n_1485),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1534),
.B(n_1485),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1534),
.B(n_1487),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1524),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1516),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1504),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1525),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_R g1575 ( 
.A(n_1520),
.B(n_1291),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1542),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1525),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_1543),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1487),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1550),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1530),
.B(n_1494),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1545),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1547),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1508),
.B(n_1489),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1508),
.B(n_1489),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1527),
.B(n_1494),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1515),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1515),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1513),
.B(n_1482),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1513),
.B(n_1480),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1506),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1510),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1517),
.B(n_1507),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1535),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1529),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1556),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1562),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1574),
.B(n_1499),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1499),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1562),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1556),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

AND2x2_ASAP7_75t_SL g1607 ( 
.A(n_1583),
.B(n_1541),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1588),
.B(n_1511),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1557),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1557),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1585),
.B(n_1507),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1577),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1557),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1551),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1491),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1580),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1586),
.B(n_1484),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1577),
.B(n_1464),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1588),
.B(n_1469),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1484),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1589),
.B(n_1469),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1551),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1583),
.B(n_1484),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1580),
.Y(n_1625)
);

O2A1O1Ixp5_ASAP7_75t_L g1626 ( 
.A1(n_1589),
.A2(n_1500),
.B(n_1505),
.C(n_1502),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1559),
.B(n_1581),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1567),
.B(n_1564),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1559),
.A2(n_1502),
.B(n_1526),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1582),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_1596),
.B(n_1521),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1558),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1582),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1566),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1553),
.B(n_1533),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1583),
.B(n_1546),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1615),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1607),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1612),
.B(n_1637),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1613),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1615),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1623),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1623),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1617),
.B(n_1566),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1599),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1611),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1612),
.B(n_1637),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1597),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1617),
.B(n_1625),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1599),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1603),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1595),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1625),
.A2(n_1587),
.B(n_1596),
.C(n_1503),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1573),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1613),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1635),
.B(n_1573),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1600),
.B(n_1595),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1627),
.B(n_1553),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1606),
.Y(n_1661)
);

NAND4xp25_ASAP7_75t_L g1662 ( 
.A(n_1630),
.B(n_1587),
.C(n_1596),
.D(n_1503),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1600),
.B(n_1595),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1629),
.B(n_1582),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1629),
.B(n_1584),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1607),
.A2(n_1519),
.B(n_1501),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1607),
.A2(n_1578),
.B(n_1581),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1630),
.B(n_1584),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1627),
.B(n_1563),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1563),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1624),
.A2(n_1563),
.B(n_1568),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1600),
.B(n_1590),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1608),
.B(n_1592),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1606),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1632),
.A2(n_1628),
.B1(n_1636),
.B2(n_1624),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1636),
.B(n_1592),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1604),
.B(n_1590),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1620),
.B(n_1593),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1628),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1604),
.B(n_1590),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1664),
.B(n_1620),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1638),
.Y(n_1682)
);

AND3x1_ASAP7_75t_L g1683 ( 
.A(n_1666),
.B(n_1624),
.C(n_1611),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1638),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1647),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1647),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1642),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1669),
.B(n_1622),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1640),
.B(n_1648),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1655),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1645),
.B(n_1622),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1655),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1650),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1657),
.B(n_1619),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1641),
.B(n_1619),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1644),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1639),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1640),
.B(n_1648),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1654),
.A2(n_1628),
.B1(n_1636),
.B2(n_1560),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1653),
.B(n_1628),
.Y(n_1702)
);

NAND2x1_ASAP7_75t_L g1703 ( 
.A(n_1679),
.B(n_1628),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1641),
.B(n_1291),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1662),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1561),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1653),
.B(n_1604),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1669),
.B(n_1601),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1646),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1651),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1652),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1661),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1656),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1658),
.B(n_1649),
.Y(n_1714)
);

AOI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1675),
.A2(n_1558),
.B1(n_1571),
.B2(n_1578),
.C1(n_1601),
.C2(n_1602),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1668),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1699),
.B(n_1649),
.Y(n_1717)
);

OAI322xp33_ASAP7_75t_L g1718 ( 
.A1(n_1705),
.A2(n_1614),
.A3(n_1610),
.B1(n_1609),
.B2(n_1605),
.C1(n_1598),
.C2(n_1660),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1705),
.A2(n_1514),
.B1(n_1605),
.B2(n_1598),
.Y(n_1719)
);

XNOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1704),
.B(n_1572),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1684),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1690),
.B(n_1659),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1688),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1691),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1694),
.B(n_1294),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1713),
.B(n_1659),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1716),
.B(n_1690),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1670),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1683),
.A2(n_1626),
.B1(n_1558),
.B2(n_1571),
.C(n_1610),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1701),
.A2(n_1671),
.B1(n_1660),
.B2(n_1670),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_R g1733 ( 
.A(n_1700),
.B(n_1321),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1714),
.A2(n_1715),
.B(n_1706),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1681),
.A2(n_1605),
.B1(n_1609),
.B2(n_1598),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1681),
.A2(n_1610),
.B1(n_1614),
.B2(n_1609),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1693),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1700),
.A2(n_1575),
.B1(n_1558),
.B2(n_1571),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1693),
.Y(n_1739)
);

OAI32xp33_ASAP7_75t_L g1740 ( 
.A1(n_1708),
.A2(n_1679),
.A3(n_1611),
.B1(n_1614),
.B2(n_1602),
.Y(n_1740)
);

NAND4xp75_ASAP7_75t_L g1741 ( 
.A(n_1685),
.B(n_1626),
.C(n_1512),
.D(n_1672),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1682),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1722),
.B(n_1707),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1726),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1721),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1720),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1717),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1730),
.B(n_1708),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1723),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1707),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1728),
.B(n_1727),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1743),
.B(n_1572),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1734),
.B(n_1663),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1743),
.B(n_1689),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1742),
.B(n_1702),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1719),
.B(n_1663),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1732),
.B(n_1672),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1677),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1735),
.B(n_1677),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1736),
.B(n_1702),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1725),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1741),
.B(n_1338),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1731),
.A2(n_1703),
.B1(n_1611),
.B2(n_1689),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1745),
.B(n_1320),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1763),
.A2(n_1738),
.B(n_1740),
.C(n_1729),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_SL g1767 ( 
.A(n_1752),
.B(n_1718),
.C(n_1733),
.Y(n_1767)
);

OAI32xp33_ASAP7_75t_L g1768 ( 
.A1(n_1754),
.A2(n_1697),
.A3(n_1696),
.B1(n_1739),
.B2(n_1737),
.Y(n_1768)
);

O2A1O1Ixp5_ASAP7_75t_L g1769 ( 
.A1(n_1764),
.A2(n_1703),
.B(n_1685),
.C(n_1686),
.Y(n_1769)
);

NOR2x1_ASAP7_75t_L g1770 ( 
.A(n_1747),
.B(n_1325),
.Y(n_1770)
);

NOR4xp25_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1686),
.C(n_1698),
.D(n_1695),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1747),
.B(n_1679),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1753),
.A2(n_1712),
.B(n_1710),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1749),
.B(n_1673),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1746),
.B(n_1712),
.C(n_1711),
.Y(n_1775)
);

O2A1O1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1748),
.A2(n_1758),
.B(n_1759),
.C(n_1757),
.Y(n_1776)
);

NOR3x1_ASAP7_75t_L g1777 ( 
.A(n_1755),
.B(n_1709),
.C(n_1676),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1766),
.A2(n_1751),
.B(n_1760),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1770),
.B(n_1756),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1767),
.A2(n_1761),
.B1(n_1756),
.B2(n_1744),
.Y(n_1780)
);

NOR3x1_ASAP7_75t_L g1781 ( 
.A(n_1772),
.B(n_1762),
.C(n_1750),
.Y(n_1781)
);

AOI211x1_ASAP7_75t_L g1782 ( 
.A1(n_1768),
.A2(n_1674),
.B(n_1678),
.C(n_1680),
.Y(n_1782)
);

AND5x1_ASAP7_75t_L g1783 ( 
.A(n_1776),
.B(n_1575),
.C(n_1350),
.D(n_1325),
.E(n_1676),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1771),
.B(n_1769),
.C(n_1765),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_SL g1785 ( 
.A(n_1765),
.B(n_1298),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1765),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1774),
.B(n_1298),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1775),
.B(n_1338),
.Y(n_1788)
);

NAND4xp25_ASAP7_75t_L g1789 ( 
.A(n_1778),
.B(n_1777),
.C(n_1773),
.D(n_1680),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1785),
.B(n_1321),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1784),
.A2(n_1633),
.B(n_1571),
.C(n_1560),
.Y(n_1791)
);

AOI211x1_ASAP7_75t_SL g1792 ( 
.A1(n_1779),
.A2(n_1633),
.B(n_1518),
.C(n_1539),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_L g1793 ( 
.A(n_1786),
.B(n_1633),
.C(n_1350),
.Y(n_1793)
);

NOR3xp33_ASAP7_75t_L g1794 ( 
.A(n_1788),
.B(n_1631),
.C(n_1634),
.Y(n_1794)
);

AND4x1_ASAP7_75t_L g1795 ( 
.A(n_1781),
.B(n_1616),
.C(n_1555),
.D(n_1560),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1787),
.A2(n_1634),
.B(n_1631),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1795),
.B(n_1780),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1793),
.A2(n_1783),
.B1(n_1782),
.B2(n_1555),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1790),
.A2(n_1555),
.B1(n_1568),
.B2(n_1579),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1792),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1789),
.A2(n_1568),
.B1(n_1579),
.B2(n_1565),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1791),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1796),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1803),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1802),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1797),
.B(n_1794),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1800),
.Y(n_1807)
);

AO22x1_ASAP7_75t_L g1808 ( 
.A1(n_1798),
.A2(n_1616),
.B1(n_1621),
.B2(n_1618),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1801),
.B(n_1616),
.Y(n_1809)
);

AND2x2_ASAP7_75t_SL g1810 ( 
.A(n_1806),
.B(n_1799),
.Y(n_1810)
);

NAND2x1p5_ASAP7_75t_L g1811 ( 
.A(n_1804),
.B(n_1618),
.Y(n_1811)
);

NOR4xp25_ASAP7_75t_L g1812 ( 
.A(n_1805),
.B(n_1567),
.C(n_1565),
.D(n_1561),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1811),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1813),
.B(n_1807),
.C(n_1808),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1810),
.B1(n_1809),
.B2(n_1812),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1814),
.A2(n_1593),
.B1(n_1618),
.B2(n_1621),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1815),
.B(n_1561),
.Y(n_1817)
);

XNOR2xp5_ASAP7_75t_L g1818 ( 
.A(n_1816),
.B(n_1365),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1817),
.A2(n_1565),
.B(n_1569),
.Y(n_1819)
);

AO21x2_ASAP7_75t_L g1820 ( 
.A1(n_1818),
.A2(n_1621),
.B(n_1570),
.Y(n_1820)
);

OAI222xp33_ASAP7_75t_L g1821 ( 
.A1(n_1819),
.A2(n_1567),
.B1(n_1579),
.B2(n_1554),
.C1(n_1552),
.C2(n_1569),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1821),
.A2(n_1820),
.B1(n_1564),
.B2(n_1576),
.Y(n_1822)
);

OAI221xp5_ASAP7_75t_R g1823 ( 
.A1(n_1822),
.A2(n_1569),
.B1(n_1570),
.B2(n_1594),
.C(n_1591),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1554),
.B(n_1552),
.C(n_1564),
.Y(n_1824)
);


endmodule