module fake_jpeg_11569_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_72),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_6),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_54),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_7),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_70),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_61),
.B(n_68),
.Y(n_92)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_23),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_77),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_13),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_36),
.Y(n_107)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_26),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_41),
.B1(n_16),
.B2(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_90),
.B1(n_102),
.B2(n_119),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_20),
.B1(n_37),
.B2(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_82),
.A2(n_99),
.B1(n_118),
.B2(n_0),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_41),
.B1(n_16),
.B2(n_31),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_37),
.B1(n_23),
.B2(n_26),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_36),
.B1(n_39),
.B2(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_47),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_114),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_57),
.A2(n_59),
.B1(n_58),
.B2(n_43),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_75),
.B1(n_73),
.B2(n_56),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_38),
.Y(n_112)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_112),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_38),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_19),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_52),
.B(n_19),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_122),
.B(n_124),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_42),
.A2(n_40),
.B1(n_33),
.B2(n_15),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_45),
.A2(n_18),
.B1(n_28),
.B2(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_18),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_60),
.B(n_28),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_33),
.B1(n_40),
.B2(n_15),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g201 ( 
.A1(n_131),
.A2(n_153),
.B1(n_155),
.B2(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_51),
.B1(n_69),
.B2(n_22),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_139),
.B1(n_144),
.B2(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_148),
.Y(n_178)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_143),
.Y(n_170)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_84),
.A2(n_48),
.B(n_72),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_147),
.Y(n_199)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_118),
.B1(n_126),
.B2(n_84),
.Y(n_142)
);

AO21x2_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_169),
.B(n_80),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_56),
.B1(n_52),
.B2(n_72),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_97),
.B(n_111),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_1),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_160),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_9),
.B(n_11),
.C(n_4),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_80),
.B(n_105),
.C(n_106),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_9),
.B1(n_11),
.B2(n_4),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_152),
.A2(n_133),
.B1(n_130),
.B2(n_168),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_94),
.Y(n_177)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_85),
.A2(n_5),
.B(n_106),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_88),
.B(n_120),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_87),
.B(n_123),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_88),
.B1(n_120),
.B2(n_113),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_96),
.A2(n_101),
.B1(n_123),
.B2(n_98),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_105),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_199),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_197),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_190),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_135),
.B(n_158),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_101),
.B1(n_98),
.B2(n_125),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_184),
.B1(n_194),
.B2(n_201),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_129),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_188),
.B(n_191),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_94),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_103),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_192),
.B(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_125),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_154),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_139),
.B(n_151),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_137),
.B1(n_140),
.B2(n_159),
.Y(n_211)
);

INVx5_ASAP7_75t_SL g196 ( 
.A(n_138),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

OR2x2_ASAP7_75t_SL g197 ( 
.A(n_128),
.B(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_132),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_162),
.B1(n_163),
.B2(n_161),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_208),
.C(n_217),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_205),
.A2(n_213),
.B1(n_171),
.B2(n_175),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_129),
.C(n_160),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_225),
.B(n_227),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_178),
.B(n_150),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_218),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_172),
.B(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_195),
.B1(n_184),
.B2(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_191),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_193),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_180),
.C(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_228),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_201),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_184),
.B1(n_203),
.B2(n_183),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_184),
.B1(n_174),
.B2(n_176),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_250),
.B1(n_216),
.B2(n_209),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_179),
.Y(n_239)
);

OAI322xp33_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_241),
.A3(n_245),
.B1(n_234),
.B2(n_237),
.C1(n_231),
.C2(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_189),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_187),
.B1(n_198),
.B2(n_181),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_222),
.B1(n_211),
.B2(n_221),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_181),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_223),
.B1(n_228),
.B2(n_227),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_247),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_171),
.A3(n_175),
.B1(n_198),
.B2(n_210),
.C1(n_217),
.C2(n_214),
.Y(n_248)
);

AOI221xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_237),
.B1(n_245),
.B2(n_241),
.C(n_239),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_229),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_257),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_235),
.B1(n_238),
.B2(n_233),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_255),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_208),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_212),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_215),
.B1(n_220),
.B2(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_234),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_260),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_242),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_264),
.Y(n_268)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_232),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_247),
.B1(n_236),
.B2(n_230),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_279),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_254),
.B1(n_262),
.B2(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_282),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_271),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_287),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_255),
.C(n_249),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_249),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_278),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_269),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_262),
.B(n_270),
.Y(n_291)
);

AO21x1_ASAP7_75t_SL g302 ( 
.A1(n_291),
.A2(n_273),
.B(n_246),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_275),
.B1(n_277),
.B2(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_295),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_275),
.B1(n_258),
.B2(n_279),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_276),
.B(n_256),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_273),
.B(n_266),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_248),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_301),
.B(n_302),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_260),
.C(n_246),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_296),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_294),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_290),
.C(n_300),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_306),
.A2(n_304),
.B(n_291),
.Y(n_308)
);

OAI311xp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_307),
.A3(n_295),
.B1(n_263),
.C1(n_240),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_240),
.C(n_263),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_243),
.Y(n_311)
);


endmodule