module fake_jpeg_2769_n_234 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_234);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_19),
.B(n_2),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_89),
.Y(n_97)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_56),
.B1(n_74),
.B2(n_67),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_80),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_61),
.B1(n_73),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_82),
.B1(n_87),
.B2(n_85),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_61),
.B1(n_74),
.B2(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_63),
.B1(n_79),
.B2(n_75),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_86),
.B1(n_87),
.B2(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_109),
.B1(n_120),
.B2(n_24),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_118),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_86),
.B1(n_88),
.B2(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_66),
.C(n_68),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_116),
.C(n_54),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_88),
.B1(n_63),
.B2(n_79),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_115),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_60),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_122),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_73),
.B1(n_54),
.B2(n_58),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_59),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_54),
.B(n_64),
.C(n_73),
.Y(n_123)
);

AO21x2_ASAP7_75t_SL g130 ( 
.A1(n_123),
.A2(n_94),
.B(n_64),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_3),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_57),
.A3(n_62),
.B1(n_70),
.B2(n_71),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_130),
.A3(n_135),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_46),
.B(n_45),
.C(n_41),
.Y(n_168)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_0),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_1),
.Y(n_138)
);

NAND2x1_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_102),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_139),
.A2(n_144),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_1),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_143),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_8),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_2),
.Y(n_143)
);

NAND2x1_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_3),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_162),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_26),
.B1(n_52),
.B2(n_51),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_156),
.B1(n_168),
.B2(n_32),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_126),
.B(n_132),
.C(n_139),
.D(n_144),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_170),
.B(n_34),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_4),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_171),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_166),
.Y(n_188)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_10),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_9),
.B(n_10),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_9),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_40),
.C(n_39),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_173),
.C(n_156),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_37),
.C(n_35),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_180),
.B(n_185),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_11),
.B(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_13),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_183),
.B(n_190),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_30),
.B(n_14),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_187),
.B(n_170),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_13),
.B(n_14),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_15),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_154),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_172),
.C(n_182),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_205),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_174),
.B1(n_189),
.B2(n_181),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_152),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_208),
.C(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_176),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_177),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_189),
.B1(n_169),
.B2(n_187),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_212),
.B1(n_195),
.B2(n_210),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_188),
.B(n_184),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_213),
.B(n_199),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_179),
.B(n_155),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_211),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_222),
.C(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_218),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

OAI31xp33_ASAP7_75t_SL g230 ( 
.A1(n_229),
.A2(n_225),
.A3(n_223),
.B(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_226),
.C(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_177),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_194),
.Y(n_234)
);


endmodule