module fake_jpeg_2519_n_227 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_7),
.B(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx6f_ASAP7_75t_SL g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_54),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_78),
.C(n_57),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_72),
.B1(n_73),
.B2(n_54),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_96),
.B1(n_100),
.B2(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_73),
.B1(n_54),
.B2(n_66),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_66),
.B1(n_60),
.B2(n_63),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_115),
.Y(n_138)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

OR2x4_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_82),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_75),
.B(n_43),
.C(n_39),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_117),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

CKINVDCx6p67_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_88),
.B(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_121),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_79),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_65),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_67),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_60),
.B1(n_64),
.B2(n_76),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_100),
.B1(n_79),
.B2(n_61),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_132),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_56),
.B(n_76),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_128),
.B(n_5),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_61),
.A3(n_56),
.B1(n_74),
.B2(n_69),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_59),
.B1(n_58),
.B2(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_51),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_50),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_0),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_22),
.Y(n_159)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_108),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_149),
.Y(n_175)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_168),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_3),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_122),
.B1(n_132),
.B2(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_159),
.Y(n_177)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_48),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_45),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_164),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_38),
.B(n_37),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_25),
.B(n_6),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_4),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_165),
.B(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_4),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_180),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_182),
.B1(n_186),
.B2(n_179),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_5),
.B(n_6),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_161),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_194),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_156),
.A3(n_158),
.B1(n_160),
.B2(n_168),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_201),
.B1(n_169),
.B2(n_182),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_151),
.B1(n_161),
.B2(n_13),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_184),
.B(n_176),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_177),
.B(n_180),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_173),
.B1(n_192),
.B2(n_188),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_183),
.C(n_170),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_210),
.C(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_173),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_214),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_216),
.C(n_210),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_203),
.B1(n_209),
.B2(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_215),
.Y(n_221)
);

XOR2x1_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_217),
.B1(n_220),
.B2(n_18),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_222),
.B(n_17),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_224),
.B(n_15),
.Y(n_225)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_19),
.B(n_20),
.Y(n_227)
);


endmodule