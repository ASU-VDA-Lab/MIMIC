module fake_ariane_2239_n_1323 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1323);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1323;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1257;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_671;
wire n_1148;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_59),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_111),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_45),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_68),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_16),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_54),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_45),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_56),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_174),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_53),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_150),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_89),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_75),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_101),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_1),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_73),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_98),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_116),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_79),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_145),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_76),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_22),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_104),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_29),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_176),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_106),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_69),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_90),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_64),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_40),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_91),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_107),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_122),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_12),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_20),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_170),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_81),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_62),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_105),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_100),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_99),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_191),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_17),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_43),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_47),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_181),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_128),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_14),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_165),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_30),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_86),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_82),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_6),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_72),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_51),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_157),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_42),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_96),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_11),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_60),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_29),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_151),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_26),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_66),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_24),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_36),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_169),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_125),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_186),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_94),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_11),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_158),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_80),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_67),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_173),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_161),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_171),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_31),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_137),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_39),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_202),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_193),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_R g317 ( 
.A(n_203),
.B(n_49),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_214),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_202),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_204),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_225),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_205),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_194),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_251),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_194),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_195),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_251),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_196),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_234),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_197),
.B(n_0),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_215),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_229),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

BUFx6f_ASAP7_75t_SL g339 ( 
.A(n_210),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_246),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_226),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_208),
.B(n_228),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_258),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_226),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_308),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_230),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_217),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_210),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_238),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_251),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_R g353 ( 
.A(n_207),
.B(n_50),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_226),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_195),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_197),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_267),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_198),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_198),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_200),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_226),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_226),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_199),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_267),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_294),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_199),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_200),
.B(n_0),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_201),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_201),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_206),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_216),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_294),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_294),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_262),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_262),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_220),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_224),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_206),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_218),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_310),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_310),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_312),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_218),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_253),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_242),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_244),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_247),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_248),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_239),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_231),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_233),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_250),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_264),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_270),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_282),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_253),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_289),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_311),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_335),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_325),
.B(n_213),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_325),
.B(n_213),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_328),
.B(n_239),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_354),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_354),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_328),
.B(n_329),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_209),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_336),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_349),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_315),
.B(n_311),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_347),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_316),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_359),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_296),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_319),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_340),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_343),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_329),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_356),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_356),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_320),
.B(n_252),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_321),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_402),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_384),
.B(n_255),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_400),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_291),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_401),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_342),
.B(n_306),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_322),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_323),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_333),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_337),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_338),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

BUFx8_ASAP7_75t_L g460 ( 
.A(n_339),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_360),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_345),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_360),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_357),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_362),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_339),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_339),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_369),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_334),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_361),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_443),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_452),
.B(n_321),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_296),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_451),
.A2(n_326),
.B1(n_318),
.B2(n_358),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_414),
.Y(n_485)
);

AND2x6_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_307),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_409),
.B(n_361),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_429),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_412),
.B(n_367),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_467),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_416),
.B(n_371),
.C(n_367),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_410),
.B(n_371),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_413),
.B(n_373),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_467),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_454),
.B(n_331),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_411),
.A2(n_324),
.B1(n_375),
.B2(n_358),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_413),
.B(n_373),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_451),
.B(n_317),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_404),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_460),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_426),
.A2(n_375),
.B1(n_324),
.B2(n_404),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_425),
.B(n_307),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_415),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_435),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_454),
.B(n_332),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

INVxp33_ASAP7_75t_SL g512 ( 
.A(n_438),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_471),
.B(n_374),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_374),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_217),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_418),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_470),
.B(n_379),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_470),
.B(n_379),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_445),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_380),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_456),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_472),
.B(n_380),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_433),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_425),
.B(n_364),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_443),
.B(n_385),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_454),
.B(n_389),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_472),
.B(n_372),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_443),
.B(n_385),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g536 ( 
.A(n_426),
.B(n_217),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_469),
.B(n_217),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_445),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_460),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_446),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_472),
.B(n_386),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_456),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_443),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_466),
.B(n_327),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_485),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_527),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_527),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_536),
.A2(n_453),
.B1(n_444),
.B2(n_426),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_536),
.B(n_426),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_446),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_439),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_485),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_519),
.B(n_439),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_540),
.B(n_440),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_473),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_522),
.B(n_422),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_513),
.B(n_422),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_515),
.B(n_440),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_524),
.B(n_466),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g562 ( 
.A(n_501),
.B(n_494),
.C(n_492),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_476),
.B(n_474),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_502),
.B(n_466),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g565 ( 
.A(n_501),
.B(n_387),
.C(n_386),
.Y(n_565)
);

OA22x2_ASAP7_75t_L g566 ( 
.A1(n_499),
.A2(n_474),
.B1(n_455),
.B2(n_459),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_496),
.B(n_449),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_502),
.B(n_466),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_483),
.B(n_440),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g570 ( 
.A1(n_487),
.A2(n_393),
.B(n_387),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_500),
.B(n_449),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_545),
.B(n_393),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_545),
.B(n_460),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_490),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_520),
.B(n_542),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_495),
.B(n_440),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_507),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_489),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_498),
.B(n_381),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_498),
.B(n_382),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_510),
.B(n_512),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_503),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_510),
.B(n_460),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_484),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_512),
.B(n_509),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_531),
.B(n_442),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_544),
.A2(n_417),
.B(n_442),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_509),
.B(n_396),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_531),
.B(n_447),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_506),
.B(n_447),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_509),
.B(n_397),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_526),
.B(n_448),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_503),
.B(n_448),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_531),
.B(n_450),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_489),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_L g600 ( 
.A(n_517),
.B(n_465),
.C(n_458),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_532),
.B(n_450),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_531),
.A2(n_417),
.B1(n_453),
.B2(n_444),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_535),
.B(n_456),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_475),
.B(n_456),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_508),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_480),
.B(n_456),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_481),
.Y(n_608)
);

AOI221xp5_ASAP7_75t_L g609 ( 
.A1(n_505),
.A2(n_330),
.B1(n_368),
.B2(n_459),
.C(n_458),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_482),
.B(n_457),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_493),
.B(n_457),
.Y(n_611)
);

O2A1O1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_529),
.A2(n_465),
.B(n_464),
.C(n_455),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_529),
.A2(n_533),
.B1(n_479),
.B2(n_486),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_533),
.B(n_457),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_511),
.B(n_457),
.Y(n_615)
);

AOI221xp5_ASAP7_75t_L g616 ( 
.A1(n_478),
.A2(n_464),
.B1(n_287),
.B2(n_280),
.C(n_295),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_497),
.B(n_457),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_518),
.B(n_405),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_491),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_479),
.B(n_457),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_518),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_521),
.B(n_405),
.Y(n_623)
);

NAND2x1_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_420),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_511),
.B(n_444),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_507),
.A2(n_453),
.B1(n_407),
.B2(n_406),
.Y(n_626)
);

BUFx8_ASAP7_75t_L g627 ( 
.A(n_539),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_491),
.B(n_350),
.Y(n_628)
);

BUFx5_ASAP7_75t_L g629 ( 
.A(n_479),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_491),
.B(n_477),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_511),
.B(n_514),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_479),
.B(n_419),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_479),
.B(n_419),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_479),
.B(n_428),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_484),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_486),
.B(n_428),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_486),
.B(n_314),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_486),
.B(n_406),
.Y(n_638)
);

AND2x4_ASAP7_75t_SL g639 ( 
.A(n_514),
.B(n_541),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_484),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_523),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_514),
.B(n_353),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_486),
.B(n_407),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_523),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_486),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_547),
.Y(n_646)
);

NOR2x1p5_ASAP7_75t_SL g647 ( 
.A(n_629),
.B(n_434),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_567),
.B(n_528),
.Y(n_648)
);

AO21x1_ASAP7_75t_L g649 ( 
.A1(n_614),
.A2(n_488),
.B(n_477),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_622),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_623),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_561),
.A2(n_534),
.B(n_488),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_571),
.B(n_541),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_630),
.A2(n_534),
.B(n_488),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_572),
.A2(n_538),
.B(n_420),
.C(n_415),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_618),
.B(n_541),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_539),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_576),
.A2(n_265),
.B(n_263),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_585),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_586),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_552),
.A2(n_420),
.B(n_429),
.C(n_434),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_576),
.B(n_427),
.C(n_424),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_585),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_574),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_562),
.B(n_523),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_630),
.A2(n_534),
.B(n_523),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_546),
.B(n_431),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_571),
.B(n_352),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_558),
.A2(n_420),
.B(n_434),
.C(n_436),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_594),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_575),
.A2(n_543),
.B(n_436),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_575),
.A2(n_537),
.B(n_516),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_564),
.A2(n_543),
.B(n_436),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_582),
.B(n_432),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_627),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_608),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_557),
.B(n_348),
.C(n_543),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_559),
.B(n_543),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_568),
.A2(n_212),
.B(n_211),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_562),
.B(n_217),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_603),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_644),
.A2(n_260),
.B(n_221),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_614),
.A2(n_537),
.B(n_516),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_589),
.A2(n_644),
.B(n_555),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_557),
.B(n_273),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_624),
.A2(n_222),
.B(n_219),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_553),
.A2(n_278),
.B(n_292),
.C(n_302),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_563),
.A2(n_537),
.B(n_516),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g690 ( 
.A1(n_559),
.A2(n_537),
.B(n_516),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_577),
.B(n_2),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_563),
.B(n_516),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_588),
.B(n_516),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_621),
.A2(n_537),
.B(n_260),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_600),
.A2(n_537),
.B1(n_269),
.B2(n_309),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_579),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_569),
.B(n_580),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_596),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_578),
.A2(n_227),
.B(n_223),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_578),
.A2(n_605),
.B(n_599),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_599),
.A2(n_235),
.B(n_232),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_605),
.A2(n_272),
.B(n_304),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_548),
.B(n_3),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_620),
.A2(n_268),
.B(n_303),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_606),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_620),
.A2(n_261),
.B(n_301),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_549),
.B(n_4),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_551),
.A2(n_236),
.B1(n_299),
.B2(n_298),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_588),
.B(n_237),
.Y(n_710)
);

AOI21x1_ASAP7_75t_L g711 ( 
.A1(n_632),
.A2(n_421),
.B(n_260),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_612),
.A2(n_260),
.B(n_297),
.C(n_293),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_591),
.B(n_240),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_595),
.A2(n_241),
.B(n_288),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_601),
.A2(n_245),
.B(n_286),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_635),
.A2(n_249),
.B(n_283),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_629),
.B(n_260),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_640),
.A2(n_259),
.B(n_281),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_641),
.A2(n_279),
.B(n_276),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_591),
.A2(n_598),
.B(n_570),
.C(n_600),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_604),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_628),
.B(n_639),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_615),
.A2(n_610),
.B(n_607),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_581),
.B(n_254),
.C(n_256),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_598),
.A2(n_257),
.B(n_421),
.C(n_7),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_560),
.A2(n_4),
.B(n_5),
.C(n_8),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_611),
.A2(n_421),
.B(n_88),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_628),
.B(n_5),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_617),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_625),
.A2(n_421),
.B(n_92),
.Y(n_731)
);

AOI21x1_ASAP7_75t_L g732 ( 
.A1(n_633),
.A2(n_421),
.B(n_87),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_626),
.B(n_9),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_556),
.A2(n_421),
.B(n_93),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_626),
.B(n_9),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_590),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_573),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_585),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_634),
.A2(n_636),
.B(n_585),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_638),
.A2(n_102),
.B(n_190),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_619),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_584),
.B(n_19),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_550),
.B(n_597),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_657),
.B(n_583),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_709),
.B(n_550),
.Y(n_745)
);

NAND2x1_ASAP7_75t_L g746 ( 
.A(n_659),
.B(n_583),
.Y(n_746)
);

NAND2x1_ASAP7_75t_L g747 ( 
.A(n_659),
.B(n_613),
.Y(n_747)
);

AND3x1_ASAP7_75t_L g748 ( 
.A(n_668),
.B(n_616),
.C(n_609),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_650),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_645),
.A2(n_565),
.B(n_619),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_676),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_SL g752 ( 
.A(n_669),
.B(n_587),
.C(n_593),
.Y(n_752)
);

AOI21xp33_ASAP7_75t_L g753 ( 
.A1(n_733),
.A2(n_566),
.B(n_602),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_681),
.A2(n_643),
.B(n_566),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_711),
.A2(n_637),
.B(n_631),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_685),
.A2(n_619),
.B(n_642),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_651),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_694),
.A2(n_629),
.B(n_619),
.Y(n_758)
);

INVx5_ASAP7_75t_L g759 ( 
.A(n_664),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_686),
.A2(n_629),
.B(n_627),
.C(n_21),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_651),
.B(n_52),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_648),
.B(n_629),
.Y(n_762)
);

OAI21xp33_ASAP7_75t_SL g763 ( 
.A1(n_653),
.A2(n_629),
.B(n_20),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_681),
.A2(n_19),
.B(n_21),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_743),
.B(n_22),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_664),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_664),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_660),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_SL g769 ( 
.A1(n_686),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C(n_27),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_739),
.A2(n_110),
.B(n_189),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_719),
.B(n_23),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_679),
.A2(n_25),
.B(n_28),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_664),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_652),
.A2(n_113),
.B(n_188),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_721),
.A2(n_658),
.B(n_729),
.C(n_697),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_732),
.A2(n_112),
.B(n_184),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_660),
.Y(n_777)
);

NOR2x1_ASAP7_75t_SL g778 ( 
.A(n_741),
.B(n_55),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_666),
.A2(n_30),
.B(n_31),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_656),
.B(n_32),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_724),
.A2(n_114),
.B(n_179),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_666),
.A2(n_32),
.B(n_33),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_654),
.A2(n_33),
.B(n_34),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_667),
.A2(n_115),
.B(n_172),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_674),
.A2(n_109),
.B(n_168),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_705),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_705),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_657),
.B(n_34),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_697),
.B(n_35),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_719),
.B(n_35),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_723),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_675),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_703),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_682),
.B(n_37),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_675),
.B(n_38),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_672),
.A2(n_121),
.B(n_167),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_738),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_692),
.A2(n_119),
.B(n_164),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_717),
.A2(n_118),
.B(n_163),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_721),
.B(n_41),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_722),
.B(n_41),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_691),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_802)
);

AOI221xp5_ASAP7_75t_SL g803 ( 
.A1(n_688),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_663),
.B(n_48),
.C(n_57),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_707),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_SL g806 ( 
.A(n_725),
.B(n_58),
.C(n_61),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_691),
.B(n_63),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_730),
.B(n_661),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_671),
.B(n_65),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_717),
.A2(n_70),
.B(n_71),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_700),
.A2(n_74),
.B(n_77),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_677),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_662),
.A2(n_78),
.B(n_83),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_728),
.A2(n_84),
.B(n_85),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_696),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_678),
.Y(n_816)
);

BUFx2_ASAP7_75t_SL g817 ( 
.A(n_749),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_744),
.B(n_647),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_757),
.B(n_710),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_744),
.B(n_759),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_762),
.A2(n_673),
.B(n_689),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_790),
.B(n_725),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_789),
.B(n_713),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_815),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_779),
.A2(n_737),
.B(n_726),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_808),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_748),
.A2(n_735),
.B1(n_742),
.B2(n_726),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_808),
.B(n_708),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_790),
.B(n_737),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_751),
.B(n_736),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_780),
.B(n_791),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_809),
.B(n_693),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_771),
.Y(n_833)
);

CKINVDCx11_ASAP7_75t_R g834 ( 
.A(n_788),
.Y(n_834)
);

NOR2x1_ASAP7_75t_SL g835 ( 
.A(n_759),
.B(n_646),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_768),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_762),
.A2(n_670),
.B(n_649),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_795),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_759),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_SL g841 ( 
.A(n_744),
.B(n_727),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_759),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_809),
.B(n_665),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_756),
.A2(n_684),
.B(n_734),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_745),
.B(n_698),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_800),
.A2(n_695),
.B1(n_690),
.B2(n_740),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_781),
.A2(n_731),
.B(n_655),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_771),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_786),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_805),
.B(n_712),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_816),
.B(n_745),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_793),
.B(n_715),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_787),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_788),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_775),
.A2(n_712),
.B(n_680),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_812),
.B(n_714),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_747),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_788),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_754),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_805),
.B(n_720),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_797),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_805),
.B(n_716),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_794),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_800),
.B(n_701),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_797),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_805),
.B(n_718),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_766),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_813),
.A2(n_706),
.B(n_704),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_752),
.B(n_702),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_797),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_794),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_801),
.B(n_699),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_801),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_766),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_792),
.B(n_683),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_807),
.A2(n_687),
.B1(n_97),
.B2(n_108),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_750),
.A2(n_95),
.B(n_123),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_765),
.B(n_129),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_765),
.B(n_130),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_767),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_772),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_772),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_761),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_779),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_824),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_836),
.Y(n_886)
);

INVx6_ASAP7_75t_L g887 ( 
.A(n_820),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_829),
.A2(n_823),
.B1(n_827),
.B2(n_839),
.Y(n_888)
);

AO21x2_ASAP7_75t_L g889 ( 
.A1(n_838),
.A2(n_753),
.B(n_813),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_854),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_820),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_861),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_831),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_837),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_837),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_878),
.A2(n_764),
.B(n_782),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_874),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_825),
.A2(n_760),
.B1(n_802),
.B2(n_782),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_853),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_853),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_874),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_859),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_822),
.A2(n_804),
.B1(n_764),
.B2(n_769),
.Y(n_904)
);

AO21x1_ASAP7_75t_L g905 ( 
.A1(n_878),
.A2(n_783),
.B(n_753),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_833),
.B(n_803),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_848),
.B(n_773),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_826),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_820),
.B(n_767),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_851),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_817),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_819),
.A2(n_783),
.B1(n_746),
.B2(n_773),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_861),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_865),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_863),
.B(n_871),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_881),
.A2(n_814),
.B(n_755),
.Y(n_916)
);

INVx4_ASAP7_75t_SL g917 ( 
.A(n_818),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_834),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_873),
.B(n_763),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_845),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_845),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_840),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_SL g923 ( 
.A1(n_875),
.A2(n_778),
.B1(n_811),
.B2(n_770),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_884),
.A2(n_774),
.B1(n_811),
.B2(n_798),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_855),
.A2(n_784),
.B(n_776),
.Y(n_925)
);

AOI21xp33_ASAP7_75t_L g926 ( 
.A1(n_872),
.A2(n_796),
.B(n_785),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_865),
.Y(n_927)
);

OAI22xp33_ASAP7_75t_L g928 ( 
.A1(n_854),
.A2(n_806),
.B1(n_810),
.B2(n_799),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_882),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_828),
.B(n_758),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_870),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_842),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_858),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_870),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_867),
.Y(n_935)
);

OAI22xp33_ASAP7_75t_L g936 ( 
.A1(n_858),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_936)
);

INVx8_ASAP7_75t_L g937 ( 
.A(n_843),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_867),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_834),
.A2(n_140),
.B1(n_141),
.B2(n_144),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_864),
.A2(n_844),
.B(n_821),
.Y(n_940)
);

BUFx2_ASAP7_75t_R g941 ( 
.A(n_842),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_867),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_874),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_858),
.B(n_146),
.Y(n_944)
);

CKINVDCx6p67_ASAP7_75t_R g945 ( 
.A(n_874),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_859),
.Y(n_946)
);

CKINVDCx6p67_ASAP7_75t_R g947 ( 
.A(n_874),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_880),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_857),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_857),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_880),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_857),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_840),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_843),
.A2(n_147),
.B1(n_148),
.B2(n_153),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_818),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_840),
.B(n_155),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_818),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_908),
.B(n_850),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_929),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_905),
.A2(n_864),
.B(n_847),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_946),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_903),
.Y(n_962)
);

NOR2x1_ASAP7_75t_L g963 ( 
.A(n_930),
.B(n_869),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_924),
.A2(n_847),
.B(n_868),
.Y(n_964)
);

NOR2x1_ASAP7_75t_R g965 ( 
.A(n_911),
.B(n_850),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_925),
.A2(n_850),
.B(n_877),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_920),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_921),
.B(n_879),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_916),
.A2(n_846),
.B(n_883),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_895),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_885),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_897),
.A2(n_869),
.B(n_846),
.Y(n_972)
);

AO21x2_ASAP7_75t_L g973 ( 
.A1(n_926),
.A2(n_856),
.B(n_852),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_899),
.A2(n_843),
.B1(n_832),
.B2(n_830),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_955),
.B(n_832),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_940),
.B(n_832),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_896),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_900),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_901),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_917),
.B(n_866),
.Y(n_980)
);

OA21x2_ASAP7_75t_L g981 ( 
.A1(n_919),
.A2(n_876),
.B(n_866),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_915),
.B(n_832),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_949),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_940),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_915),
.B(n_957),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_949),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_955),
.B(n_866),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_950),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_950),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_888),
.B(n_841),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_952),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_952),
.A2(n_862),
.B(n_860),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_886),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_945),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_916),
.A2(n_860),
.B(n_862),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_893),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_916),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_957),
.B(n_894),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_917),
.B(n_860),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_898),
.B(n_862),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_931),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_934),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_889),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_907),
.B(n_835),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_963),
.B(n_976),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_959),
.B(n_889),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_960),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_959),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_988),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_983),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_988),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_960),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_995),
.B(n_917),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_989),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_963),
.Y(n_1016)
);

OA222x2_ASAP7_75t_L g1017 ( 
.A1(n_998),
.A2(n_910),
.B1(n_938),
.B2(n_935),
.C1(n_942),
.C2(n_951),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_989),
.Y(n_1018)
);

AOI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_972),
.A2(n_906),
.B1(n_904),
.B2(n_936),
.C(n_933),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_972),
.B(n_948),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_976),
.B(n_984),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_995),
.B(n_902),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_976),
.B(n_923),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_984),
.B(n_890),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_984),
.B(n_945),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_997),
.B(n_947),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_983),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_997),
.B(n_960),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_990),
.A2(n_939),
.B1(n_936),
.B2(n_933),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_1003),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_986),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_986),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_980),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_971),
.B(n_918),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_989),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_973),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_962),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_980),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_991),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_960),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_960),
.B(n_947),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_962),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_971),
.B(n_914),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_985),
.B(n_943),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_962),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_967),
.B(n_902),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_991),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_961),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_985),
.B(n_943),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1003),
.B(n_898),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_967),
.B(n_912),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1016),
.B(n_973),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_L g1053 ( 
.A(n_1019),
.B(n_974),
.C(n_939),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1023),
.B(n_995),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1020),
.B(n_993),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_1033),
.B(n_911),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_SL g1057 ( 
.A1(n_1019),
.A2(n_954),
.B(n_944),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_L g1058 ( 
.A(n_1029),
.B(n_968),
.C(n_993),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1023),
.B(n_982),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1029),
.B(n_968),
.C(n_996),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1023),
.B(n_982),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1047),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1005),
.A2(n_981),
.B1(n_958),
.B2(n_1004),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1016),
.B(n_973),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1044),
.B(n_973),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1044),
.B(n_1004),
.Y(n_1066)
);

OAI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_1028),
.A2(n_954),
.B(n_958),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1044),
.B(n_992),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1005),
.A2(n_981),
.B1(n_937),
.B2(n_987),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1049),
.B(n_992),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1049),
.B(n_992),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1049),
.B(n_992),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_1036),
.A2(n_1040),
.B(n_1028),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1020),
.B(n_928),
.C(n_969),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1005),
.B(n_1033),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1006),
.B(n_996),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_SL g1077 ( 
.A(n_1051),
.B(n_928),
.C(n_1001),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_SL g1078 ( 
.A1(n_1028),
.A2(n_969),
.B(n_922),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_L g1079 ( 
.A(n_1040),
.B(n_981),
.C(n_1002),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1034),
.B(n_998),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_1014),
.B(n_965),
.Y(n_1081)
);

OAI221xp5_ASAP7_75t_L g1082 ( 
.A1(n_1034),
.A2(n_1002),
.B1(n_1001),
.B2(n_981),
.C(n_961),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1062),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1075),
.B(n_1033),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1076),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1075),
.B(n_1033),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_1080),
.B(n_1034),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1054),
.B(n_1038),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1054),
.B(n_1038),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1055),
.B(n_1051),
.Y(n_1090)
);

NAND4xp25_ASAP7_75t_L g1091 ( 
.A(n_1053),
.B(n_1028),
.C(n_1040),
.D(n_1046),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1076),
.B(n_1006),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1073),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1068),
.B(n_1038),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1065),
.B(n_1068),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1070),
.B(n_1071),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1065),
.B(n_1024),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1062),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1073),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1070),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1071),
.B(n_1006),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1072),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1073),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1072),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1073),
.B(n_1030),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1088),
.B(n_1066),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1088),
.B(n_1066),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1087),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1087),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_SL g1111 ( 
.A(n_1105),
.B(n_1038),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1090),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1085),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1091),
.B(n_1059),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_1105),
.B(n_1014),
.Y(n_1115)
);

NAND2x1_ASAP7_75t_L g1116 ( 
.A(n_1089),
.B(n_1094),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1093),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1106),
.B(n_1061),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1083),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1083),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_1116),
.B(n_1014),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1111),
.B(n_1093),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1109),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1117),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1117),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1116),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1110),
.B(n_1092),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1111),
.B(n_1107),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1123),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1128),
.B(n_1107),
.Y(n_1130)
);

INVx6_ASAP7_75t_L g1131 ( 
.A(n_1127),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1128),
.B(n_1108),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1121),
.B(n_1108),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1131),
.Y(n_1134)
);

AOI21xp33_ASAP7_75t_SL g1135 ( 
.A1(n_1130),
.A2(n_1126),
.B(n_1121),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1130),
.B(n_1121),
.Y(n_1136)
);

AOI33xp33_ASAP7_75t_L g1137 ( 
.A1(n_1131),
.A2(n_1126),
.A3(n_1113),
.B1(n_1122),
.B2(n_1103),
.B3(n_1099),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1131),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1129),
.Y(n_1139)
);

NAND4xp25_ASAP7_75t_L g1140 ( 
.A(n_1129),
.B(n_1114),
.C(n_1122),
.D(n_1053),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1132),
.Y(n_1141)
);

AND4x1_ASAP7_75t_L g1142 ( 
.A(n_1133),
.B(n_1081),
.C(n_1077),
.D(n_1060),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1131),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1129),
.A2(n_1125),
.B(n_1124),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1129),
.A2(n_1099),
.B1(n_1103),
.B2(n_1122),
.C(n_1124),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1134),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1138),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_1136),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1143),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1136),
.B(n_1118),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1141),
.B(n_1127),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1139),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1144),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1137),
.B(n_1115),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1140),
.B(n_1112),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1137),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1145),
.Y(n_1157)
);

AOI222xp33_ASAP7_75t_L g1158 ( 
.A1(n_1142),
.A2(n_1125),
.B1(n_1060),
.B2(n_1058),
.C1(n_1079),
.C2(n_1057),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1135),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1134),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1134),
.B(n_1095),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1134),
.B(n_1096),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1148),
.B(n_1096),
.Y(n_1163)
);

NOR4xp25_ASAP7_75t_SL g1164 ( 
.A(n_1157),
.B(n_1057),
.C(n_1120),
.D(n_1119),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1153),
.B(n_1064),
.C(n_1052),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1156),
.A2(n_1115),
.B(n_1064),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1151),
.B(n_1095),
.Y(n_1167)
);

OAI211xp5_ASAP7_75t_L g1168 ( 
.A1(n_1148),
.A2(n_1056),
.B(n_1078),
.C(n_1058),
.Y(n_1168)
);

AOI211xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1147),
.A2(n_1082),
.B(n_1081),
.C(n_1074),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1155),
.A2(n_1115),
.B(n_1052),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1155),
.A2(n_1104),
.B1(n_1102),
.B2(n_1100),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1151),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1146),
.B(n_1100),
.Y(n_1173)
);

OAI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1158),
.A2(n_1079),
.B1(n_1067),
.B2(n_1078),
.C(n_1036),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1154),
.A2(n_1067),
.B(n_1101),
.Y(n_1175)
);

AOI211xp5_ASAP7_75t_L g1176 ( 
.A1(n_1154),
.A2(n_1102),
.B(n_1104),
.C(n_1101),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1146),
.B(n_1092),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_1149),
.B(n_944),
.C(n_965),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1159),
.A2(n_1098),
.B(n_1013),
.C(n_1007),
.Y(n_1179)
);

AOI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1160),
.A2(n_1007),
.B1(n_1013),
.B2(n_1063),
.C(n_1097),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1148),
.A2(n_1098),
.B(n_1089),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1172),
.B(n_1148),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1177),
.B(n_1152),
.C(n_1161),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_SL g1184 ( 
.A(n_1164),
.B(n_1150),
.C(n_1162),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1163),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1169),
.B(n_1150),
.C(n_1030),
.Y(n_1186)
);

NOR2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1167),
.B(n_1094),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1173),
.Y(n_1188)
);

NOR3x1_ASAP7_75t_L g1189 ( 
.A(n_1168),
.B(n_1046),
.C(n_1043),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1174),
.B(n_1084),
.Y(n_1190)
);

NOR3x1_ASAP7_75t_L g1191 ( 
.A(n_1176),
.B(n_1043),
.C(n_1008),
.Y(n_1191)
);

NOR2x1_ASAP7_75t_SL g1192 ( 
.A(n_1171),
.B(n_1084),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_1166),
.B(n_1007),
.C(n_1013),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_L g1194 ( 
.A(n_1179),
.B(n_1007),
.C(n_1013),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1181),
.B(n_1086),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1178),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_L g1197 ( 
.A(n_1175),
.B(n_1007),
.C(n_1013),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1170),
.B(n_1008),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1182),
.Y(n_1199)
);

OAI211xp5_ASAP7_75t_L g1200 ( 
.A1(n_1184),
.A2(n_1180),
.B(n_1165),
.C(n_1086),
.Y(n_1200)
);

NAND4xp25_ASAP7_75t_SL g1201 ( 
.A(n_1183),
.B(n_1026),
.C(n_953),
.D(n_1061),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1186),
.B(n_956),
.C(n_953),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1196),
.B(n_1008),
.C(n_941),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1192),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1188),
.B(n_1007),
.C(n_1013),
.Y(n_1205)
);

NAND4xp75_ASAP7_75t_L g1206 ( 
.A(n_1185),
.B(n_1024),
.C(n_1041),
.D(n_1026),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1187),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1190),
.A2(n_1043),
.B1(n_1026),
.B2(n_1048),
.Y(n_1208)
);

OAI211xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1195),
.A2(n_1069),
.B(n_1048),
.C(n_1017),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1198),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1197),
.B(n_922),
.Y(n_1211)
);

NOR3xp33_ASAP7_75t_L g1212 ( 
.A(n_1193),
.B(n_969),
.C(n_966),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1191),
.B(n_1048),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1194),
.B(n_956),
.C(n_922),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1198),
.A2(n_1189),
.B1(n_1041),
.B2(n_981),
.Y(n_1215)
);

NAND4xp25_ASAP7_75t_L g1216 ( 
.A(n_1184),
.B(n_1041),
.C(n_1050),
.D(n_927),
.Y(n_1216)
);

AOI311xp33_ASAP7_75t_L g1217 ( 
.A1(n_1183),
.A2(n_1039),
.A3(n_1032),
.B(n_1031),
.C(n_1027),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1182),
.Y(n_1218)
);

AND4x2_ASAP7_75t_L g1219 ( 
.A(n_1190),
.B(n_1017),
.C(n_994),
.D(n_964),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_L g1220 ( 
.A(n_1182),
.B(n_927),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1183),
.B(n_994),
.Y(n_1221)
);

OAI211xp5_ASAP7_75t_L g1222 ( 
.A1(n_1182),
.A2(n_994),
.B(n_966),
.C(n_964),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1210),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1199),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1218),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1204),
.A2(n_994),
.B1(n_1014),
.B2(n_1050),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1207),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1220),
.B(n_994),
.Y(n_1228)
);

NOR2x1_ASAP7_75t_L g1229 ( 
.A(n_1216),
.B(n_892),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1221),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1202),
.B(n_994),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1213),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1208),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1200),
.B(n_932),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1215),
.B(n_1050),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1201),
.Y(n_1236)
);

NOR3xp33_ASAP7_75t_L g1237 ( 
.A(n_1209),
.B(n_913),
.C(n_914),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1219),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1203),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1211),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1206),
.Y(n_1241)
);

AO22x2_ASAP7_75t_L g1242 ( 
.A1(n_1205),
.A2(n_1017),
.B1(n_892),
.B2(n_913),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1205),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1212),
.A2(n_1022),
.B1(n_1014),
.B2(n_932),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1217),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1214),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1225),
.B(n_1222),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1224),
.B(n_1022),
.Y(n_1248)
);

XNOR2xp5_ASAP7_75t_L g1249 ( 
.A(n_1239),
.B(n_1014),
.Y(n_1249)
);

NOR2x1_ASAP7_75t_L g1250 ( 
.A(n_1223),
.B(n_932),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1234),
.A2(n_964),
.B(n_1039),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1227),
.B(n_932),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1236),
.A2(n_1022),
.B(n_1039),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1241),
.A2(n_1022),
.B(n_909),
.Y(n_1254)
);

XNOR2xp5_ASAP7_75t_L g1255 ( 
.A(n_1240),
.B(n_909),
.Y(n_1255)
);

XNOR2x1_ASAP7_75t_L g1256 ( 
.A(n_1246),
.B(n_1238),
.Y(n_1256)
);

NAND4xp75_ASAP7_75t_L g1257 ( 
.A(n_1230),
.B(n_1025),
.C(n_1032),
.D(n_1031),
.Y(n_1257)
);

NOR4xp75_ASAP7_75t_SL g1258 ( 
.A(n_1226),
.B(n_1022),
.C(n_887),
.D(n_937),
.Y(n_1258)
);

NOR3xp33_ASAP7_75t_L g1259 ( 
.A(n_1232),
.B(n_1027),
.C(n_1010),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1233),
.A2(n_1032),
.B1(n_1031),
.B2(n_1027),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1243),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1242),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1228),
.Y(n_1263)
);

NAND4xp25_ASAP7_75t_L g1264 ( 
.A(n_1245),
.B(n_1022),
.C(n_1010),
.D(n_999),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1229),
.Y(n_1265)
);

NAND4xp75_ASAP7_75t_L g1266 ( 
.A(n_1244),
.B(n_1025),
.C(n_1010),
.D(n_1021),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1235),
.B(n_1047),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1242),
.Y(n_1268)
);

XOR2x2_ASAP7_75t_L g1269 ( 
.A(n_1256),
.B(n_1237),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1252),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1261),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1261),
.Y(n_1272)
);

XNOR2x1_ASAP7_75t_L g1273 ( 
.A(n_1247),
.B(n_1244),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1262),
.A2(n_1231),
.B1(n_1047),
.B2(n_979),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1263),
.B(n_1231),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1268),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1250),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1257),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1248),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1255),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1267),
.Y(n_1281)
);

XNOR2x1_ASAP7_75t_L g1282 ( 
.A(n_1249),
.B(n_980),
.Y(n_1282)
);

XNOR2xp5_ASAP7_75t_L g1283 ( 
.A(n_1264),
.B(n_156),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1271),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1275),
.B(n_1265),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1272),
.Y(n_1286)
);

AOI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1272),
.A2(n_1278),
.B1(n_1270),
.B2(n_1277),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1281),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1282),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1279),
.A2(n_1253),
.B1(n_1251),
.B2(n_1260),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1273),
.A2(n_1254),
.B1(n_1259),
.B2(n_1266),
.Y(n_1291)
);

OR3x1_ASAP7_75t_L g1292 ( 
.A(n_1277),
.B(n_1258),
.C(n_979),
.Y(n_1292)
);

XOR2xp5_ASAP7_75t_L g1293 ( 
.A(n_1269),
.B(n_159),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1276),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1274),
.A2(n_1047),
.B1(n_887),
.B2(n_1000),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1283),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1280),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1272),
.Y(n_1298)
);

AOI211xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1285),
.A2(n_162),
.B(n_192),
.C(n_1025),
.Y(n_1299)
);

NOR4xp25_ASAP7_75t_L g1300 ( 
.A(n_1294),
.B(n_978),
.C(n_977),
.D(n_1011),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1288),
.B(n_1286),
.Y(n_1301)
);

AOI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1290),
.A2(n_978),
.B1(n_977),
.B2(n_970),
.C(n_1011),
.Y(n_1302)
);

OAI322xp33_ASAP7_75t_L g1303 ( 
.A1(n_1297),
.A2(n_1009),
.A3(n_1035),
.B1(n_1018),
.B2(n_1015),
.C1(n_1011),
.C2(n_1012),
.Y(n_1303)
);

NAND4xp25_ASAP7_75t_L g1304 ( 
.A(n_1284),
.B(n_999),
.C(n_980),
.D(n_1021),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1287),
.B(n_1298),
.C(n_1296),
.Y(n_1305)
);

NAND4xp25_ASAP7_75t_L g1306 ( 
.A(n_1291),
.B(n_999),
.C(n_1021),
.D(n_975),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1289),
.B(n_1293),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_SL g1308 ( 
.A(n_1291),
.B(n_1000),
.C(n_1035),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_L g1309 ( 
.A(n_1305),
.B(n_1295),
.C(n_1292),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1301),
.A2(n_887),
.B1(n_1000),
.B2(n_1009),
.Y(n_1310)
);

OA22x2_ASAP7_75t_L g1311 ( 
.A1(n_1307),
.A2(n_999),
.B1(n_1035),
.B2(n_1018),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1299),
.A2(n_1000),
.B(n_1035),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1302),
.A2(n_1304),
.B1(n_1306),
.B2(n_1308),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1300),
.B(n_1009),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_L g1315 ( 
.A(n_1309),
.B(n_1303),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1313),
.A2(n_937),
.B(n_1009),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1312),
.A2(n_937),
.B(n_1011),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1314),
.A2(n_1310),
.B(n_1311),
.Y(n_1318)
);

AOI222xp33_ASAP7_75t_L g1319 ( 
.A1(n_1315),
.A2(n_1012),
.B1(n_1018),
.B2(n_1015),
.C1(n_970),
.C2(n_1045),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1319),
.A2(n_1318),
.B(n_1316),
.Y(n_1320)
);

AOI322xp5_ASAP7_75t_L g1321 ( 
.A1(n_1320),
.A2(n_1317),
.A3(n_1012),
.B1(n_1015),
.B2(n_1018),
.C1(n_1042),
.C2(n_1037),
.Y(n_1321)
);

AOI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1321),
.A2(n_891),
.B1(n_1015),
.B2(n_1012),
.C(n_1045),
.Y(n_1322)
);

AOI211xp5_ASAP7_75t_L g1323 ( 
.A1(n_1322),
.A2(n_891),
.B(n_975),
.C(n_987),
.Y(n_1323)
);


endmodule