module fake_jpeg_20420_n_395 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_38),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_49),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_22),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_15),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_60),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_63),
.Y(n_101)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_65),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_33),
.B1(n_23),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_90),
.B1(n_102),
.B2(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_81),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_33),
.B1(n_23),
.B2(n_29),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_89),
.B1(n_25),
.B2(n_24),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_26),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_37),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_96),
.Y(n_142)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_33),
.B1(n_23),
.B2(n_26),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_33),
.B1(n_58),
.B2(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_46),
.A2(n_29),
.B1(n_16),
.B2(n_17),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_29),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_16),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_36),
.B(n_17),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_17),
.B1(n_32),
.B2(n_28),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_110),
.B1(n_112),
.B2(n_125),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_109),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_32),
.B1(n_20),
.B2(n_28),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_32),
.B1(n_20),
.B2(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_30),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_71),
.C(n_74),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_129),
.B1(n_134),
.B2(n_141),
.Y(n_150)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_22),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_82),
.Y(n_152)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_99),
.B1(n_70),
.B2(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_22),
.B1(n_30),
.B2(n_14),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_136),
.B1(n_145),
.B2(n_146),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_66),
.Y(n_179)
);

BUFx24_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_91),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_144),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_72),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_71),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_81),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_148),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_68),
.B(n_88),
.C(n_97),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_80),
.A3(n_68),
.B1(n_88),
.B2(n_79),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_153),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_133),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_108),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_159),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_102),
.B1(n_100),
.B2(n_69),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_163),
.B1(n_165),
.B2(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_127),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_69),
.B1(n_85),
.B2(n_84),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_115),
.C(n_140),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_93),
.B1(n_104),
.B2(n_98),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_98),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_92),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_92),
.B1(n_82),
.B2(n_75),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_92),
.B1(n_86),
.B2(n_103),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_177),
.B1(n_180),
.B2(n_137),
.Y(n_210)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_117),
.A2(n_86),
.B1(n_103),
.B2(n_66),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_137),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_66),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_107),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_119),
.B(n_138),
.C(n_139),
.D(n_137),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_136),
.B1(n_138),
.B2(n_107),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_186),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_142),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_142),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_188),
.B(n_196),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_167),
.C(n_147),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_139),
.B(n_115),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_194),
.A2(n_217),
.B(n_10),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_139),
.B1(n_125),
.B2(n_146),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_195),
.A2(n_201),
.B1(n_219),
.B2(n_221),
.Y(n_248)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_204),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_208),
.C(n_163),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_155),
.B(n_110),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_199),
.B(n_202),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_223),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_132),
.B1(n_112),
.B2(n_143),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_143),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_131),
.B1(n_126),
.B2(n_123),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_210),
.B1(n_182),
.B2(n_168),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_111),
.C(n_123),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_130),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_205),
.B(n_206),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_111),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_66),
.C(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_218),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_150),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_214),
.A2(n_154),
.B1(n_161),
.B2(n_162),
.Y(n_227)
);

BUFx24_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_5),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_156),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_152),
.B(n_7),
.C(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_152),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_154),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_10),
.Y(n_223)
);

OAI211xp5_ASAP7_75t_L g274 ( 
.A1(n_224),
.A2(n_234),
.B(n_190),
.C(n_173),
.Y(n_274)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_237),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_227),
.A2(n_229),
.B1(n_230),
.B2(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_150),
.B1(n_176),
.B2(n_149),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_157),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_233),
.A2(n_258),
.B1(n_190),
.B2(n_10),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_148),
.Y(n_234)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_241),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_152),
.B(n_181),
.C(n_165),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_214),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_172),
.B1(n_174),
.B2(n_169),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_247),
.B1(n_197),
.B2(n_186),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_178),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_249),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_201),
.B1(n_186),
.B2(n_222),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_178),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_180),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_257),
.Y(n_285)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_182),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_261),
.A2(n_271),
.B1(n_230),
.B2(n_227),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_218),
.C(n_194),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_232),
.C(n_231),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_202),
.A3(n_198),
.B1(n_193),
.B2(n_192),
.C1(n_221),
.C2(n_212),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g312 ( 
.A(n_266),
.B(n_282),
.C(n_263),
.Y(n_312)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_251),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_217),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_274),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_200),
.B1(n_220),
.B2(n_211),
.Y(n_271)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_228),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_284),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_256),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_246),
.B1(n_256),
.B2(n_236),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_272),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_283),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_232),
.C(n_239),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_299),
.C(n_284),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_248),
.B1(n_252),
.B2(n_235),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_293),
.A2(n_287),
.B1(n_263),
.B2(n_285),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_235),
.B(n_233),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_296),
.A2(n_306),
.B(n_309),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_233),
.C(n_247),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_311),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_271),
.A2(n_243),
.B1(n_249),
.B2(n_241),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_300),
.B1(n_296),
.B2(n_299),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_265),
.A2(n_226),
.B(n_237),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_253),
.B(n_12),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_262),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_265),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_324),
.Y(n_340)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_315),
.A2(n_333),
.B1(n_314),
.B2(n_324),
.Y(n_338)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_330),
.C(n_332),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_318),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_321),
.Y(n_347)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_322),
.B(n_323),
.Y(n_341)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_285),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_308),
.Y(n_325)
);

INVx11_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_326),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_329),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_270),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_260),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_259),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_303),
.C(n_311),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_343),
.C(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_306),
.B(n_292),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_290),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_308),
.C(n_294),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_319),
.A2(n_293),
.B1(n_309),
.B2(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_344),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_328),
.A2(n_279),
.B(n_278),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_348),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_349),
.B(n_330),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_350),
.B(n_334),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_335),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_355),
.Y(n_373)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_362),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_334),
.Y(n_363)
);

AO221x1_ASAP7_75t_L g358 ( 
.A1(n_345),
.A2(n_260),
.B1(n_297),
.B2(n_273),
.C(n_331),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_359),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_346),
.A2(n_322),
.B1(n_288),
.B2(n_268),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_361),
.A2(n_342),
.B1(n_336),
.B2(n_295),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_317),
.C(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_363),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_338),
.B1(n_347),
.B2(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_366),
.B(n_367),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_347),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_368),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_340),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_369),
.A2(n_370),
.B(n_372),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_340),
.Y(n_370)
);

NAND4xp25_ASAP7_75t_SL g375 ( 
.A(n_371),
.B(n_352),
.C(n_346),
.D(n_354),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_376),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_373),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_380),
.B(n_371),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_378),
.A2(n_362),
.B1(n_337),
.B2(n_339),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_384),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_381),
.A2(n_342),
.B1(n_336),
.B2(n_366),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_385),
.B(n_386),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_379),
.A2(n_374),
.B(n_377),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_367),
.C(n_363),
.Y(n_387)
);

OAI311xp33_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_365),
.A3(n_359),
.B1(n_313),
.C1(n_315),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_390),
.B(n_382),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_391),
.A2(n_392),
.B(n_389),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_385),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_393),
.A2(n_281),
.B1(n_276),
.B2(n_277),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_327),
.Y(n_395)
);


endmodule