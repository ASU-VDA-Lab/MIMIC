module fake_jpeg_22657_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_23),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_58),
.B1(n_32),
.B2(n_20),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_18),
.B1(n_25),
.B2(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_65),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_31),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_25),
.B1(n_18),
.B2(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_76),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_22),
.B1(n_30),
.B2(n_35),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_77),
.A2(n_86),
.B1(n_90),
.B2(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_36),
.Y(n_78)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_40),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_60),
.C(n_48),
.Y(n_102)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_24),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_42),
.B1(n_41),
.B2(n_43),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_0),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_20),
.B(n_24),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_89),
.B(n_87),
.Y(n_133)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_74),
.C(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_112),
.Y(n_137)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_110),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_108),
.Y(n_156)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_66),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_124),
.B1(n_91),
.B2(n_93),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_50),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_40),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_93),
.B1(n_17),
.B2(n_79),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_34),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_19),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_61),
.B1(n_57),
.B2(n_51),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_83),
.B1(n_88),
.B2(n_84),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_143),
.B1(n_145),
.B2(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_153),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_136),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_142),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_87),
.B(n_89),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_84),
.B(n_80),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_93),
.B1(n_87),
.B2(n_75),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_75),
.B1(n_91),
.B2(n_76),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_69),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_102),
.B1(n_112),
.B2(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_152),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_121),
.B(n_114),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_120),
.C(n_100),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_175),
.C(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_121),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_134),
.B(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_189),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_125),
.C(n_123),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_130),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_118),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_185),
.B(n_138),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_114),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_111),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_111),
.B(n_126),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_36),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_149),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_188),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_135),
.B1(n_152),
.B2(n_148),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_216),
.B1(n_158),
.B2(n_160),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_199),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_212),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_144),
.B(n_133),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_208),
.B(n_185),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_151),
.B1(n_116),
.B2(n_79),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_158),
.B1(n_166),
.B2(n_168),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_49),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_17),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_21),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_162),
.A2(n_104),
.B1(n_113),
.B2(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_167),
.B(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_227),
.B1(n_228),
.B2(n_233),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_190),
.A2(n_169),
.B1(n_175),
.B2(n_177),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_167),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_235),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_190),
.A2(n_169),
.B1(n_174),
.B2(n_179),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_132),
.B1(n_128),
.B2(n_104),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_239),
.B1(n_243),
.B2(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_242),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_107),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_43),
.B1(n_49),
.B2(n_69),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_107),
.B1(n_109),
.B2(n_23),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_204),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_204),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_194),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_267),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_207),
.B1(n_216),
.B2(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_213),
.B1(n_200),
.B2(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_198),
.C(n_196),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_260),
.C(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_197),
.C(n_208),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_241),
.C(n_219),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_208),
.C(n_205),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_212),
.C(n_201),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_266),
.C(n_23),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_192),
.C(n_109),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_192),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_221),
.B1(n_245),
.B2(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_272),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_250),
.A2(n_234),
.B1(n_214),
.B2(n_23),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_278),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_9),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_107),
.C(n_1),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_283),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_262),
.B(n_260),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_285),
.A2(n_286),
.B(n_9),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_274),
.B(n_284),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_295),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_288),
.B(n_289),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_267),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_258),
.B(n_248),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_296),
.B(n_10),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_276),
.B(n_263),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_271),
.B(n_270),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_247),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_263),
.C(n_9),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_8),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_279),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_300),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_302),
.B(n_309),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_0),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_11),
.B(n_15),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_306),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_312),
.B1(n_5),
.B2(n_7),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_11),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_311),
.B(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_289),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_12),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_322),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_293),
.C(n_2),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_320),
.C(n_321),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_303),
.C(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_1),
.C(n_2),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_5),
.C(n_7),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_328),
.B(n_329),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_330),
.B(n_4),
.C(n_326),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_327),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_15),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_14),
.C(n_4),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_314),
.B1(n_321),
.B2(n_14),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.C(n_333),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_330),
.CI(n_335),
.CON(n_337),
.SN(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_317),
.Y(n_338)
);


endmodule