module fake_jpeg_24206_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_20),
.Y(n_57)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_38),
.B(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_64),
.B(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_17),
.B1(n_33),
.B2(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_79),
.B1(n_40),
.B2(n_47),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_23),
.B1(n_33),
.B2(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_26),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_26),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_89),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_70),
.B1(n_75),
.B2(n_58),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_96),
.B1(n_108),
.B2(n_109),
.Y(n_132)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_30),
.B1(n_19),
.B2(n_22),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_49),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_56),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_30),
.B1(n_19),
.B2(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_31),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_44),
.C(n_34),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_83),
.C(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_102),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_34),
.B1(n_27),
.B2(n_18),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_27),
.B1(n_18),
.B2(n_44),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_95),
.B1(n_86),
.B2(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_121),
.B1(n_123),
.B2(n_133),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_60),
.Y(n_115)
);

OAI221xp5_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_116),
.B1(n_122),
.B2(n_129),
.C(n_15),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_75),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_67),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_56),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_134),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_74),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_89),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_58),
.B1(n_48),
.B2(n_31),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_48),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_85),
.A2(n_31),
.B(n_20),
.C(n_68),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_105),
.B1(n_87),
.B2(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_97),
.B1(n_91),
.B2(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_1),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_158),
.B(n_134),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_140),
.B(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_151),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_97),
.B1(n_80),
.B2(n_20),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_159),
.B1(n_161),
.B2(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_63),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_160),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_124),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_20),
.B1(n_101),
.B2(n_98),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_98),
.B1(n_101),
.B2(n_3),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_98),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_101),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_166),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_171),
.B1(n_116),
.B2(n_143),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_126),
.B(n_120),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_167),
.B(n_161),
.Y(n_188)
);

XNOR2x2_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_129),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_116),
.B1(n_151),
.B2(n_122),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_129),
.B1(n_132),
.B2(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_115),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_110),
.C(n_113),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

OAI322xp33_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_141),
.A3(n_147),
.B1(n_144),
.B2(n_142),
.C1(n_153),
.C2(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_183),
.Y(n_207)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_138),
.B1(n_152),
.B2(n_154),
.C(n_139),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_139),
.C(n_123),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_189),
.C(n_179),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_195),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_148),
.C(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_159),
.B1(n_145),
.B2(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_168),
.B1(n_173),
.B2(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_196),
.B1(n_7),
.B2(n_8),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_149),
.B(n_115),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_172),
.B(n_175),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_166),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_174),
.B1(n_173),
.B2(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_210),
.B1(n_10),
.B2(n_11),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_172),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_204),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_164),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_193),
.B(n_188),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_1),
.C(n_4),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_185),
.B1(n_189),
.B2(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_10),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_194),
.B1(n_191),
.B2(n_185),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_186),
.B1(n_183),
.B2(n_182),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_218),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_207),
.A2(n_186),
.B(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_11),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_205),
.B1(n_207),
.B2(n_202),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_226),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_208),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_213),
.Y(n_229)
);

AOI31xp67_ASAP7_75t_SL g228 ( 
.A1(n_226),
.A2(n_215),
.A3(n_217),
.B(n_216),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_214),
.B(n_222),
.C(n_232),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_225),
.B(n_221),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_218),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_213),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_235),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_13),
.C(n_15),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_11),
.C(n_13),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_13),
.B(n_15),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_240),
.Y(n_242)
);


endmodule