module fake_jpeg_7687_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_62),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_2),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_46),
.B1(n_53),
.B2(n_52),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_46),
.B1(n_54),
.B2(n_50),
.Y(n_72)
);

AOI222xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.C1(n_77),
.C2(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_52),
.B1(n_50),
.B2(n_45),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_45),
.B1(n_43),
.B2(n_26),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_24),
.B1(n_36),
.B2(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_13),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_38),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_89),
.B(n_92),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_17),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_90),
.B(n_93),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_90),
.B1(n_95),
.B2(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_97),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_87),
.B1(n_78),
.B2(n_68),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_91),
.B1(n_75),
.B2(n_70),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_89),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_67),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_18),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_20),
.C(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_22),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_27),
.B(n_28),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_30),
.B(n_31),
.Y(n_110)
);

NAND2x1_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_94),
.Y(n_111)
);


endmodule