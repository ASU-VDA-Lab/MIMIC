module fake_jpeg_2225_n_162 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_29),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_45),
.B(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_18),
.B1(n_16),
.B2(n_22),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_24),
.A2(n_13),
.B1(n_26),
.B2(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_57),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_14),
.C(n_26),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_58),
.C(n_7),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_14),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_35),
.C(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_22),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_18),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_2),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_5),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_47),
.Y(n_101)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_95),
.B1(n_73),
.B2(n_55),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_96),
.B1(n_60),
.B2(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_9),
.B1(n_10),
.B2(n_48),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_52),
.A3(n_72),
.B1(n_51),
.B2(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_85),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_48),
.B1(n_62),
.B2(n_59),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_91),
.B1(n_90),
.B2(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_62),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_80),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_59),
.B(n_61),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_61),
.B(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_75),
.C(n_88),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_125),
.C(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_127),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_112),
.B(n_106),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_84),
.C(n_74),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_113),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_136),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_104),
.B(n_97),
.C(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_137),
.Y(n_138)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_100),
.A3(n_97),
.B1(n_115),
.B2(n_123),
.C(n_126),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_103),
.B1(n_118),
.B2(n_107),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_144),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_130),
.A2(n_118),
.B(n_122),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_143),
.B(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_132),
.C(n_131),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_143),
.B1(n_136),
.B2(n_138),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_137),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_141),
.C(n_113),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_140),
.B(n_128),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_103),
.B1(n_110),
.B2(n_114),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_146),
.A3(n_148),
.B1(n_153),
.B2(n_94),
.C1(n_86),
.C2(n_55),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_86),
.A3(n_102),
.B1(n_10),
.B2(n_93),
.C1(n_89),
.C2(n_69),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_156),
.B(n_159),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_156),
.Y(n_162)
);


endmodule