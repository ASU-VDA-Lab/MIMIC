module fake_netlist_5_2490_n_1811 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1811);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1811;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g161 ( 
.A(n_47),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_26),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_68),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_57),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_113),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_98),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_27),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_34),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_109),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_46),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_15),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_79),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_145),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_35),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_55),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_64),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_33),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_24),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_126),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_51),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_140),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_38),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_25),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_90),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_70),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_45),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_39),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_28),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_111),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_43),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_4),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_43),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_25),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_89),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_120),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_27),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_36),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_41),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_5),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_154),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_76),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_18),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_55),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_149),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_15),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_107),
.Y(n_230)
);

BUFx2_ASAP7_75t_SL g231 ( 
.A(n_56),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_155),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_2),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_72),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_18),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_86),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_67),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_29),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_100),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_121),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_4),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_73),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_46),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_53),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_78),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_36),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_96),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_84),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_53),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_93),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_102),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_153),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_88),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_40),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_115),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_105),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_159),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_135),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_60),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_32),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_57),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_104),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_85),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_74),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_60),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_129),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_118),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_142),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_12),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_134),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_77),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_64),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_136),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_54),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_39),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_58),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_29),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_103),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_48),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_10),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_94),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_71),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_110),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_147),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_69),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_108),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_17),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_19),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_13),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_66),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_119),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_137),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_22),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_48),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_92),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_9),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_24),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_165),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_203),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_203),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_203),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_185),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_186),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_167),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_203),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_173),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_R g329 ( 
.A(n_163),
.B(n_0),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_203),
.B(n_0),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_174),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_177),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_229),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_179),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_184),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_203),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_161),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_194),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_161),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_190),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_196),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_193),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_201),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_161),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_197),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_202),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_188),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_197),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_168),
.B(n_1),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_228),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_208),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_214),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_188),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_222),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_188),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_227),
.Y(n_358)
);

BUFx6f_ASAP7_75t_SL g359 ( 
.A(n_172),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_210),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_232),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_168),
.B(n_1),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_210),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_239),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_240),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_172),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_235),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_295),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_307),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_247),
.B(n_305),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_245),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_210),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_175),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_265),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_314),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_252),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_258),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_260),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_233),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_266),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_175),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_265),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_265),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_193),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_193),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_215),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_189),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_229),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_270),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_271),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_207),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_274),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_276),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_247),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

BUFx8_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_221),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_305),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_337),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_393),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_162),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_172),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_182),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_351),
.B(n_233),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_205),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_286),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_362),
.B(n_315),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_330),
.B(n_182),
.Y(n_426)
);

AOI22x1_ASAP7_75t_L g427 ( 
.A1(n_345),
.A2(n_350),
.B1(n_370),
.B2(n_369),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_360),
.A2(n_192),
.B(n_189),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_337),
.B(n_277),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_320),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_281),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_363),
.A2(n_200),
.B(n_192),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_280),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_333),
.B(n_315),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_333),
.B(n_182),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_339),
.B(n_182),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_385),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_385),
.B(n_207),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_207),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_330),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_326),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_278),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_328),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_375),
.B(n_288),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_347),
.B(n_216),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_426),
.A2(n_368),
.B1(n_347),
.B2(n_236),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_370),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_430),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_331),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_412),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_464),
.A2(n_417),
.B1(n_423),
.B2(n_415),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_231),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_464),
.B(n_332),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_458),
.B(n_462),
.Y(n_482)
);

BUFx4f_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_458),
.B(n_334),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_164),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_397),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_458),
.B(n_335),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_415),
.B(n_340),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_458),
.B(n_462),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_458),
.B(n_341),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_423),
.A2(n_329),
.B1(n_294),
.B2(n_285),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_437),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_433),
.B(n_401),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_426),
.A2(n_368),
.B1(n_259),
.B2(n_236),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_411),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_458),
.B(n_343),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_411),
.Y(n_502)
);

OR2x6_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_231),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_443),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_402),
.B(n_346),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_437),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_449),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_397),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_462),
.B(n_353),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_426),
.A2(n_259),
.B1(n_236),
.B2(n_204),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_462),
.B(n_354),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVx3_ASAP7_75t_R g520 ( 
.A(n_454),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_433),
.B(n_381),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_402),
.B(n_356),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_459),
.B(n_278),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

INVx6_ASAP7_75t_L g527 ( 
.A(n_401),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

BUFx4f_ASAP7_75t_L g529 ( 
.A(n_462),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_462),
.B(n_358),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_455),
.B(n_361),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_455),
.B(n_364),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_455),
.B(n_389),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_456),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_449),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_416),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_431),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_404),
.B(n_365),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_432),
.B(n_373),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_431),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_432),
.B(n_378),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_434),
.B(n_379),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_456),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_434),
.B(n_380),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_412),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_460),
.B(n_390),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_449),
.B(n_382),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_396),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_446),
.B(n_391),
.Y(n_554)
);

AND3x1_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_204),
.C(n_200),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_414),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_459),
.B(n_278),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

AO21x2_ASAP7_75t_L g560 ( 
.A1(n_420),
.A2(n_170),
.B(n_164),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_449),
.B(n_392),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_416),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_449),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_426),
.B(n_394),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_412),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_414),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_462),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_453),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_454),
.B(n_170),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_426),
.B(n_395),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_416),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_453),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_409),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_454),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_416),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_446),
.B(n_390),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_462),
.B(n_359),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_457),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_462),
.B(n_299),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_409),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_457),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_460),
.B(n_403),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_454),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_440),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_414),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_427),
.B(n_463),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_457),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_457),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_416),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_463),
.B(n_324),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_426),
.B(n_286),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_426),
.B(n_216),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_398),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_461),
.B(n_325),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_461),
.B(n_338),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_416),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_414),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_454),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_400),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_465),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_259),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_465),
.B(n_348),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_465),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

BUFx4f_ASAP7_75t_L g612 ( 
.A(n_426),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_466),
.B(n_352),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_398),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_451),
.Y(n_615)
);

OAI21xp33_ASAP7_75t_L g616 ( 
.A1(n_403),
.A2(n_219),
.B(n_212),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_466),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_460),
.B(n_171),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_612),
.B(n_401),
.Y(n_619)
);

BUFx6f_ASAP7_75t_SL g620 ( 
.A(n_512),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_552),
.B(n_426),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_511),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_475),
.B(n_445),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_509),
.B(n_426),
.Y(n_624)
);

AO221x1_ASAP7_75t_L g625 ( 
.A1(n_470),
.A2(n_169),
.B1(n_313),
.B2(n_286),
.C(n_251),
.Y(n_625)
);

AND2x4_ASAP7_75t_SL g626 ( 
.A(n_607),
.B(n_367),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_470),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_511),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_612),
.B(n_401),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_535),
.A2(n_426),
.B1(n_420),
.B2(n_427),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_478),
.A2(n_426),
.B1(n_371),
.B2(n_377),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_541),
.B(n_460),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_470),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_601),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_550),
.B(n_460),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_602),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_607),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_470),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_478),
.A2(n_183),
.B1(n_282),
.B2(n_283),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_612),
.B(n_401),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_569),
.B(n_401),
.Y(n_641)
);

AOI22x1_ASAP7_75t_L g642 ( 
.A1(n_468),
.A2(n_171),
.B1(n_176),
.B2(n_269),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_569),
.B(n_459),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_470),
.B(n_412),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_492),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_564),
.B(n_459),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_537),
.B(n_459),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_543),
.B(n_388),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_609),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_485),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_574),
.B(n_440),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_485),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_485),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_492),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_499),
.B(n_398),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_564),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_485),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_577),
.Y(n_659)
);

AOI221xp5_ASAP7_75t_L g660 ( 
.A1(n_616),
.A2(n_218),
.B1(n_217),
.B2(n_248),
.C(n_311),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_499),
.B(n_399),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_485),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_502),
.B(n_399),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_468),
.B(n_459),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_523),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_599),
.B(n_467),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_540),
.B(n_440),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_607),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_502),
.B(n_399),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_523),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_589),
.B(n_410),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_611),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_523),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_589),
.B(n_410),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_583),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_611),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_523),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_576),
.B(n_410),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_600),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_583),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_467),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_590),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_587),
.B(n_467),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_614),
.Y(n_686)
);

O2A1O1Ixp5_ASAP7_75t_L g687 ( 
.A1(n_593),
.A2(n_467),
.B(n_396),
.C(n_451),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_587),
.B(n_467),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_544),
.B(n_282),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_547),
.B(n_467),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_512),
.B(n_212),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_590),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_614),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_531),
.B(n_283),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_506),
.B(n_406),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_473),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_551),
.B(n_406),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_561),
.B(n_406),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_491),
.A2(n_303),
.B1(n_306),
.B2(n_317),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_610),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_532),
.B(n_486),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_557),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_611),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_486),
.B(n_406),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_486),
.B(n_524),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_486),
.B(n_406),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_481),
.B(n_554),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_473),
.B(n_406),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_474),
.B(n_407),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_515),
.B(n_286),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_610),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_483),
.A2(n_396),
.B(n_400),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_581),
.B(n_217),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_516),
.A2(n_427),
.B1(n_412),
.B2(n_451),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_534),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_504),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_515),
.B(n_286),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_534),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_605),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_563),
.B(n_218),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_495),
.A2(n_329),
.B1(n_261),
.B2(n_257),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_474),
.B(n_477),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_566),
.A2(n_253),
.B1(n_312),
.B2(n_181),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_477),
.B(n_407),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_489),
.B(n_407),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_597),
.B(n_617),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_489),
.B(n_407),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_546),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_490),
.B(n_407),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_515),
.B(n_476),
.Y(n_731)
);

NAND3x1_ASAP7_75t_L g732 ( 
.A(n_495),
.B(n_220),
.C(n_219),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_490),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_496),
.B(n_407),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_496),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_L g736 ( 
.A(n_469),
.B(n_178),
.C(n_166),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_510),
.B(n_513),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_546),
.Y(n_738)
);

NOR3xp33_ASAP7_75t_L g739 ( 
.A(n_487),
.B(n_248),
.C(n_191),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_515),
.B(n_476),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_539),
.B(n_180),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_504),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_515),
.B(n_286),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_539),
.B(n_195),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_515),
.B(n_476),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_548),
.B(n_451),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_510),
.B(n_428),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_513),
.B(n_428),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_542),
.B(n_198),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_548),
.B(n_451),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_483),
.A2(n_400),
.B(n_451),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_542),
.B(n_206),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_549),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_518),
.B(n_428),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_518),
.B(n_412),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_548),
.B(n_308),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_605),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_526),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_471),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_526),
.B(n_428),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_567),
.B(n_176),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_567),
.B(n_181),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_550),
.B(n_209),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_575),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_471),
.B(n_211),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_567),
.B(n_187),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_570),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_428),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_549),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_572),
.B(n_187),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_608),
.B(n_428),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_570),
.B(n_223),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_533),
.B(n_224),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_487),
.B(n_225),
.C(n_319),
.Y(n_774)
);

BUFx6f_ASAP7_75t_SL g775 ( 
.A(n_571),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_591),
.B(n_234),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_483),
.B(n_213),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_484),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_529),
.B(n_213),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_575),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_553),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_529),
.B(n_226),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_533),
.B(n_237),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_555),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_618),
.B(n_438),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_559),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_742),
.Y(n_787)
);

O2A1O1Ixp5_ASAP7_75t_L g788 ( 
.A1(n_777),
.A2(n_482),
.B(n_493),
.C(n_529),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_623),
.B(n_522),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_708),
.B(n_689),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_624),
.A2(n_672),
.B(n_643),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_703),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_621),
.A2(n_598),
.B(n_584),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_722),
.A2(n_616),
.B(n_501),
.C(n_517),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_703),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_634),
.B(n_488),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_672),
.A2(n_503),
.B(n_480),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_694),
.A2(n_514),
.B1(n_530),
.B2(n_494),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_702),
.A2(n_605),
.B1(n_615),
.B2(n_586),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_681),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_672),
.A2(n_503),
.B(n_480),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_717),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_723),
.A2(n_503),
.B(n_480),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_643),
.A2(n_503),
.B(n_480),
.Y(n_804)
);

OR2x2_ASAP7_75t_SL g805 ( 
.A(n_652),
.B(n_220),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_737),
.A2(n_503),
.B(n_480),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_706),
.A2(n_605),
.B1(n_615),
.B2(n_618),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_681),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_632),
.B(n_571),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_767),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_636),
.B(n_605),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_714),
.A2(n_498),
.B(n_571),
.C(n_565),
.Y(n_812)
);

OAI21xp33_ASAP7_75t_L g813 ( 
.A1(n_773),
.A2(n_555),
.B(n_243),
.Y(n_813)
);

OAI21xp33_ASAP7_75t_L g814 ( 
.A1(n_721),
.A2(n_246),
.B(n_238),
.Y(n_814)
);

O2A1O1Ixp5_ASAP7_75t_L g815 ( 
.A1(n_777),
.A2(n_571),
.B(n_559),
.C(n_565),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_628),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_650),
.B(n_615),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_628),
.B(n_615),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_746),
.A2(n_615),
.B(n_520),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_746),
.A2(n_520),
.B(n_560),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_750),
.A2(n_560),
.B(n_508),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_701),
.B(n_712),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_687),
.A2(n_579),
.B(n_578),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_750),
.A2(n_560),
.B(n_508),
.Y(n_824)
);

AO21x1_ASAP7_75t_L g825 ( 
.A1(n_779),
.A2(n_782),
.B(n_770),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_645),
.A2(n_508),
.B(n_472),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_645),
.A2(n_519),
.B(n_472),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_653),
.A2(n_519),
.B(n_472),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_635),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_759),
.B(n_497),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_727),
.B(n_680),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_647),
.A2(n_579),
.B(n_578),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_646),
.B(n_226),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_691),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_696),
.B(n_582),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_631),
.A2(n_527),
.B1(n_253),
.B2(n_267),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_668),
.A2(n_558),
.B1(n_525),
.B2(n_582),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_696),
.B(n_585),
.Y(n_838)
);

OAI321xp33_ASAP7_75t_L g839 ( 
.A1(n_639),
.A2(n_284),
.A3(n_275),
.B1(n_301),
.B2(n_300),
.C(n_289),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_673),
.A2(n_585),
.B(n_588),
.C(n_594),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_733),
.B(n_588),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_630),
.A2(n_527),
.B1(n_269),
.B2(n_256),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_731),
.A2(n_745),
.B(n_740),
.Y(n_843)
);

BUFx8_ASAP7_75t_L g844 ( 
.A(n_620),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_779),
.A2(n_782),
.B(n_770),
.C(n_666),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_699),
.B(n_249),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_763),
.A2(n_256),
.B(n_290),
.C(n_302),
.Y(n_847)
);

CKINVDCx10_ASAP7_75t_R g848 ( 
.A(n_620),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_784),
.B(n_254),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_731),
.A2(n_536),
.B(n_562),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_740),
.A2(n_536),
.B(n_562),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_745),
.A2(n_536),
.B(n_562),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_644),
.A2(n_558),
.B1(n_525),
.B2(n_595),
.Y(n_853)
);

OAI22x1_ASAP7_75t_L g854 ( 
.A1(n_649),
.A2(n_273),
.B1(n_255),
.B2(n_316),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_768),
.A2(n_594),
.B(n_595),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_776),
.B(n_262),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_751),
.A2(n_519),
.B(n_603),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_765),
.B(n_263),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_778),
.B(n_268),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_635),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_772),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_646),
.B(n_230),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_SL g863 ( 
.A1(n_761),
.A2(n_312),
.B(n_304),
.C(n_267),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_733),
.B(n_735),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_628),
.B(n_580),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_735),
.B(n_573),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_758),
.B(n_693),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_676),
.A2(n_257),
.B(n_304),
.C(n_302),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_783),
.B(n_272),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_622),
.A2(n_527),
.B1(n_290),
.B2(n_241),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_758),
.B(n_573),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_628),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_771),
.A2(n_558),
.B(n_525),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_747),
.A2(n_754),
.B(n_748),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_686),
.Y(n_875)
);

BUFx2_ASAP7_75t_SL g876 ( 
.A(n_775),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_666),
.A2(n_603),
.B(n_596),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_622),
.B(n_573),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_691),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_697),
.A2(n_603),
.B(n_596),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_622),
.B(n_596),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_698),
.A2(n_580),
.B(n_400),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_647),
.A2(n_580),
.B(n_405),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_657),
.A2(n_250),
.B1(n_241),
.B2(n_242),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_716),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_635),
.A2(n_525),
.B1(n_558),
.B2(n_412),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_757),
.A2(n_580),
.B(n_405),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_655),
.A2(n_230),
.B(n_250),
.C(n_244),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_651),
.B(n_654),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_651),
.B(n_479),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_741),
.B(n_287),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_720),
.B(n_580),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_756),
.A2(n_507),
.B(n_604),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_744),
.B(n_291),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_757),
.A2(n_405),
.B(n_606),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_651),
.B(n_479),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_749),
.B(n_292),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_757),
.A2(n_405),
.B(n_606),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_690),
.A2(n_405),
.B(n_592),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_720),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_654),
.B(n_500),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_L g902 ( 
.A1(n_752),
.A2(n_242),
.B(n_261),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_755),
.A2(n_405),
.B(n_592),
.Y(n_903)
);

OAI321xp33_ASAP7_75t_L g904 ( 
.A1(n_660),
.A2(n_289),
.A3(n_251),
.B1(n_264),
.B2(n_275),
.C(n_284),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_654),
.B(n_500),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_627),
.B(n_604),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_755),
.A2(n_568),
.B(n_505),
.Y(n_907)
);

OAI21xp33_ASAP7_75t_L g908 ( 
.A1(n_691),
.A2(n_310),
.B(n_309),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_764),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_683),
.A2(n_568),
.B(n_505),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_720),
.B(n_507),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_719),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_627),
.B(n_633),
.Y(n_913)
);

NOR2x1_ASAP7_75t_L g914 ( 
.A(n_635),
.B(n_244),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_729),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_700),
.B(n_298),
.C(n_293),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_637),
.B(n_521),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_764),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_633),
.B(n_521),
.Y(n_919)
);

AOI21xp33_ASAP7_75t_L g920 ( 
.A1(n_659),
.A2(n_318),
.B(n_301),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_667),
.A2(n_558),
.B1(n_525),
.B2(n_412),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_638),
.B(n_528),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_785),
.A2(n_528),
.B(n_556),
.C(n_545),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_685),
.A2(n_556),
.B(n_545),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_669),
.B(n_674),
.Y(n_925)
);

BUFx8_ASAP7_75t_L g926 ( 
.A(n_775),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_738),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_638),
.B(n_538),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_720),
.B(n_538),
.Y(n_929)
);

AND2x2_ASAP7_75t_SL g930 ( 
.A(n_715),
.B(n_264),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_658),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_658),
.B(n_525),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_662),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_688),
.A2(n_558),
.B(n_525),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_678),
.B(n_3),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_L g936 ( 
.A1(n_739),
.A2(n_293),
.B(n_297),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_662),
.B(n_438),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_704),
.B(n_3),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_724),
.A2(n_297),
.B(n_300),
.C(n_318),
.Y(n_939)
);

AO22x1_ASAP7_75t_L g940 ( 
.A1(n_774),
.A2(n_558),
.B1(n_412),
.B2(n_442),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_677),
.A2(n_412),
.B1(n_450),
.B2(n_421),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_665),
.B(n_450),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_682),
.A2(n_438),
.B(n_435),
.C(n_429),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_760),
.A2(n_438),
.B(n_421),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_684),
.A2(n_692),
.B(n_705),
.C(n_707),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_626),
.B(n_648),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_695),
.A2(n_419),
.B(n_447),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_665),
.B(n_438),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_671),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_671),
.A2(n_450),
.B1(n_421),
.B2(n_424),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_709),
.A2(n_438),
.B(n_425),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_675),
.B(n_435),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_675),
.B(n_679),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_736),
.B(n_435),
.C(n_424),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_679),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_756),
.A2(n_447),
.B(n_444),
.Y(n_956)
);

OAI22xp33_ASAP7_75t_L g957 ( 
.A1(n_656),
.A2(n_429),
.B1(n_424),
.B2(n_442),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_661),
.B(n_436),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_710),
.A2(n_436),
.B(n_425),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_761),
.A2(n_447),
.B(n_444),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_663),
.B(n_436),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_762),
.A2(n_447),
.B(n_444),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_762),
.A2(n_444),
.B(n_419),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_670),
.B(n_442),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_753),
.B(n_441),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_780),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_766),
.A2(n_441),
.B(n_439),
.C(n_429),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_766),
.A2(n_422),
.B(n_419),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_769),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_725),
.A2(n_422),
.B(n_419),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_726),
.A2(n_422),
.B(n_418),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_781),
.B(n_441),
.Y(n_972)
);

OAI321xp33_ASAP7_75t_L g973 ( 
.A1(n_641),
.A2(n_439),
.A3(n_425),
.B1(n_422),
.B2(n_418),
.C(n_9),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_626),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_809),
.A2(n_793),
.B(n_804),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_790),
.B(n_786),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_789),
.A2(n_641),
.B1(n_629),
.B2(n_619),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_810),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_787),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_791),
.A2(n_820),
.B(n_801),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_926),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_926),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_876),
.B(n_732),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_902),
.A2(n_640),
.B(n_629),
.C(n_619),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_831),
.A2(n_640),
.B(n_730),
.C(n_734),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_861),
.B(n_728),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_800),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_789),
.A2(n_798),
.B1(n_861),
.B2(n_796),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_844),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_802),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_966),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_811),
.B(n_732),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_955),
.B(n_664),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_811),
.B(n_625),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_900),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_L g996 ( 
.A(n_796),
.B(n_141),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_797),
.A2(n_713),
.B(n_718),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_966),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_909),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_817),
.B(n_891),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_918),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_808),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_794),
.A2(n_718),
.B(n_711),
.C(n_743),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_803),
.A2(n_743),
.B(n_711),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_806),
.A2(n_642),
.B(n_664),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_847),
.A2(n_439),
.B(n_418),
.C(n_7),
.Y(n_1006)
);

BUFx2_ASAP7_75t_SL g1007 ( 
.A(n_792),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_877),
.A2(n_418),
.B(n_664),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_829),
.B(n_664),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_795),
.B(n_664),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_858),
.B(n_5),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_879),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_821),
.A2(n_124),
.B(n_152),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_900),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_817),
.B(n_6),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_805),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_834),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_894),
.B(n_6),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_830),
.B(n_158),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_946),
.B(n_146),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_813),
.A2(n_7),
.B(n_8),
.C(n_11),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_930),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_SL g1023 ( 
.A(n_844),
.B(n_144),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_R g1024 ( 
.A(n_848),
.B(n_139),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_872),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_897),
.B(n_133),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_904),
.A2(n_14),
.B(n_16),
.C(n_20),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_930),
.B(n_21),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_859),
.B(n_114),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_846),
.B(n_822),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_859),
.B(n_21),
.C(n_22),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_869),
.A2(n_112),
.B1(n_95),
.B2(n_87),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_888),
.A2(n_23),
.B(n_26),
.C(n_30),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_957),
.A2(n_23),
.B(n_30),
.C(n_31),
.Y(n_1034)
);

O2A1O1Ixp5_ASAP7_75t_L g1035 ( 
.A1(n_825),
.A2(n_80),
.B(n_35),
.C(n_37),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_869),
.A2(n_812),
.B(n_845),
.C(n_856),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_925),
.B(n_31),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_974),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_955),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_846),
.B(n_37),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_824),
.A2(n_38),
.B(n_40),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_807),
.A2(n_799),
.B1(n_867),
.B2(n_933),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_849),
.B(n_41),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_833),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_849),
.B(n_42),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_856),
.A2(n_63),
.B1(n_49),
.B2(n_50),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_SL g1047 ( 
.A(n_936),
.B(n_45),
.C(n_50),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_933),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_885),
.B(n_52),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_842),
.A2(n_58),
.B(n_59),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_912),
.B(n_59),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_875),
.Y(n_1052)
);

NAND2x1p5_ASAP7_75t_L g1053 ( 
.A(n_816),
.B(n_61),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_916),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_915),
.B(n_62),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_927),
.B(n_969),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_788),
.A2(n_855),
.B(n_843),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_972),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_864),
.A2(n_837),
.B1(n_955),
.B2(n_945),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_931),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_955),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_958),
.B(n_961),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_957),
.A2(n_973),
.B(n_964),
.C(n_839),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_SL g1064 ( 
.A(n_829),
.B(n_860),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_913),
.A2(n_953),
.B(n_874),
.Y(n_1065)
);

INVx6_ASAP7_75t_L g1066 ( 
.A(n_833),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_965),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_944),
.A2(n_951),
.B(n_873),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_814),
.A2(n_938),
.B(n_935),
.C(n_819),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_925),
.B(n_908),
.Y(n_1070)
);

INVxp67_ASAP7_75t_SL g1071 ( 
.A(n_931),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_860),
.B(n_862),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_816),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_917),
.B(n_862),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_949),
.A2(n_836),
.B1(n_889),
.B2(n_818),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_935),
.A2(n_938),
.B(n_815),
.C(n_914),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_917),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_965),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_854),
.B(n_920),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_884),
.A2(n_870),
.A3(n_823),
.B1(n_868),
.B2(n_959),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_939),
.A2(n_954),
.B(n_943),
.C(n_863),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_934),
.A2(n_857),
.B(n_907),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_893),
.A2(n_865),
.B(n_911),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_826),
.A2(n_827),
.B(n_882),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_818),
.A2(n_932),
.B1(n_835),
.B2(n_838),
.Y(n_1085)
);

CKINVDCx6p67_ASAP7_75t_R g1086 ( 
.A(n_865),
.Y(n_1086)
);

INVx8_ASAP7_75t_L g1087 ( 
.A(n_940),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_954),
.A2(n_952),
.B1(n_886),
.B2(n_853),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_SL g1089 ( 
.A1(n_952),
.A2(n_948),
.B(n_937),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_937),
.B(n_948),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_950),
.B(n_841),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_942),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_878),
.A2(n_881),
.B(n_903),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_866),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_840),
.A2(n_880),
.B(n_956),
.C(n_883),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_929),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_906),
.B(n_919),
.Y(n_1097)
);

NAND2x1_ASAP7_75t_L g1098 ( 
.A(n_890),
.B(n_896),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_923),
.A2(n_967),
.B(n_911),
.C(n_892),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_892),
.A2(n_929),
.B1(n_871),
.B2(n_905),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_SL g1101 ( 
.A1(n_947),
.A2(n_899),
.B(n_924),
.C(n_910),
.Y(n_1101)
);

INVx3_ASAP7_75t_SL g1102 ( 
.A(n_832),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_970),
.A2(n_971),
.B(n_928),
.C(n_922),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_850),
.B(n_851),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_L g1105 ( 
.A(n_901),
.B(n_921),
.C(n_887),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_941),
.B(n_852),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_R g1107 ( 
.A(n_828),
.B(n_960),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_895),
.B(n_898),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_962),
.B(n_963),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_968),
.B(n_790),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_790),
.B(n_831),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_800),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_L g1113 ( 
.A1(n_790),
.A2(n_708),
.B(n_623),
.C(n_902),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_809),
.A2(n_612),
.B(n_529),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_790),
.B(n_634),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_790),
.A2(n_708),
.B1(n_623),
.B2(n_789),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_790),
.B(n_634),
.Y(n_1117)
);

CKINVDCx8_ASAP7_75t_R g1118 ( 
.A(n_848),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_966),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_790),
.B(n_831),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_966),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_966),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_978),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_975),
.A2(n_980),
.B(n_1114),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_1039),
.B(n_1009),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1084),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1061),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_979),
.B(n_1038),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_1022),
.B(n_1028),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1116),
.B(n_1115),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1061),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_988),
.A2(n_1113),
.B(n_1040),
.C(n_1117),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1058),
.B(n_976),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1000),
.B(n_1062),
.Y(n_1135)
);

AOI221x1_ASAP7_75t_L g1136 ( 
.A1(n_1041),
.A2(n_977),
.B1(n_1050),
.B2(n_1082),
.C(n_1005),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_1008),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1114),
.A2(n_1068),
.B(n_1005),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1030),
.B(n_990),
.Y(n_1139)
);

AO21x2_ASAP7_75t_L g1140 ( 
.A1(n_1057),
.A2(n_1068),
.B(n_997),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1093),
.A2(n_997),
.B(n_1098),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1103),
.A2(n_1109),
.B(n_1108),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1007),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1065),
.A2(n_1095),
.B(n_1004),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_984),
.A2(n_1110),
.B(n_985),
.Y(n_1145)
);

AO32x2_ASAP7_75t_L g1146 ( 
.A1(n_1059),
.A2(n_1042),
.A3(n_1075),
.B1(n_1048),
.B2(n_1085),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1076),
.A2(n_1100),
.A3(n_1069),
.B(n_1004),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1070),
.A2(n_1016),
.B1(n_1026),
.B2(n_1043),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1018),
.A2(n_1037),
.B(n_1054),
.C(n_1045),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_978),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1103),
.A2(n_1106),
.B(n_1099),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1041),
.A2(n_994),
.A3(n_1013),
.B(n_1015),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_984),
.A2(n_985),
.B(n_1101),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1092),
.B(n_986),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_993),
.A2(n_1091),
.B(n_1097),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1099),
.A2(n_1013),
.B(n_1003),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1104),
.A2(n_1003),
.B(n_1087),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1072),
.B(n_1009),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1063),
.A2(n_1056),
.B1(n_1074),
.B2(n_1027),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1021),
.A2(n_992),
.A3(n_1050),
.B(n_1090),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1039),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1012),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1077),
.B(n_1044),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1087),
.A2(n_1104),
.B(n_1105),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1010),
.A2(n_1081),
.B(n_1067),
.Y(n_1166)
);

AOI211x1_ASAP7_75t_L g1167 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1051),
.C(n_1055),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1081),
.A2(n_1078),
.B(n_1088),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1087),
.A2(n_1104),
.B(n_996),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1094),
.B(n_1002),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1063),
.A2(n_1029),
.B(n_1089),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1052),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_987),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1071),
.A2(n_1006),
.B(n_1039),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_982),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1112),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1107),
.A2(n_1019),
.B(n_1006),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_1025),
.B(n_995),
.Y(n_1178)
);

AOI21xp33_ASAP7_75t_L g1179 ( 
.A1(n_1027),
.A2(n_1034),
.B(n_1079),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1072),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_999),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1001),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1011),
.A2(n_1046),
.B(n_1032),
.C(n_1034),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_991),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1060),
.A2(n_1122),
.B(n_1121),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_989),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1020),
.A2(n_1035),
.B(n_1025),
.Y(n_1187)
);

AOI221x1_ASAP7_75t_L g1188 ( 
.A1(n_1080),
.A2(n_1119),
.B1(n_998),
.B2(n_1096),
.C(n_1073),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_983),
.A2(n_1102),
.B(n_1017),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1047),
.A2(n_1080),
.B(n_1086),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1061),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_995),
.B(n_1073),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1096),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1064),
.A2(n_1066),
.B1(n_983),
.B2(n_1023),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1053),
.A2(n_1033),
.B(n_1080),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1096),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_983),
.B(n_981),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1066),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1014),
.B(n_1053),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1014),
.B(n_1033),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1080),
.B(n_1024),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1118),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_990),
.Y(n_1203)
);

AO32x2_ASAP7_75t_L g1204 ( 
.A1(n_988),
.A2(n_1116),
.A3(n_977),
.B1(n_1059),
.B2(n_1042),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1056),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1084),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_975),
.A2(n_529),
.B(n_483),
.Y(n_1209)
);

OAI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1116),
.A2(n_790),
.B1(n_631),
.B2(n_636),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_975),
.A2(n_529),
.B(n_483),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_975),
.A2(n_529),
.B(n_483),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_L g1213 ( 
.A1(n_1113),
.A2(n_790),
.B(n_623),
.C(n_708),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1113),
.A2(n_708),
.B(n_623),
.C(n_790),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1072),
.B(n_1009),
.Y(n_1216)
);

O2A1O1Ixp5_ASAP7_75t_SL g1217 ( 
.A1(n_1116),
.A2(n_902),
.B(n_455),
.C(n_988),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_SL g1218 ( 
.A1(n_1041),
.A2(n_1050),
.B(n_1081),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1056),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1084),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1116),
.A2(n_623),
.B1(n_789),
.B2(n_708),
.Y(n_1221)
);

AO21x1_ASAP7_75t_L g1222 ( 
.A1(n_1116),
.A2(n_988),
.B(n_977),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1072),
.B(n_1009),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_1036),
.A2(n_790),
.B(n_1069),
.C(n_1021),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_980),
.A2(n_1036),
.A3(n_1057),
.B(n_975),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1039),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1057),
.A2(n_980),
.B(n_975),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1056),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1056),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_L g1231 ( 
.A(n_979),
.B(n_787),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1036),
.A2(n_569),
.B(n_619),
.Y(n_1232)
);

INVx4_ASAP7_75t_SL g1233 ( 
.A(n_1061),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1113),
.A2(n_708),
.B(n_623),
.C(n_790),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_988),
.A2(n_1116),
.A3(n_977),
.B1(n_1059),
.B2(n_1042),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1052),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1113),
.A2(n_1036),
.B(n_1116),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1116),
.B(n_634),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1056),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1116),
.B(n_634),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_980),
.A2(n_1057),
.B(n_975),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1057),
.A2(n_980),
.B(n_975),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_978),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1052),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1061),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_990),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_SL g1248 ( 
.A1(n_1041),
.A2(n_1050),
.B(n_1081),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_975),
.A2(n_529),
.B(n_483),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_978),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1115),
.B(n_1117),
.Y(n_1251)
);

AOI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1116),
.A2(n_623),
.B1(n_789),
.B2(n_714),
.C(n_988),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_975),
.A2(n_529),
.B(n_483),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1022),
.A2(n_649),
.B1(n_789),
.B2(n_623),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1056),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1084),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1257)
);

AOI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1116),
.A2(n_790),
.B(n_1113),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1072),
.B(n_1009),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_990),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1009),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_990),
.Y(n_1262)
);

OAI22x1_ASAP7_75t_L g1263 ( 
.A1(n_1046),
.A2(n_789),
.B1(n_478),
.B2(n_623),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1116),
.B(n_789),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_L g1265 ( 
.A(n_989),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1057),
.A2(n_980),
.B(n_975),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_1070),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_975),
.A2(n_529),
.B(n_483),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1084),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1084),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_978),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1226),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1251),
.B(n_1130),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1130),
.B(n_1205),
.Y(n_1274)
);

INVx6_ASAP7_75t_L g1275 ( 
.A(n_1226),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1163),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1168),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1254),
.A2(n_1252),
.B1(n_1131),
.B2(n_1221),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1263),
.A2(n_1240),
.B1(n_1238),
.B2(n_1134),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1180),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1252),
.A2(n_1129),
.B1(n_1148),
.B2(n_1264),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1183),
.A2(n_1179),
.B(n_1149),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1222),
.A2(n_1179),
.B1(n_1210),
.B2(n_1258),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1133),
.A2(n_1194),
.B(n_1237),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1258),
.A2(n_1237),
.B1(n_1190),
.B2(n_1160),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1176),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1190),
.A2(n_1160),
.B1(n_1135),
.B2(n_1171),
.Y(n_1287)
);

CKINVDCx11_ASAP7_75t_R g1288 ( 
.A(n_1202),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1205),
.A2(n_1207),
.B1(n_1247),
.B2(n_1257),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1172),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1135),
.A2(n_1171),
.B1(n_1134),
.B2(n_1247),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1202),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1158),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1214),
.B(n_1234),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1202),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1207),
.A2(n_1229),
.B1(n_1215),
.B2(n_1257),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1215),
.A2(n_1229),
.B1(n_1267),
.B2(n_1231),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1175),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1206),
.B(n_1219),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1218),
.A2(n_1248),
.B1(n_1267),
.B2(n_1228),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1201),
.A2(n_1143),
.B1(n_1177),
.B2(n_1255),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1216),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1230),
.B(n_1239),
.Y(n_1303)
);

INVx6_ASAP7_75t_L g1304 ( 
.A(n_1226),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1236),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1244),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1139),
.A2(n_1201),
.B1(n_1154),
.B2(n_1170),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1181),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_SL g1309 ( 
.A(n_1150),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1182),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1177),
.A2(n_1157),
.B1(n_1165),
.B2(n_1250),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1154),
.A2(n_1144),
.B1(n_1145),
.B2(n_1157),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1164),
.A2(n_1259),
.B1(n_1223),
.B2(n_1261),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1246),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1223),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1170),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1184),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1186),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1185),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1200),
.A2(n_1195),
.B1(n_1243),
.B2(n_1156),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1128),
.B2(n_1260),
.Y(n_1321)
);

INVxp33_ASAP7_75t_SL g1322 ( 
.A(n_1203),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1159),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1125),
.Y(n_1324)
);

INVx4_ASAP7_75t_L g1325 ( 
.A(n_1162),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1144),
.A2(n_1145),
.B1(n_1200),
.B2(n_1140),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1191),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1167),
.B(n_1203),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1193),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1260),
.A2(n_1197),
.B1(n_1265),
.B2(n_1271),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_1123),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1233),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1140),
.A2(n_1155),
.B1(n_1151),
.B2(n_1153),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1196),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1262),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1233),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1192),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1265),
.Y(n_1338)
);

OAI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1217),
.A2(n_1187),
.B(n_1189),
.Y(n_1339)
);

BUFx10_ASAP7_75t_L g1340 ( 
.A(n_1198),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1233),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1125),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1136),
.A2(n_1188),
.B1(n_1199),
.B2(n_1235),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1127),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1166),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1199),
.A2(n_1204),
.B1(n_1235),
.B2(n_1187),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1162),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1127),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1153),
.A2(n_1241),
.B1(n_1138),
.B2(n_1169),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1127),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1174),
.A2(n_1124),
.B(n_1235),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1232),
.A2(n_1174),
.B1(n_1192),
.B2(n_1178),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1224),
.A2(n_1211),
.B(n_1268),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1178),
.A2(n_1268),
.B1(n_1249),
.B2(n_1253),
.Y(n_1354)
);

CKINVDCx11_ASAP7_75t_R g1355 ( 
.A(n_1132),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1241),
.A2(n_1266),
.B1(n_1242),
.B2(n_1227),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1204),
.A2(n_1209),
.B(n_1253),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1225),
.Y(n_1358)
);

BUFx8_ASAP7_75t_SL g1359 ( 
.A(n_1132),
.Y(n_1359)
);

BUFx8_ASAP7_75t_L g1360 ( 
.A(n_1132),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1245),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1245),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1245),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1142),
.B(n_1266),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1227),
.A2(n_1242),
.B1(n_1204),
.B2(n_1213),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1146),
.A2(n_1126),
.B1(n_1269),
.B2(n_1256),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1161),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1161),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1209),
.A2(n_1212),
.B1(n_1249),
.B2(n_1211),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1208),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1220),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1152),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1270),
.B(n_1141),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1146),
.A2(n_1147),
.B1(n_1137),
.B2(n_1152),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1147),
.A2(n_1152),
.B1(n_1254),
.B2(n_1252),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1147),
.Y(n_1376)
);

INVx6_ASAP7_75t_L g1377 ( 
.A(n_1226),
.Y(n_1377)
);

BUFx8_ASAP7_75t_SL g1378 ( 
.A(n_1202),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1175),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1143),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1143),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1173),
.Y(n_1382)
);

BUFx8_ASAP7_75t_L g1383 ( 
.A(n_1202),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1173),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1202),
.Y(n_1385)
);

BUFx2_ASAP7_75t_SL g1386 ( 
.A(n_1231),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1202),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1163),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1254),
.A2(n_1252),
.B1(n_1131),
.B2(n_1221),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1173),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1252),
.A2(n_790),
.B1(n_478),
.B2(n_1116),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1221),
.A2(n_649),
.B(n_623),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1202),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1251),
.B(n_1130),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1254),
.A2(n_649),
.B1(n_789),
.B2(n_623),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1163),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1175),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1202),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1163),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1254),
.A2(n_1252),
.B1(n_1131),
.B2(n_1221),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1351),
.A2(n_1357),
.B(n_1353),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1367),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1339),
.A2(n_1285),
.B(n_1333),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1369),
.A2(n_1294),
.B(n_1343),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_SL g1405 ( 
.A1(n_1391),
.A2(n_1392),
.B(n_1328),
.C(n_1274),
.Y(n_1405)
);

INVx5_ASAP7_75t_L g1406 ( 
.A(n_1372),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1373),
.A2(n_1354),
.B(n_1364),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1285),
.A2(n_1333),
.B(n_1365),
.Y(n_1408)
);

BUFx4f_ASAP7_75t_SL g1409 ( 
.A(n_1398),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1368),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1277),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1277),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1376),
.Y(n_1413)
);

INVx5_ASAP7_75t_SL g1414 ( 
.A(n_1385),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1296),
.B(n_1289),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1288),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_L g1417 ( 
.A(n_1284),
.B(n_1282),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1349),
.A2(n_1372),
.B(n_1356),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1296),
.B(n_1291),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1337),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1298),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1391),
.A2(n_1294),
.B(n_1349),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.B(n_1287),
.Y(n_1423)
);

AO21x1_ASAP7_75t_L g1424 ( 
.A1(n_1281),
.A2(n_1343),
.B(n_1346),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1356),
.A2(n_1370),
.B(n_1366),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1287),
.B(n_1279),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1286),
.B(n_1320),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1307),
.B(n_1358),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1286),
.B(n_1291),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1319),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1345),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1316),
.B(n_1307),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1297),
.A2(n_1394),
.B1(n_1273),
.B2(n_1313),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1366),
.A2(n_1326),
.B(n_1365),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1395),
.A2(n_1400),
.B1(n_1389),
.B2(n_1278),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1326),
.A2(n_1352),
.B(n_1312),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1346),
.A2(n_1310),
.B(n_1308),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1312),
.A2(n_1300),
.B(n_1283),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1278),
.B(n_1389),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1283),
.B(n_1382),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1400),
.B(n_1299),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1303),
.A2(n_1330),
.B1(n_1322),
.B2(n_1321),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1272),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1371),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1300),
.B(n_1384),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1275),
.B(n_1304),
.Y(n_1446)
);

CKINVDCx8_ASAP7_75t_R g1447 ( 
.A(n_1386),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1374),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1390),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1324),
.A2(n_1342),
.B(n_1327),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1301),
.B(n_1306),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1290),
.B(n_1305),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1380),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1272),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1272),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1317),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1311),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1329),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1388),
.A2(n_1399),
.B1(n_1396),
.B2(n_1280),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1381),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1324),
.A2(n_1342),
.B(n_1362),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1275),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1304),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1377),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1314),
.B(n_1276),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1293),
.B(n_1315),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1363),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1302),
.B(n_1323),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1276),
.Y(n_1469)
);

INVx8_ASAP7_75t_L g1470 ( 
.A(n_1359),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1335),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_SL g1472 ( 
.A1(n_1325),
.A2(n_1347),
.B(n_1336),
.Y(n_1472)
);

NOR3xp33_ASAP7_75t_SL g1473 ( 
.A(n_1309),
.B(n_1338),
.C(n_1383),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1340),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1438),
.B(n_1422),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1461),
.B(n_1361),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1416),
.B(n_1378),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1405),
.A2(n_1347),
.B1(n_1325),
.B2(n_1344),
.C(n_1348),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1461),
.B(n_1348),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1434),
.A2(n_1418),
.B(n_1436),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1417),
.A2(n_1344),
.B(n_1361),
.C(n_1332),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1441),
.B(n_1361),
.Y(n_1482)
);

AO32x2_ASAP7_75t_L g1483 ( 
.A1(n_1442),
.A2(n_1424),
.A3(n_1455),
.B1(n_1443),
.B2(n_1462),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1417),
.A2(n_1398),
.B1(n_1397),
.B2(n_1379),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1435),
.A2(n_1309),
.B1(n_1295),
.B2(n_1292),
.Y(n_1485)
);

AO32x1_ASAP7_75t_L g1486 ( 
.A1(n_1448),
.A2(n_1350),
.A3(n_1360),
.B1(n_1332),
.B2(n_1336),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1469),
.B(n_1340),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1420),
.B(n_1341),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1441),
.B(n_1360),
.Y(n_1489)
);

AO22x2_ASAP7_75t_L g1490 ( 
.A1(n_1422),
.A2(n_1341),
.B1(n_1332),
.B2(n_1355),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1423),
.B(n_1331),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1433),
.B(n_1334),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1415),
.B(n_1383),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1438),
.B(n_1318),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1416),
.A2(n_1393),
.B1(n_1387),
.B2(n_1331),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1439),
.A2(n_1426),
.B(n_1438),
.C(n_1457),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1420),
.B(n_1437),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1439),
.A2(n_1442),
.B(n_1415),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1461),
.B(n_1427),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1469),
.B(n_1426),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1424),
.A2(n_1419),
.B1(n_1423),
.B2(n_1457),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1432),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1434),
.A2(n_1418),
.B(n_1425),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1471),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1451),
.B(n_1427),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1447),
.A2(n_1459),
.B1(n_1471),
.B2(n_1465),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1432),
.A2(n_1428),
.B(n_1451),
.C(n_1429),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_SL g1508 ( 
.A1(n_1472),
.A2(n_1449),
.B(n_1443),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1402),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1404),
.B(n_1429),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1440),
.B(n_1449),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1404),
.B(n_1437),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1404),
.A2(n_1416),
.B1(n_1403),
.B2(n_1408),
.Y(n_1513)
);

O2A1O1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1453),
.A2(n_1460),
.B(n_1404),
.C(n_1465),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1437),
.B(n_1401),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1401),
.A2(n_1446),
.B(n_1403),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1452),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1430),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1437),
.B(n_1401),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1430),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1401),
.B(n_1408),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1428),
.B(n_1449),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1444),
.B(n_1413),
.Y(n_1523)
);

NAND2xp33_ASAP7_75t_R g1524 ( 
.A(n_1473),
.B(n_1403),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1408),
.B(n_1444),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1408),
.B(n_1444),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1456),
.B(n_1452),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1447),
.A2(n_1409),
.B1(n_1474),
.B2(n_1414),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1445),
.B(n_1450),
.Y(n_1529)
);

NOR2x1_ASAP7_75t_R g1530 ( 
.A(n_1470),
.B(n_1468),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1456),
.B(n_1411),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1499),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1509),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1499),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1510),
.B(n_1411),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1498),
.A2(n_1464),
.B1(n_1463),
.B2(n_1466),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1495),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_L g1539 ( 
.A(n_1501),
.B(n_1403),
.C(n_1463),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1529),
.B(n_1407),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1523),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1412),
.Y(n_1542)
);

INVx4_ASAP7_75t_SL g1543 ( 
.A(n_1494),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1497),
.B(n_1412),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1525),
.B(n_1431),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1492),
.B(n_1468),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1520),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1522),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1488),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1531),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1505),
.B(n_1458),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1527),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1511),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1525),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1517),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1406),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1476),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1476),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1500),
.B(n_1467),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1526),
.B(n_1410),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1496),
.B(n_1502),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1479),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1559),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1544),
.Y(n_1567)
);

AOI211xp5_ASAP7_75t_L g1568 ( 
.A1(n_1564),
.A2(n_1506),
.B(n_1492),
.C(n_1496),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1559),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1539),
.A2(n_1501),
.B(n_1513),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1532),
.B(n_1521),
.Y(n_1571)
);

AOI221xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1545),
.A2(n_1507),
.B1(n_1513),
.B2(n_1514),
.C(n_1481),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1556),
.B(n_1526),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1546),
.Y(n_1574)
);

OAI321xp33_ASAP7_75t_L g1575 ( 
.A1(n_1537),
.A2(n_1475),
.A3(n_1512),
.B1(n_1507),
.B2(n_1485),
.C(n_1494),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1552),
.A2(n_1481),
.B(n_1530),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1557),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1546),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1547),
.Y(n_1580)
);

OAI31xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1549),
.A2(n_1528),
.A3(n_1478),
.B(n_1512),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1563),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1563),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1538),
.A2(n_1475),
.B1(n_1494),
.B2(n_1489),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1548),
.B(n_1475),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1547),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1548),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1536),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1550),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1559),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1556),
.B(n_1515),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1536),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1540),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1554),
.A2(n_1490),
.B1(n_1493),
.B2(n_1491),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1534),
.Y(n_1596)
);

AO221x1_ASAP7_75t_L g1597 ( 
.A1(n_1534),
.A2(n_1490),
.B1(n_1508),
.B2(n_1483),
.C(n_1454),
.Y(n_1597)
);

AO221x2_ASAP7_75t_L g1598 ( 
.A1(n_1565),
.A2(n_1483),
.B1(n_1524),
.B2(n_1490),
.C(n_1486),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1543),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1595),
.B(n_1487),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1594),
.B(n_1535),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1574),
.Y(n_1603)
);

OR2x2_ASAP7_75t_SL g1604 ( 
.A(n_1581),
.B(n_1503),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1578),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1574),
.Y(n_1606)
);

AND2x4_ASAP7_75t_SL g1607 ( 
.A(n_1599),
.B(n_1494),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1594),
.B(n_1560),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1592),
.B(n_1555),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1579),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1596),
.B(n_1555),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1580),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1596),
.B(n_1553),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1580),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1560),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1567),
.B(n_1553),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1586),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1576),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1589),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1578),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1599),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1566),
.B(n_1540),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1576),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1567),
.B(n_1542),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1582),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1573),
.B(n_1558),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1570),
.A2(n_1491),
.B1(n_1519),
.B2(n_1515),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1573),
.B(n_1558),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1582),
.B(n_1551),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1587),
.B(n_1588),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1561),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1603),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1632),
.B(n_1585),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1632),
.B(n_1585),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1568),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1630),
.A2(n_1570),
.B(n_1575),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1608),
.B(n_1566),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1608),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1568),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1566),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1604),
.B(n_1624),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1625),
.B(n_1566),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.B(n_1585),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1604),
.B(n_1477),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1572),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1602),
.B(n_1562),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1605),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1604),
.B(n_1624),
.Y(n_1656)
);

O2A1O1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1624),
.A2(n_1575),
.B(n_1482),
.C(n_1519),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1605),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1606),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1631),
.B(n_1587),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1610),
.B(n_1583),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1610),
.B(n_1583),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1606),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1541),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1615),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1626),
.B(n_1577),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1612),
.B(n_1588),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1611),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1615),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1621),
.B(n_1593),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1612),
.B(n_1593),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1611),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1613),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1621),
.B(n_1619),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1619),
.B(n_1578),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1626),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1677),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1667),
.B(n_1625),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1645),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1641),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1660),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1641),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1646),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1664),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1638),
.B(n_1599),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1667),
.B(n_1625),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1651),
.B(n_1628),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1642),
.B(n_1470),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1669),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1667),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1667),
.B(n_1625),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1640),
.B(n_1625),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1673),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1628),
.Y(n_1697)
);

OAI31xp67_ASAP7_75t_L g1698 ( 
.A1(n_1639),
.A2(n_1623),
.A3(n_1597),
.B(n_1483),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1649),
.B(n_1598),
.C(n_1484),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1675),
.B(n_1633),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1646),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1470),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1654),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1654),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1616),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1675),
.B(n_1633),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1616),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1650),
.B(n_1599),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1658),
.B(n_1613),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1644),
.B(n_1599),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_1633),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1643),
.B(n_1601),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1680),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1689),
.B(n_1636),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1680),
.Y(n_1716)
);

OAI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1699),
.A2(n_1656),
.B1(n_1644),
.B2(n_1671),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1681),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1681),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1678),
.B(n_1689),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1683),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1678),
.Y(n_1722)
);

AOI321xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1698),
.A2(n_1656),
.A3(n_1657),
.B1(n_1597),
.B2(n_1643),
.C(n_1648),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1699),
.A2(n_1597),
.B1(n_1672),
.B2(n_1668),
.C(n_1662),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1698),
.A2(n_1470),
.B(n_1598),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1683),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1686),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1697),
.A2(n_1584),
.B(n_1516),
.Y(n_1729)
);

OAI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1697),
.A2(n_1665),
.B1(n_1637),
.B2(n_1590),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1686),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1712),
.B(n_1655),
.Y(n_1732)
);

AOI322xp5_ASAP7_75t_L g1733 ( 
.A1(n_1705),
.A2(n_1627),
.A3(n_1584),
.B1(n_1601),
.B2(n_1647),
.C1(n_1634),
.C2(n_1617),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1712),
.B(n_1661),
.Y(n_1734)
);

NAND2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1687),
.B(n_1421),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1710),
.B(n_1659),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1653),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1691),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1722),
.B(n_1711),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1722),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1717),
.B(n_1711),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1720),
.B(n_1713),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1737),
.B(n_1702),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1724),
.A2(n_1708),
.B1(n_1692),
.B2(n_1710),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1720),
.B(n_1713),
.Y(n_1746)
);

OAI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1735),
.A2(n_1692),
.B1(n_1709),
.B2(n_1707),
.C(n_1705),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1725),
.A2(n_1729),
.B(n_1736),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1726),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1723),
.A2(n_1688),
.B1(n_1693),
.B2(n_1679),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1729),
.A2(n_1688),
.B1(n_1693),
.B2(n_1679),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1714),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1715),
.A2(n_1709),
.B1(n_1707),
.B2(n_1706),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1716),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1730),
.A2(n_1690),
.B1(n_1598),
.B2(n_1694),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1732),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1726),
.B(n_1694),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1718),
.B(n_1695),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1741),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1756),
.B(n_1719),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1745),
.A2(n_1700),
.B1(n_1706),
.B2(n_1734),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1749),
.B(n_1721),
.Y(n_1762)
);

XOR2x2_ASAP7_75t_L g1763 ( 
.A(n_1742),
.B(n_1470),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1740),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1758),
.Y(n_1765)
);

OAI31xp33_ASAP7_75t_L g1766 ( 
.A1(n_1748),
.A2(n_1739),
.A3(n_1738),
.B(n_1727),
.Y(n_1766)
);

AOI31xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1743),
.A2(n_1682),
.A3(n_1684),
.B(n_1733),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1753),
.B(n_1750),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1758),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1768),
.B(n_1747),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1757),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1766),
.B(n_1744),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1768),
.B(n_1746),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1759),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1762),
.B(n_1753),
.C(n_1755),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1763),
.A2(n_1751),
.B1(n_1754),
.B2(n_1752),
.Y(n_1776)
);

XOR2x2_ASAP7_75t_L g1777 ( 
.A(n_1760),
.B(n_1728),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1762),
.B(n_1731),
.Y(n_1778)
);

NOR3xp33_ASAP7_75t_L g1779 ( 
.A(n_1764),
.B(n_1684),
.C(n_1682),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1774),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1770),
.A2(n_1765),
.B(n_1769),
.C(n_1759),
.Y(n_1781)
);

OAI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1771),
.A2(n_1767),
.B(n_1684),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1775),
.A2(n_1773),
.B1(n_1772),
.B2(n_1778),
.C(n_1776),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1777),
.B(n_1695),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1780),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1782),
.B(n_1779),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1783),
.A2(n_1704),
.B1(n_1682),
.B2(n_1696),
.C(n_1701),
.Y(n_1787)
);

NOR3x1_ASAP7_75t_L g1788 ( 
.A(n_1781),
.B(n_1704),
.C(n_1696),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1784),
.B(n_1647),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1783),
.A2(n_1701),
.B1(n_1703),
.B2(n_1685),
.C(n_1659),
.Y(n_1790)
);

AO22x2_ASAP7_75t_L g1791 ( 
.A1(n_1786),
.A2(n_1703),
.B1(n_1685),
.B2(n_1676),
.Y(n_1791)
);

NAND4xp75_ASAP7_75t_L g1792 ( 
.A(n_1788),
.B(n_1703),
.C(n_1685),
.D(n_1609),
.Y(n_1792)
);

OR2x6_ASAP7_75t_L g1793 ( 
.A(n_1785),
.B(n_1789),
.Y(n_1793)
);

OR3x2_ASAP7_75t_L g1794 ( 
.A(n_1787),
.B(n_1414),
.C(n_1676),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1790),
.B(n_1634),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_L g1796 ( 
.A1(n_1793),
.A2(n_1607),
.B(n_1609),
.Y(n_1796)
);

NOR2xp67_ASAP7_75t_L g1797 ( 
.A(n_1795),
.B(n_1623),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1794),
.A2(n_1590),
.B(n_1569),
.C(n_1620),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1797),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1799),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1800),
.B(n_1796),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1800),
.A2(n_1792),
.B1(n_1794),
.B2(n_1798),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1801),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1802),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1804),
.A2(n_1791),
.B1(n_1414),
.B2(n_1607),
.Y(n_1806)
);

BUFx4_ASAP7_75t_R g1807 ( 
.A(n_1805),
.Y(n_1807)
);

AO21x2_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1806),
.B(n_1472),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1808),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1620),
.B1(n_1618),
.B2(n_1614),
.C(n_1622),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1618),
.B(n_1614),
.C(n_1622),
.Y(n_1811)
);


endmodule