module fake_jpeg_10337_n_47 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_47);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_32;

BUFx12_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_9),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_12),
.B1(n_14),
.B2(n_19),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_31),
.B1(n_42),
.B2(n_39),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_40),
.C(n_30),
.Y(n_45)
);

A2O1A1O1Ixp25_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_40),
.B(n_34),
.C(n_26),
.D(n_21),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_R g47 ( 
.A(n_46),
.B(n_28),
.Y(n_47)
);


endmodule