module fake_jpeg_28304_n_95 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_0),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_38),
.B(n_22),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_60),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_53),
.C(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_43),
.B1(n_46),
.B2(n_44),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_25),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_51),
.B1(n_50),
.B2(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_40),
.B1(n_47),
.B2(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_76),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_75),
.B1(n_70),
.B2(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_76),
.B1(n_72),
.B2(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_73),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_80),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_82),
.A3(n_83),
.B1(n_6),
.B2(n_7),
.C1(n_11),
.C2(n_12),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_5),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_29),
.B1(n_15),
.B2(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_84),
.B1(n_17),
.B2(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_33),
.C(n_24),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_28),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_31),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_32),
.C(n_35),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_36),
.C(n_7),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_69),
.Y(n_95)
);


endmodule