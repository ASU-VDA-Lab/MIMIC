module real_aes_11745_n_361 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_361);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_361;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1802;
wire n_727;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_729;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_0), .A2(n_161), .B1(n_570), .B2(n_904), .Y(n_1510) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_0), .A2(n_161), .B1(n_505), .B2(n_884), .Y(n_1517) );
INVxp67_ASAP7_75t_SL g1098 ( .A(n_1), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_1), .A2(n_8), .B1(n_514), .B2(n_889), .Y(n_1118) );
INVxp33_ASAP7_75t_L g754 ( .A(n_2), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_2), .A2(n_731), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g638 ( .A(n_3), .Y(n_638) );
INVx1_ASAP7_75t_L g1332 ( .A(n_4), .Y(n_1332) );
INVx1_ASAP7_75t_L g1459 ( .A(n_5), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_6), .A2(n_228), .B1(n_586), .B2(n_912), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_6), .A2(n_228), .B1(n_547), .B2(n_599), .Y(n_1126) );
INVx1_ASAP7_75t_L g1089 ( .A(n_7), .Y(n_1089) );
INVx1_ASAP7_75t_L g1097 ( .A(n_8), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_9), .A2(n_294), .B1(n_716), .B2(n_718), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_9), .A2(n_294), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g1595 ( .A(n_10), .Y(n_1595) );
INVxp33_ASAP7_75t_SL g450 ( .A(n_11), .Y(n_450) );
AOI22xp5_ASAP7_75t_SL g542 ( .A1(n_11), .A2(n_288), .B1(n_543), .B2(n_547), .Y(n_542) );
AO22x1_ASAP7_75t_L g391 ( .A1(n_12), .A2(n_392), .B1(n_393), .B2(n_555), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_12), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g1515 ( .A1(n_13), .A2(n_303), .B1(n_531), .B2(n_1045), .Y(n_1515) );
INVxp67_ASAP7_75t_L g1524 ( .A(n_13), .Y(n_1524) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_14), .A2(n_225), .B1(n_499), .B2(n_503), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_14), .A2(n_225), .B1(n_536), .B2(n_539), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_15), .A2(n_215), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_15), .A2(n_215), .B1(n_595), .B2(n_598), .Y(n_594) );
INVx1_ASAP7_75t_L g708 ( .A(n_16), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_16), .A2(n_60), .B1(n_722), .B2(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_17), .A2(n_244), .B1(n_886), .B2(n_915), .Y(n_996) );
AOI221xp5_ASAP7_75t_SL g1008 ( .A1(n_17), .A2(n_526), .B1(n_816), .B2(n_1009), .C(n_1010), .Y(n_1008) );
INVx1_ASAP7_75t_L g1088 ( .A(n_18), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_18), .A2(n_69), .B1(n_1103), .B2(n_1116), .Y(n_1119) );
INVx1_ASAP7_75t_L g571 ( .A(n_19), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_19), .A2(n_237), .B1(n_618), .B2(n_619), .Y(n_617) );
INVxp33_ASAP7_75t_SL g699 ( .A(n_20), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_20), .A2(n_103), .B1(n_426), .B2(n_661), .Y(n_744) );
AO221x2_ASAP7_75t_L g1593 ( .A1(n_21), .A2(n_263), .B1(n_1558), .B2(n_1577), .C(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1188 ( .A(n_22), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_22), .A2(n_323), .B1(n_860), .B2(n_862), .Y(n_1201) );
CKINVDCx16_ASAP7_75t_R g1570 ( .A(n_23), .Y(n_1570) );
INVx1_ASAP7_75t_L g1227 ( .A(n_24), .Y(n_1227) );
INVxp67_ASAP7_75t_SL g1472 ( .A(n_25), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_25), .A2(n_214), .B1(n_543), .B2(n_825), .Y(n_1492) );
OAI211xp5_ASAP7_75t_L g1418 ( .A1(n_26), .A2(n_712), .B(n_832), .C(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1437 ( .A(n_26), .Y(n_1437) );
INVx1_ASAP7_75t_L g1153 ( .A(n_27), .Y(n_1153) );
AOI22xp33_ASAP7_75t_SL g1166 ( .A1(n_27), .A2(n_200), .B1(n_531), .B2(n_1130), .Y(n_1166) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_28), .Y(n_1274) );
INVx1_ASAP7_75t_L g1502 ( .A(n_29), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_29), .A2(n_32), .B1(n_618), .B2(n_619), .Y(n_1521) );
AOI22xp33_ASAP7_75t_SL g1391 ( .A1(n_30), .A2(n_90), .B1(n_583), .B2(n_1392), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_30), .A2(n_90), .B1(n_825), .B2(n_836), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_31), .Y(n_1443) );
INVx1_ASAP7_75t_L g1503 ( .A(n_32), .Y(n_1503) );
INVx1_ASAP7_75t_L g1221 ( .A(n_33), .Y(n_1221) );
INVx1_ASAP7_75t_L g1064 ( .A(n_34), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_34), .A2(n_219), .B1(n_860), .B2(n_963), .Y(n_1069) );
INVx1_ASAP7_75t_L g695 ( .A(n_35), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_36), .A2(n_132), .B1(n_543), .B2(n_1037), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_36), .Y(n_1050) );
XNOR2xp5_ASAP7_75t_L g1830 ( .A(n_37), .B(n_1831), .Y(n_1830) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_38), .A2(n_350), .B1(n_608), .B2(n_609), .Y(n_607) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_38), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g966 ( .A1(n_39), .A2(n_486), .B(n_967), .C(n_969), .Y(n_966) );
INVx1_ASAP7_75t_L g1004 ( .A(n_39), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_40), .A2(n_116), .B1(n_455), .B2(n_720), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_40), .A2(n_116), .B1(n_543), .B2(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g367 ( .A(n_41), .Y(n_367) );
OAI211xp5_ASAP7_75t_L g1025 ( .A1(n_42), .A2(n_486), .B(n_1026), .C(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1043 ( .A(n_42), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_43), .A2(n_67), .B1(n_376), .B2(n_485), .Y(n_937) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_43), .A2(n_344), .B1(n_860), .B2(n_862), .Y(n_948) );
XNOR2xp5_ASAP7_75t_L g1324 ( .A(n_44), .B(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g429 ( .A(n_45), .Y(n_429) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_46), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_46), .A2(n_193), .B1(n_790), .B2(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g1505 ( .A(n_47), .Y(n_1505) );
INVxp67_ASAP7_75t_L g1805 ( .A(n_48), .Y(n_1805) );
AOI22xp33_ASAP7_75t_L g1819 ( .A1(n_48), .A2(n_276), .B1(n_825), .B2(n_1820), .Y(n_1819) );
INVxp67_ASAP7_75t_SL g1796 ( .A(n_49), .Y(n_1796) );
OAI22xp5_ASAP7_75t_L g1802 ( .A1(n_49), .A2(n_360), .B1(n_618), .B2(n_1105), .Y(n_1802) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_50), .A2(n_187), .B1(n_517), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_50), .A2(n_187), .B1(n_426), .B2(n_601), .Y(n_600) );
INVxp33_ASAP7_75t_L g1388 ( .A(n_51), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_51), .A2(n_290), .B1(n_895), .B2(n_1257), .Y(n_1408) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_52), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_52), .A2(n_287), .B1(n_716), .B2(n_725), .Y(n_724) );
INVxp33_ASAP7_75t_SL g482 ( .A(n_53), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_53), .A2(n_285), .B1(n_536), .B2(n_550), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_54), .A2(n_340), .B1(n_860), .B2(n_963), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_54), .A2(n_242), .B1(n_677), .B2(n_1291), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_55), .A2(n_312), .B1(n_912), .B2(n_913), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_55), .A2(n_312), .B1(n_597), .B2(n_923), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_56), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_57), .A2(n_196), .B1(n_915), .B2(n_1103), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_57), .A2(n_196), .B1(n_570), .B2(n_904), .Y(n_1162) );
INVxp33_ASAP7_75t_SL g1460 ( .A(n_58), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_58), .A2(n_199), .B1(n_790), .B2(n_889), .Y(n_1477) );
INVxp33_ASAP7_75t_SL g1474 ( .A(n_59), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_59), .A2(n_74), .B1(n_606), .B2(n_1488), .Y(n_1491) );
INVxp33_ASAP7_75t_SL g703 ( .A(n_60), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_61), .A2(n_85), .B1(n_866), .B2(n_870), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_61), .A2(n_85), .B1(n_597), .B2(n_598), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g1576 ( .A1(n_62), .A2(n_325), .B1(n_1558), .B2(n_1577), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g1809 ( .A1(n_63), .A2(n_65), .B1(n_1402), .B2(n_1810), .Y(n_1809) );
AOI22xp33_ASAP7_75t_L g1815 ( .A1(n_63), .A2(n_65), .B1(n_737), .B2(n_1345), .Y(n_1815) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_64), .A2(n_111), .B1(n_866), .B2(n_870), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_64), .A2(n_101), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_66), .A2(n_355), .B1(n_866), .B2(n_870), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_66), .A2(n_355), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_67), .A2(n_182), .B1(n_709), .B2(n_928), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_68), .A2(n_139), .B1(n_376), .B2(n_485), .Y(n_972) );
INVx1_ASAP7_75t_L g1001 ( .A(n_68), .Y(n_1001) );
INVx1_ASAP7_75t_L g1092 ( .A(n_69), .Y(n_1092) );
INVx1_ASAP7_75t_L g1101 ( .A(n_70), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_70), .A2(n_246), .B1(n_541), .B2(n_895), .Y(n_1128) );
INVx1_ASAP7_75t_L g641 ( .A(n_71), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_72), .A2(n_952), .B1(n_1018), .B2(n_1019), .Y(n_951) );
INVxp67_ASAP7_75t_SL g1019 ( .A(n_72), .Y(n_1019) );
INVx1_ASAP7_75t_L g635 ( .A(n_73), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_73), .A2(n_162), .B1(n_543), .B2(n_648), .Y(n_663) );
INVxp67_ASAP7_75t_SL g1468 ( .A(n_74), .Y(n_1468) );
AOI22xp33_ASAP7_75t_L g1808 ( .A1(n_75), .A2(n_142), .B1(n_677), .B2(n_1439), .Y(n_1808) );
AOI22xp33_ASAP7_75t_L g1816 ( .A1(n_75), .A2(n_142), .B1(n_598), .B2(n_826), .Y(n_1816) );
INVx1_ASAP7_75t_L g1219 ( .A(n_76), .Y(n_1219) );
INVx1_ASAP7_75t_L g935 ( .A(n_77), .Y(n_935) );
AO22x2_ASAP7_75t_L g1267 ( .A1(n_78), .A2(n_1268), .B1(n_1269), .B2(n_1319), .Y(n_1267) );
INVxp67_ASAP7_75t_L g1319 ( .A(n_78), .Y(n_1319) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_79), .Y(n_1205) );
INVxp33_ASAP7_75t_SL g650 ( .A(n_80), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_80), .A2(n_154), .B1(n_507), .B2(n_674), .Y(n_679) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_81), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_81), .A2(n_266), .B1(n_825), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g425 ( .A(n_82), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_82), .A2(n_118), .B1(n_499), .B2(n_517), .Y(n_516) );
INVxp67_ASAP7_75t_SL g992 ( .A(n_83), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_83), .A2(n_97), .B1(n_1013), .B2(n_1016), .Y(n_1012) );
INVx1_ASAP7_75t_L g1034 ( .A(n_84), .Y(n_1034) );
AOI221xp5_ASAP7_75t_L g1438 ( .A1(n_86), .A2(n_252), .B1(n_1439), .B2(n_1440), .C(n_1441), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_86), .A2(n_252), .B1(n_1130), .B2(n_1235), .Y(n_1446) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_87), .A2(n_95), .B1(n_892), .B2(n_1484), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_87), .A2(n_95), .B1(n_606), .B2(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g415 ( .A(n_88), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_89), .A2(n_239), .B1(n_866), .B2(n_870), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_89), .A2(n_239), .B1(n_599), .B2(n_1235), .Y(n_1449) );
BUFx2_ASAP7_75t_L g447 ( .A(n_91), .Y(n_447) );
BUFx2_ASAP7_75t_L g491 ( .A(n_91), .Y(n_491) );
INVx1_ASAP7_75t_L g521 ( .A(n_91), .Y(n_521) );
INVx1_ASAP7_75t_L g568 ( .A(n_92), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_92), .A2(n_194), .B1(n_579), .B2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g1338 ( .A1(n_93), .A2(n_233), .B1(n_467), .B2(n_579), .Y(n_1338) );
AOI22xp33_ASAP7_75t_SL g1344 ( .A1(n_93), .A2(n_233), .B1(n_426), .B2(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1462 ( .A(n_94), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1478 ( .A1(n_94), .A2(n_114), .B1(n_886), .B2(n_1116), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_96), .A2(n_322), .B1(n_886), .B2(n_915), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_96), .A2(n_322), .B1(n_570), .B2(n_666), .Y(n_921) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_97), .Y(n_995) );
INVx1_ASAP7_75t_L g1139 ( .A(n_98), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_98), .A2(n_354), .B1(n_509), .B2(n_586), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1480 ( .A1(n_99), .A2(n_273), .B1(n_889), .B2(n_1481), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_99), .A2(n_273), .B1(n_534), .B2(n_1006), .Y(n_1489) );
XNOR2xp5_ASAP7_75t_L g846 ( .A(n_100), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g1278 ( .A(n_101), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g1428 ( .A(n_102), .Y(n_1428) );
INVx1_ASAP7_75t_L g694 ( .A(n_103), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_104), .A2(n_352), .B1(n_666), .B2(n_709), .Y(n_1514) );
INVxp33_ASAP7_75t_L g1526 ( .A(n_104), .Y(n_1526) );
INVx1_ASAP7_75t_L g1258 ( .A(n_105), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_106), .A2(n_107), .B1(n_866), .B2(n_870), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_106), .A2(n_107), .B1(n_597), .B2(n_1045), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_108), .A2(n_117), .B1(n_1095), .B2(n_1144), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_108), .A2(n_117), .B1(n_876), .B2(n_1105), .Y(n_1148) );
INVx1_ASAP7_75t_L g436 ( .A(n_109), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g1572 ( .A(n_110), .Y(n_1572) );
INVx1_ASAP7_75t_L g1314 ( .A(n_111), .Y(n_1314) );
INVx1_ASAP7_75t_L g949 ( .A(n_112), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_113), .A2(n_137), .B1(n_660), .B2(n_662), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_113), .A2(n_137), .B1(n_636), .B2(n_674), .Y(n_673) );
INVxp33_ASAP7_75t_SL g1456 ( .A(n_114), .Y(n_1456) );
INVx1_ASAP7_75t_L g1251 ( .A(n_115), .Y(n_1251) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_118), .Y(n_396) );
INVxp33_ASAP7_75t_SL g632 ( .A(n_119), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_119), .A2(n_164), .B1(n_657), .B2(n_665), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_120), .Y(n_1442) );
INVx1_ASAP7_75t_L g1231 ( .A(n_121), .Y(n_1231) );
OAI22xp33_ASAP7_75t_SL g1264 ( .A1(n_121), .A2(n_216), .B1(n_376), .B2(n_866), .Y(n_1264) );
AO22x2_ASAP7_75t_L g1494 ( .A1(n_122), .A2(n_1495), .B1(n_1527), .B2(n_1528), .Y(n_1494) );
INVx1_ASAP7_75t_L g1527 ( .A(n_122), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_123), .A2(n_224), .B1(n_608), .B2(n_1354), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_123), .A2(n_224), .B1(n_866), .B2(n_870), .Y(n_1362) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_124), .A2(n_319), .B1(n_1558), .B2(n_1577), .Y(n_1592) );
INVxp33_ASAP7_75t_SL g1384 ( .A(n_125), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_125), .A2(n_217), .B1(n_1410), .B2(n_1411), .Y(n_1409) );
INVxp67_ASAP7_75t_SL g1799 ( .A(n_126), .Y(n_1799) );
AOI22xp33_ASAP7_75t_L g1818 ( .A1(n_126), .A2(n_301), .B1(n_737), .B2(n_895), .Y(n_1818) );
XOR2xp5_ASAP7_75t_L g1168 ( .A(n_127), .B(n_1169), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_128), .A2(n_309), .B1(n_1130), .B2(n_1235), .Y(n_1509) );
AOI22xp33_ASAP7_75t_SL g1516 ( .A1(n_128), .A2(n_309), .B1(n_586), .B2(n_912), .Y(n_1516) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_129), .A2(n_242), .B1(n_862), .B2(n_955), .Y(n_1328) );
INVxp33_ASAP7_75t_SL g1361 ( .A(n_129), .Y(n_1361) );
AOI22xp33_ASAP7_75t_SL g1393 ( .A1(n_130), .A2(n_298), .B1(n_730), .B2(n_1394), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_130), .A2(n_298), .B1(n_734), .B2(n_1257), .Y(n_1405) );
INVxp33_ASAP7_75t_SL g1371 ( .A(n_131), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_131), .A2(n_341), .B1(n_1397), .B2(n_1399), .Y(n_1396) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_132), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1539 ( .A1(n_133), .A2(n_136), .B1(n_1540), .B2(n_1548), .Y(n_1539) );
INVxp67_ASAP7_75t_SL g1501 ( .A(n_134), .Y(n_1501) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_134), .A2(n_212), .B1(n_505), .B2(n_915), .Y(n_1512) );
INVx1_ASAP7_75t_L g1247 ( .A(n_135), .Y(n_1247) );
OAI22xp33_ASAP7_75t_L g1253 ( .A1(n_135), .A2(n_143), .B1(n_860), .B2(n_963), .Y(n_1253) );
XNOR2xp5_ASAP7_75t_L g1783 ( .A(n_136), .B(n_1784), .Y(n_1783) );
AOI22xp5_ASAP7_75t_L g1828 ( .A1(n_136), .A2(n_1829), .B1(n_1832), .B2(n_1835), .Y(n_1828) );
AOI22xp5_ASAP7_75t_L g1551 ( .A1(n_138), .A2(n_338), .B1(n_1552), .B2(n_1556), .Y(n_1551) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_139), .A2(n_345), .B1(n_862), .B2(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g1185 ( .A(n_140), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_140), .A2(n_291), .B1(n_955), .B2(n_963), .Y(n_1207) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_141), .A2(n_688), .B1(n_748), .B2(n_749), .Y(n_687) );
INVxp67_ASAP7_75t_L g748 ( .A(n_141), .Y(n_748) );
INVx1_ASAP7_75t_L g1250 ( .A(n_143), .Y(n_1250) );
INVxp33_ASAP7_75t_SL g1499 ( .A(n_144), .Y(n_1499) );
AOI22xp33_ASAP7_75t_SL g1511 ( .A1(n_144), .A2(n_316), .B1(n_586), .B2(n_912), .Y(n_1511) );
AO221x2_ASAP7_75t_L g1612 ( .A1(n_145), .A2(n_209), .B1(n_1552), .B2(n_1558), .C(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1544 ( .A(n_146), .Y(n_1544) );
OAI211xp5_ASAP7_75t_L g871 ( .A1(n_147), .A2(n_486), .B(n_872), .C(n_874), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_147), .A2(n_251), .B1(n_896), .B2(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g1668 ( .A(n_148), .Y(n_1668) );
CKINVDCx5p33_ASAP7_75t_R g1137 ( .A(n_149), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_150), .A2(n_357), .B1(n_376), .B2(n_485), .Y(n_1024) );
INVx1_ASAP7_75t_L g1040 ( .A(n_150), .Y(n_1040) );
XOR2x2_ASAP7_75t_L g557 ( .A(n_151), .B(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_152), .A2(n_226), .B1(n_791), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_152), .A2(n_226), .B1(n_597), .B2(n_598), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_153), .A2(n_238), .B1(n_614), .B2(n_1116), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_153), .A2(n_238), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_154), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g750 ( .A(n_155), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g1575 ( .A1(n_155), .A2(n_353), .B1(n_1540), .B2(n_1548), .Y(n_1575) );
INVx1_ASAP7_75t_L g1377 ( .A(n_156), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_156), .A2(n_282), .B1(n_619), .B2(n_971), .Y(n_1382) );
OAI211xp5_ASAP7_75t_L g1282 ( .A1(n_157), .A2(n_712), .B(n_1002), .C(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1303 ( .A(n_157), .Y(n_1303) );
INVx1_ASAP7_75t_L g1197 ( .A(n_158), .Y(n_1197) );
OAI22xp33_ASAP7_75t_SL g1212 ( .A1(n_158), .A2(n_169), .B1(n_376), .B2(n_866), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_159), .A2(n_295), .B1(n_507), .B2(n_510), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_159), .A2(n_295), .B1(n_530), .B2(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g1545 ( .A(n_160), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1550 ( .A(n_160), .B(n_1543), .Y(n_1550) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_162), .Y(n_633) );
INVxp33_ASAP7_75t_SL g408 ( .A(n_163), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_163), .A2(n_234), .B1(n_507), .B2(n_514), .Y(n_513) );
INVxp33_ASAP7_75t_SL g640 ( .A(n_164), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g1416 ( .A1(n_165), .A2(n_176), .B1(n_860), .B2(n_963), .Y(n_1416) );
AOI221xp5_ASAP7_75t_L g1432 ( .A1(n_165), .A2(n_306), .B1(n_507), .B2(n_1433), .C(n_1435), .Y(n_1432) );
INVxp67_ASAP7_75t_SL g1791 ( .A(n_166), .Y(n_1791) );
AOI22xp33_ASAP7_75t_SL g1812 ( .A1(n_166), .A2(n_221), .B1(n_718), .B2(n_1439), .Y(n_1812) );
INVx2_ASAP7_75t_L g379 ( .A(n_167), .Y(n_379) );
INVxp33_ASAP7_75t_L g1370 ( .A(n_168), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_168), .A2(n_330), .B1(n_505), .B2(n_1402), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_169), .A2(n_281), .B1(n_597), .B2(n_599), .Y(n_1199) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_170), .A2(n_307), .B1(n_604), .B2(n_606), .Y(n_603) );
INVxp33_ASAP7_75t_SL g624 ( .A(n_170), .Y(n_624) );
INVx1_ASAP7_75t_L g1059 ( .A(n_171), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1074 ( .A1(n_171), .A2(n_357), .B1(n_862), .B2(n_955), .Y(n_1074) );
BUFx3_ASAP7_75t_L g405 ( .A(n_172), .Y(n_405) );
INVx1_ASAP7_75t_L g423 ( .A(n_172), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_173), .A2(n_179), .B1(n_426), .B2(n_601), .Y(n_1352) );
INVx1_ASAP7_75t_L g1360 ( .A(n_173), .Y(n_1360) );
INVx1_ASAP7_75t_L g760 ( .A(n_174), .Y(n_760) );
INVx1_ASAP7_75t_L g1614 ( .A(n_175), .Y(n_1614) );
INVx1_ASAP7_75t_L g1436 ( .A(n_176), .Y(n_1436) );
AOI22xp33_ASAP7_75t_SL g1156 ( .A1(n_177), .A2(n_231), .B1(n_586), .B2(n_912), .Y(n_1156) );
AOI22xp33_ASAP7_75t_SL g1163 ( .A1(n_177), .A2(n_231), .B1(n_531), .B2(n_599), .Y(n_1163) );
INVx1_ASAP7_75t_L g757 ( .A(n_178), .Y(n_757) );
INVx1_ASAP7_75t_L g1358 ( .A(n_179), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_180), .A2(n_336), .B1(n_860), .B2(n_963), .Y(n_1286) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_180), .A2(n_336), .B1(n_507), .B2(n_674), .C(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1136 ( .A(n_181), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_181), .A2(n_308), .B1(n_915), .B2(n_1103), .Y(n_1160) );
OAI211xp5_ASAP7_75t_SL g931 ( .A1(n_182), .A2(n_486), .B(n_932), .C(n_934), .Y(n_931) );
INVxp33_ASAP7_75t_L g755 ( .A(n_183), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_183), .A2(n_299), .B1(n_790), .B2(n_791), .C(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g1666 ( .A(n_184), .Y(n_1666) );
INVx1_ASAP7_75t_L g1066 ( .A(n_185), .Y(n_1066) );
OAI211xp5_ASAP7_75t_L g1070 ( .A1(n_185), .A2(n_712), .B(n_1071), .C(n_1073), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_186), .A2(n_324), .B1(n_1291), .B2(n_1336), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_186), .A2(n_324), .B1(n_609), .B2(n_1348), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_188), .A2(n_344), .B1(n_884), .B2(n_886), .Y(n_919) );
INVx1_ASAP7_75t_L g941 ( .A(n_188), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_189), .A2(n_284), .B1(n_543), .B2(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_189), .A2(n_284), .B1(n_507), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g1793 ( .A(n_190), .Y(n_1793) );
AOI22xp33_ASAP7_75t_L g1813 ( .A1(n_190), .A2(n_198), .B1(n_467), .B2(n_1402), .Y(n_1813) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_191), .A2(n_1022), .B1(n_1075), .B2(n_1076), .Y(n_1021) );
INVx1_ASAP7_75t_L g1076 ( .A(n_191), .Y(n_1076) );
INVx1_ASAP7_75t_L g855 ( .A(n_192), .Y(n_855) );
INVx1_ASAP7_75t_L g858 ( .A(n_193), .Y(n_858) );
INVxp33_ASAP7_75t_SL g561 ( .A(n_194), .Y(n_561) );
XNOR2xp5_ASAP7_75t_L g1413 ( .A(n_195), .B(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1615 ( .A(n_195), .Y(n_1615) );
INVx1_ASAP7_75t_L g1232 ( .A(n_197), .Y(n_1232) );
OAI211xp5_ASAP7_75t_SL g1262 ( .A1(n_197), .A2(n_486), .B(n_872), .C(n_1263), .Y(n_1262) );
INVxp33_ASAP7_75t_SL g1787 ( .A(n_198), .Y(n_1787) );
INVxp33_ASAP7_75t_SL g1457 ( .A(n_199), .Y(n_1457) );
INVx1_ASAP7_75t_L g1151 ( .A(n_200), .Y(n_1151) );
INVx1_ASAP7_75t_L g445 ( .A(n_201), .Y(n_445) );
INVx1_ASAP7_75t_L g936 ( .A(n_202), .Y(n_936) );
INVx1_ASAP7_75t_L g1035 ( .A(n_203), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_204), .A2(n_206), .B1(n_580), .B2(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_204), .A2(n_206), .B1(n_734), .B2(n_737), .Y(n_733) );
INVxp67_ASAP7_75t_L g1110 ( .A(n_205), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_205), .A2(n_293), .B1(n_531), .B2(n_1130), .Y(n_1129) );
INVxp67_ASAP7_75t_SL g1180 ( .A(n_207), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_207), .A2(n_329), .B1(n_599), .B2(n_658), .Y(n_1194) );
INVx1_ASAP7_75t_L g1587 ( .A(n_208), .Y(n_1587) );
INVx1_ASAP7_75t_L g565 ( .A(n_210), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g1591 ( .A1(n_211), .A2(n_296), .B1(n_1540), .B2(n_1548), .Y(n_1591) );
INVxp33_ASAP7_75t_SL g1498 ( .A(n_212), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_213), .A2(n_302), .B1(n_534), .B2(n_658), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_213), .A2(n_302), .B1(n_866), .B2(n_870), .Y(n_930) );
INVxp33_ASAP7_75t_L g1471 ( .A(n_214), .Y(n_1471) );
INVx1_ASAP7_75t_L g1236 ( .A(n_216), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1386 ( .A(n_217), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_218), .A2(n_306), .B1(n_862), .B2(n_955), .Y(n_1417) );
INVx1_ASAP7_75t_L g1429 ( .A(n_218), .Y(n_1429) );
INVx1_ASAP7_75t_L g1057 ( .A(n_219), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g1293 ( .A(n_220), .Y(n_1293) );
INVxp33_ASAP7_75t_SL g1788 ( .A(n_221), .Y(n_1788) );
INVx1_ASAP7_75t_L g1176 ( .A(n_222), .Y(n_1176) );
INVx1_ASAP7_75t_L g854 ( .A(n_223), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_227), .A2(n_304), .B1(n_860), .B2(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g983 ( .A(n_227), .Y(n_983) );
CKINVDCx16_ASAP7_75t_R g1584 ( .A(n_229), .Y(n_1584) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_230), .A2(n_258), .B1(n_884), .B2(n_886), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_230), .A2(n_258), .B1(n_895), .B2(n_896), .Y(n_894) );
INVx1_ASAP7_75t_L g961 ( .A(n_232), .Y(n_961) );
INVxp33_ASAP7_75t_SL g419 ( .A(n_234), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g1285 ( .A1(n_235), .A2(n_241), .B1(n_862), .B2(n_955), .Y(n_1285) );
INVx1_ASAP7_75t_L g1301 ( .A(n_235), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_236), .A2(n_268), .B1(n_912), .B2(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g947 ( .A(n_236), .Y(n_947) );
INVx1_ASAP7_75t_L g573 ( .A(n_237), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_240), .Y(n_787) );
INVx1_ASAP7_75t_L g1279 ( .A(n_241), .Y(n_1279) );
INVx1_ASAP7_75t_L g647 ( .A(n_243), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_243), .A2(n_292), .B1(n_505), .B2(n_588), .Y(n_680) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_244), .Y(n_1011) );
INVx1_ASAP7_75t_L g1238 ( .A(n_245), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_245), .A2(n_253), .B1(n_485), .B2(n_870), .Y(n_1261) );
INVxp33_ASAP7_75t_L g1107 ( .A(n_246), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_247), .Y(n_1425) );
INVx1_ASAP7_75t_L g637 ( .A(n_248), .Y(n_637) );
BUFx3_ASAP7_75t_L g407 ( .A(n_249), .Y(n_407) );
INVx1_ASAP7_75t_L g413 ( .A(n_249), .Y(n_413) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_250), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_250), .A2(n_257), .B1(n_507), .B2(n_588), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_251), .A2(n_328), .B1(n_376), .B2(n_485), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g1254 ( .A1(n_253), .A2(n_261), .B1(n_862), .B2(n_955), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_254), .Y(n_375) );
INVx1_ASAP7_75t_L g523 ( .A(n_254), .Y(n_523) );
AND2x2_ASAP7_75t_L g767 ( .A(n_254), .B(n_454), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_254), .B(n_334), .Y(n_781) );
INVx1_ASAP7_75t_L g762 ( .A(n_255), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g774 ( .A1(n_255), .A2(n_358), .B1(n_775), .B2(n_782), .C(n_784), .Y(n_774) );
AOI221xp5_ASAP7_75t_SL g1289 ( .A1(n_256), .A2(n_270), .B1(n_677), .B2(n_1290), .C(n_1292), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_256), .A2(n_270), .B1(n_598), .B2(n_1310), .Y(n_1309) );
INVxp33_ASAP7_75t_SL g563 ( .A(n_257), .Y(n_563) );
INVx1_ASAP7_75t_L g1672 ( .A(n_259), .Y(n_1672) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_260), .Y(n_1206) );
INVx1_ASAP7_75t_L g1248 ( .A(n_261), .Y(n_1248) );
INVx1_ASAP7_75t_L g960 ( .A(n_262), .Y(n_960) );
XNOR2xp5_ASAP7_75t_L g1213 ( .A(n_264), .B(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1588 ( .A(n_264), .Y(n_1588) );
INVx2_ASAP7_75t_L g400 ( .A(n_265), .Y(n_400) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_266), .Y(n_768) );
INVx1_ASAP7_75t_L g1084 ( .A(n_267), .Y(n_1084) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_268), .Y(n_946) );
INVx1_ASAP7_75t_L g1670 ( .A(n_269), .Y(n_1670) );
INVx1_ASAP7_75t_L g1373 ( .A(n_271), .Y(n_1373) );
INVx1_ASAP7_75t_L g1464 ( .A(n_272), .Y(n_1464) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_272), .A2(n_315), .B1(n_618), .B2(n_1105), .Y(n_1469) );
INVxp33_ASAP7_75t_SL g691 ( .A(n_274), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_274), .A2(n_279), .B1(n_746), .B2(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g1259 ( .A(n_275), .Y(n_1259) );
INVxp67_ASAP7_75t_L g1804 ( .A(n_276), .Y(n_1804) );
CKINVDCx16_ASAP7_75t_R g1585 ( .A(n_277), .Y(n_1585) );
OAI211xp5_ASAP7_75t_L g956 ( .A1(n_278), .A2(n_712), .B(n_957), .C(n_959), .Y(n_956) );
INVx1_ASAP7_75t_L g985 ( .A(n_278), .Y(n_985) );
INVxp33_ASAP7_75t_SL g692 ( .A(n_279), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g1329 ( .A1(n_280), .A2(n_712), .B(n_833), .C(n_1330), .Y(n_1329) );
AOI22xp33_ASAP7_75t_SL g1342 ( .A1(n_280), .A2(n_340), .B1(n_467), .B2(n_580), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_281), .A2(n_323), .B1(n_485), .B2(n_870), .Y(n_1209) );
INVx1_ASAP7_75t_L g1378 ( .A(n_282), .Y(n_1378) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_283), .Y(n_1296) );
INVx1_ASAP7_75t_L g466 ( .A(n_285), .Y(n_466) );
INVx1_ASAP7_75t_L g1563 ( .A(n_286), .Y(n_1563) );
INVxp33_ASAP7_75t_SL g704 ( .A(n_287), .Y(n_704) );
INVxp33_ASAP7_75t_SL g459 ( .A(n_288), .Y(n_459) );
INVx1_ASAP7_75t_L g1790 ( .A(n_289), .Y(n_1790) );
INVxp67_ASAP7_75t_SL g1381 ( .A(n_290), .Y(n_1381) );
INVx1_ASAP7_75t_L g1183 ( .A(n_291), .Y(n_1183) );
INVxp33_ASAP7_75t_SL g645 ( .A(n_292), .Y(n_645) );
INVx1_ASAP7_75t_L g1108 ( .A(n_293), .Y(n_1108) );
INVx1_ASAP7_75t_L g1198 ( .A(n_297), .Y(n_1198) );
OAI211xp5_ASAP7_75t_SL g1210 ( .A1(n_297), .A2(n_486), .B(n_872), .C(n_1211), .Y(n_1210) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_299), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_300), .A2(n_332), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_300), .A2(n_332), .B1(n_618), .B2(n_1105), .Y(n_1104) );
INVxp67_ASAP7_75t_SL g1801 ( .A(n_301), .Y(n_1801) );
INVxp33_ASAP7_75t_L g1523 ( .A(n_303), .Y(n_1523) );
INVx1_ASAP7_75t_L g976 ( .A(n_304), .Y(n_976) );
INVx1_ASAP7_75t_L g1150 ( .A(n_305), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_305), .A2(n_337), .B1(n_541), .B2(n_904), .Y(n_1165) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_307), .Y(n_616) );
INVx1_ASAP7_75t_L g1142 ( .A(n_308), .Y(n_1142) );
INVx1_ASAP7_75t_L g1596 ( .A(n_310), .Y(n_1596) );
INVx1_ASAP7_75t_L g696 ( .A(n_311), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_313), .A2(n_328), .B1(n_860), .B2(n_862), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_313), .A2(n_343), .B1(n_891), .B2(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g1224 ( .A(n_314), .Y(n_1224) );
INVx1_ASAP7_75t_L g1463 ( .A(n_315), .Y(n_1463) );
INVxp33_ASAP7_75t_SL g1506 ( .A(n_316), .Y(n_1506) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_317), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_317), .B(n_367), .Y(n_1547) );
AND3x2_ASAP7_75t_L g1555 ( .A(n_317), .B(n_367), .C(n_1544), .Y(n_1555) );
INVx2_ASAP7_75t_L g380 ( .A(n_318), .Y(n_380) );
INVx1_ASAP7_75t_L g1029 ( .A(n_320), .Y(n_1029) );
AOI21xp33_ASAP7_75t_L g785 ( .A1(n_321), .A2(n_469), .B(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_321), .Y(n_823) );
INVx1_ASAP7_75t_L g806 ( .A(n_326), .Y(n_806) );
INVx1_ASAP7_75t_L g700 ( .A(n_327), .Y(n_700) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_329), .Y(n_1178) );
INVxp67_ASAP7_75t_SL g1376 ( .A(n_330), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1420 ( .A(n_331), .Y(n_1420) );
INVx1_ASAP7_75t_L g1173 ( .A(n_333), .Y(n_1173) );
INVx1_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
INVx2_ASAP7_75t_L g454 ( .A(n_334), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g1132 ( .A(n_335), .B(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1147 ( .A(n_337), .Y(n_1147) );
INVx1_ASAP7_75t_L g803 ( .A(n_339), .Y(n_803) );
INVxp33_ASAP7_75t_L g1374 ( .A(n_341), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_342), .Y(n_1276) );
INVx1_ASAP7_75t_L g851 ( .A(n_343), .Y(n_851) );
INVx1_ASAP7_75t_L g980 ( .A(n_345), .Y(n_980) );
CKINVDCx5p33_ASAP7_75t_R g1421 ( .A(n_346), .Y(n_1421) );
AO22x2_ASAP7_75t_L g627 ( .A1(n_347), .A2(n_628), .B1(n_629), .B2(n_684), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_347), .Y(n_628) );
INVx1_ASAP7_75t_L g1028 ( .A(n_348), .Y(n_1028) );
INVx1_ASAP7_75t_L g1331 ( .A(n_349), .Y(n_1331) );
INVxp33_ASAP7_75t_SL g621 ( .A(n_350), .Y(n_621) );
XOR2x2_ASAP7_75t_L g1452 ( .A(n_351), .B(n_1453), .Y(n_1452) );
INVxp67_ASAP7_75t_SL g1520 ( .A(n_352), .Y(n_1520) );
INVx1_ASAP7_75t_L g1140 ( .A(n_354), .Y(n_1140) );
INVx1_ASAP7_75t_L g1189 ( .A(n_356), .Y(n_1189) );
INVx1_ASAP7_75t_L g761 ( .A(n_358), .Y(n_761) );
AO22x1_ASAP7_75t_L g1365 ( .A1(n_359), .A2(n_1366), .B1(n_1367), .B2(n_1412), .Y(n_1365) );
INVxp67_ASAP7_75t_L g1366 ( .A(n_359), .Y(n_1366) );
INVxp67_ASAP7_75t_SL g1795 ( .A(n_360), .Y(n_1795) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_383), .B(n_1531), .Y(n_361) );
INVx3_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_370), .Y(n_364) );
AND2x4_ASAP7_75t_L g1827 ( .A(n_365), .B(n_371), .Y(n_1827) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_SL g1834 ( .A(n_366), .Y(n_1834) );
NAND2xp5_ASAP7_75t_L g1838 ( .A(n_366), .B(n_368), .Y(n_1838) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g1833 ( .A(n_368), .B(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_376), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x6_ASAP7_75t_L g490 ( .A(n_373), .B(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_373), .B(n_491), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g497 ( .A(n_374), .B(n_382), .Y(n_497) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g998 ( .A(n_375), .B(n_453), .Y(n_998) );
INVx8_ASAP7_75t_L g483 ( .A(n_376), .Y(n_483) );
OR2x6_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
OR2x6_ASAP7_75t_L g485 ( .A(n_377), .B(n_452), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_377), .A2(n_497), .B(n_787), .Y(n_786) );
BUFx6f_ASAP7_75t_L g984 ( .A(n_377), .Y(n_984) );
INVx1_ASAP7_75t_L g1063 ( .A(n_377), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1187 ( .A(n_377), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_377), .Y(n_1243) );
INVx2_ASAP7_75t_SL g1295 ( .A(n_377), .Y(n_1295) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g456 ( .A(n_379), .Y(n_456) );
AND2x4_ASAP7_75t_L g463 ( .A(n_379), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g471 ( .A(n_379), .Y(n_471) );
INVx1_ASAP7_75t_L g477 ( .A(n_379), .Y(n_477) );
AND2x2_ASAP7_75t_L g502 ( .A(n_379), .B(n_380), .Y(n_502) );
INVx1_ASAP7_75t_L g458 ( .A(n_380), .Y(n_458) );
INVx2_ASAP7_75t_L g464 ( .A(n_380), .Y(n_464) );
INVx1_ASAP7_75t_L g473 ( .A(n_380), .Y(n_473) );
INVx1_ASAP7_75t_L g795 ( .A(n_380), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_380), .B(n_456), .Y(n_869) );
AND2x4_ASAP7_75t_L g472 ( .A(n_381), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g619 ( .A(n_382), .B(n_476), .Y(n_619) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_382), .B(n_476), .Y(n_1105) );
XNOR2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_1363), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_1322), .B2(n_1323), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
XNOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_842), .Y(n_386) );
XOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_626), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_556), .B2(n_557), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g555 ( .A(n_393), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_443), .B1(n_448), .B2(n_489), .C(n_492), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_414), .C(n_424), .D(n_439), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_408), .B2(n_409), .Y(n_395) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_397), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_397), .A2(n_409), .B1(n_703), .B2(n_704), .Y(n_702) );
AOI22xp5_ASAP7_75t_SL g1087 ( .A1(n_397), .A2(n_416), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_397), .A2(n_409), .B1(n_1456), .B2(n_1457), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_397), .A2(n_409), .B1(n_1498), .B2(n_1499), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g1786 ( .A1(n_397), .A2(n_409), .B1(n_1787), .B2(n_1788), .Y(n_1786) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
AND2x6_ASAP7_75t_L g420 ( .A(n_398), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g562 ( .A(n_398), .B(n_401), .Y(n_562) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g943 ( .A(n_399), .B(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g411 ( .A(n_400), .Y(n_411) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
AND2x2_ASAP7_75t_L g528 ( .A(n_400), .B(n_445), .Y(n_528) );
INVx2_ASAP7_75t_L g554 ( .A(n_400), .Y(n_554) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g538 ( .A(n_402), .Y(n_538) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_402), .Y(n_602) );
INVx2_ASAP7_75t_L g605 ( .A(n_402), .Y(n_605) );
INVx2_ASAP7_75t_SL g736 ( .A(n_402), .Y(n_736) );
INVx1_ASAP7_75t_L g928 ( .A(n_402), .Y(n_928) );
INVx1_ASAP7_75t_L g1123 ( .A(n_402), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g1346 ( .A(n_402), .Y(n_1346) );
INVx6_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g416 ( .A(n_403), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g667 ( .A(n_403), .Y(n_667) );
BUFx2_ASAP7_75t_L g895 ( .A(n_403), .Y(n_895) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g412 ( .A(n_405), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g428 ( .A(n_405), .B(n_407), .Y(n_428) );
INVx1_ASAP7_75t_L g435 ( .A(n_406), .Y(n_435) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g422 ( .A(n_407), .B(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_409), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_409), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_409), .A2(n_562), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_409), .A2(n_420), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_409), .A2(n_420), .B1(n_946), .B2(n_947), .Y(n_945) );
CKINVDCx6p67_ASAP7_75t_R g963 ( .A(n_409), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g1096 ( .A1(n_409), .A2(n_420), .B1(n_1097), .B2(n_1098), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_409), .A2(n_420), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_409), .A2(n_562), .B1(n_1370), .B2(n_1371), .Y(n_1369) );
AND2x6_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g441 ( .A(n_410), .Y(n_441) );
INVx1_ASAP7_75t_L g861 ( .A(n_410), .Y(n_861) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_410), .B(n_570), .Y(n_1091) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x6_ASAP7_75t_L g437 ( .A(n_411), .B(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g531 ( .A(n_412), .Y(n_531) );
INVx2_ASAP7_75t_SL g548 ( .A(n_412), .Y(n_548) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_412), .Y(n_597) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_412), .Y(n_658) );
BUFx2_ASAP7_75t_L g740 ( .A(n_412), .Y(n_740) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_412), .Y(n_826) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_412), .Y(n_1006) );
BUFx6f_ASAP7_75t_L g1235 ( .A(n_412), .Y(n_1235) );
HB1xp67_ASAP7_75t_L g1410 ( .A(n_412), .Y(n_1410) );
INVx1_ASAP7_75t_L g820 ( .A(n_413), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_419), .B2(n_420), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_415), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_416), .A2(n_420), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_416), .A2(n_420), .B1(n_641), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_416), .A2(n_420), .B1(n_700), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_416), .A2(n_420), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx4_ASAP7_75t_L g862 ( .A(n_416), .Y(n_862) );
AOI22xp5_ASAP7_75t_SL g1135 ( .A1(n_416), .A2(n_562), .B1(n_1136), .B2(n_1137), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_416), .A2(n_420), .B1(n_1373), .B2(n_1374), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_416), .A2(n_420), .B1(n_1459), .B2(n_1460), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1504 ( .A1(n_416), .A2(n_420), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
AOI22xp33_ASAP7_75t_L g1789 ( .A1(n_416), .A2(n_420), .B1(n_1790), .B2(n_1791), .Y(n_1789) );
AND2x4_ASAP7_75t_L g432 ( .A(n_417), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_417), .B(n_433), .Y(n_711) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx4_ASAP7_75t_L g955 ( .A(n_420), .Y(n_955) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_421), .Y(n_534) );
INVx1_ASAP7_75t_L g837 ( .A(n_421), .Y(n_837) );
BUFx6f_ASAP7_75t_L g1130 ( .A(n_421), .Y(n_1130) );
INVx2_ASAP7_75t_L g1237 ( .A(n_421), .Y(n_1237) );
INVx1_ASAP7_75t_L g1821 ( .A(n_421), .Y(n_1821) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g546 ( .A(n_422), .Y(n_546) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_422), .Y(n_599) );
INVx1_ASAP7_75t_L g742 ( .A(n_422), .Y(n_742) );
INVx1_ASAP7_75t_L g924 ( .A(n_422), .Y(n_924) );
INVx1_ASAP7_75t_L g819 ( .A(n_423), .Y(n_819) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_429), .B2(n_430), .C1(n_436), .C2(n_437), .Y(n_424) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_426), .A2(n_437), .B1(n_711), .B2(n_760), .C1(n_761), .C2(n_762), .Y(n_759) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_427), .Y(n_541) );
INVx1_ASAP7_75t_L g551 ( .A(n_427), .Y(n_551) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_427), .Y(n_606) );
INVx1_ASAP7_75t_L g853 ( .A(n_427), .Y(n_853) );
INVx2_ASAP7_75t_SL g897 ( .A(n_427), .Y(n_897) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_428), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_429), .A2(n_436), .B1(n_466), .B2(n_467), .C1(n_472), .C2(n_474), .Y(n_465) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx4f_ASAP7_75t_L g572 ( .A(n_432), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_432), .A2(n_437), .B1(n_960), .B2(n_961), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_432), .A2(n_437), .B1(n_1028), .B2(n_1029), .Y(n_1073) );
AOI22xp33_ASAP7_75t_SL g1330 ( .A1(n_432), .A2(n_437), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_432), .A2(n_437), .B1(n_1420), .B2(n_1421), .Y(n_1419) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g944 ( .A(n_434), .Y(n_944) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g1015 ( .A(n_435), .Y(n_1015) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_437), .A2(n_568), .B1(n_569), .B2(n_571), .C1(n_572), .C2(n_573), .Y(n_567) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_437), .A2(n_572), .B1(n_637), .B2(n_638), .C1(n_647), .C2(n_648), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g707 ( .A1(n_437), .A2(n_695), .B1(n_696), .B2(n_708), .C1(n_709), .C2(n_711), .Y(n_707) );
AOI222xp33_ASAP7_75t_L g850 ( .A1(n_437), .A2(n_711), .B1(n_851), .B2(n_852), .C1(n_854), .C2(n_855), .Y(n_850) );
AOI222xp33_ASAP7_75t_L g940 ( .A1(n_437), .A2(n_935), .B1(n_936), .B2(n_941), .C1(n_942), .C2(n_943), .Y(n_940) );
INVx3_ASAP7_75t_L g1095 ( .A(n_437), .Y(n_1095) );
AOI222xp33_ASAP7_75t_L g1203 ( .A1(n_437), .A2(n_943), .B1(n_1189), .B2(n_1204), .C1(n_1205), .C2(n_1206), .Y(n_1203) );
AOI222xp33_ASAP7_75t_L g1256 ( .A1(n_437), .A2(n_943), .B1(n_1251), .B2(n_1257), .C1(n_1258), .C2(n_1259), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_437), .A2(n_572), .B1(n_1274), .B2(n_1276), .Y(n_1283) );
AOI222xp33_ASAP7_75t_L g1375 ( .A1(n_437), .A2(n_541), .B1(n_711), .B2(n_1376), .C1(n_1377), .C2(n_1378), .Y(n_1375) );
AOI222xp33_ASAP7_75t_L g1461 ( .A1(n_437), .A2(n_711), .B1(n_737), .B2(n_1462), .C1(n_1463), .C2(n_1464), .Y(n_1461) );
AOI222xp33_ASAP7_75t_L g1500 ( .A1(n_437), .A2(n_550), .B1(n_711), .B2(n_1501), .C1(n_1502), .C2(n_1503), .Y(n_1500) );
AOI222xp33_ASAP7_75t_L g1792 ( .A1(n_437), .A2(n_711), .B1(n_1793), .B2(n_1794), .C1(n_1795), .C2(n_1796), .Y(n_1792) );
BUFx3_ASAP7_75t_L g1017 ( .A(n_438), .Y(n_1017) );
NAND4xp25_ASAP7_75t_SL g559 ( .A(n_439), .B(n_560), .C(n_564), .D(n_567), .Y(n_559) );
BUFx2_ASAP7_75t_L g643 ( .A(n_439), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g752 ( .A(n_439), .B(n_753), .C(n_756), .D(n_759), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g1086 ( .A(n_439), .B(n_1087), .C(n_1090), .D(n_1096), .Y(n_1086) );
NAND4xp25_ASAP7_75t_L g1134 ( .A(n_439), .B(n_1135), .C(n_1138), .D(n_1141), .Y(n_1134) );
NAND4xp25_ASAP7_75t_SL g1368 ( .A(n_439), .B(n_1369), .C(n_1372), .D(n_1375), .Y(n_1368) );
INVx5_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx8_ASAP7_75t_R g712 ( .A(n_440), .Y(n_712) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_442), .Y(n_570) );
INVx2_ASAP7_75t_L g710 ( .A(n_442), .Y(n_710) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_442), .Y(n_738) );
INVx1_ASAP7_75t_L g1125 ( .A(n_442), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_443), .Y(n_574) );
AOI221x1_ASAP7_75t_L g629 ( .A1(n_443), .A2(n_489), .B1(n_630), .B2(n_642), .C(n_653), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_443), .A2(n_489), .B1(n_689), .B2(n_701), .C(n_713), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g1453 ( .A1(n_443), .A2(n_489), .B1(n_1454), .B2(n_1465), .C(n_1475), .Y(n_1453) );
AO211x2_ASAP7_75t_L g1784 ( .A1(n_443), .A2(n_1785), .B(n_1797), .C(n_1806), .Y(n_1784) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
AND2x4_ASAP7_75t_L g863 ( .A(n_444), .B(n_446), .Y(n_863) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g553 ( .A(n_445), .B(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
OR2x6_ASAP7_75t_L g997 ( .A(n_447), .B(n_998), .Y(n_997) );
NAND4xp25_ASAP7_75t_SL g448 ( .A(n_449), .B(n_465), .C(n_481), .D(n_486), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_459), .B2(n_460), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_451), .A2(n_460), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_451), .A2(n_460), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_451), .A2(n_460), .B1(n_691), .B2(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g1106 ( .A1(n_451), .A2(n_483), .B1(n_1107), .B2(n_1108), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_451), .A2(n_483), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_451), .A2(n_1384), .B1(n_1385), .B2(n_1386), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_451), .A2(n_1385), .B1(n_1471), .B2(n_1472), .Y(n_1470) );
AOI22xp33_ASAP7_75t_SL g1522 ( .A1(n_451), .A2(n_1385), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
AOI22xp5_ASAP7_75t_SL g1803 ( .A1(n_451), .A2(n_460), .B1(n_1804), .B2(n_1805), .Y(n_1803) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
AND2x4_ASAP7_75t_L g460 ( .A(n_452), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g867 ( .A(n_452), .Y(n_867) );
AND2x4_ASAP7_75t_L g1385 ( .A(n_452), .B(n_461), .Y(n_1385) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g480 ( .A(n_454), .Y(n_480) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
BUFx2_ASAP7_75t_L g583 ( .A(n_455), .Y(n_583) );
INVx1_ASAP7_75t_L g717 ( .A(n_455), .Y(n_717) );
AND2x2_ASAP7_75t_L g766 ( .A(n_455), .B(n_767), .Y(n_766) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_455), .Y(n_889) );
BUFx6f_ASAP7_75t_L g912 ( .A(n_455), .Y(n_912) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_455), .Y(n_1291) );
INVx1_ASAP7_75t_L g1398 ( .A(n_455), .Y(n_1398) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g783 ( .A(n_456), .Y(n_783) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx5_ASAP7_75t_SL g870 ( .A(n_460), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g1109 ( .A1(n_460), .A2(n_484), .B1(n_1089), .B2(n_1110), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_460), .A2(n_484), .B1(n_1137), .B2(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_462), .Y(n_515) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_463), .Y(n_586) );
INVx1_ASAP7_75t_L g728 ( .A(n_463), .Y(n_728) );
AND2x4_ASAP7_75t_L g470 ( .A(n_464), .B(n_471), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g1146 ( .A1(n_467), .A2(n_487), .B(n_1147), .C(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g892 ( .A(n_468), .Y(n_892) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g693 ( .A1(n_469), .A2(n_472), .B1(n_694), .B2(n_695), .C1(n_696), .C2(n_697), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g1357 ( .A1(n_469), .A2(n_472), .B1(n_697), .B2(n_1331), .C1(n_1332), .C2(n_1358), .Y(n_1357) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_469), .Y(n_1394) );
BUFx2_ASAP7_75t_L g1810 ( .A(n_469), .Y(n_1810) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g487 ( .A(n_470), .B(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_470), .Y(n_505) );
BUFx2_ASAP7_75t_L g592 ( .A(n_470), .Y(n_592) );
INVx1_ASAP7_75t_L g615 ( .A(n_470), .Y(n_615) );
BUFx3_ASAP7_75t_L g805 ( .A(n_470), .Y(n_805) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_470), .Y(n_1103) );
INVx2_ASAP7_75t_L g618 ( .A(n_472), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_472), .A2(n_474), .B1(n_635), .B2(n_636), .C1(n_637), .C2(n_638), .Y(n_634) );
INVx2_ASAP7_75t_L g876 ( .A(n_472), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_472), .A2(n_474), .B1(n_935), .B2(n_936), .Y(n_934) );
INVx2_ASAP7_75t_L g971 ( .A(n_472), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_472), .A2(n_474), .B1(n_1205), .B2(n_1206), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_472), .A2(n_474), .B1(n_1258), .B2(n_1259), .Y(n_1263) );
AOI222xp33_ASAP7_75t_L g1273 ( .A1(n_472), .A2(n_474), .B1(n_505), .B2(n_1274), .C1(n_1275), .C2(n_1276), .Y(n_1273) );
AOI222xp33_ASAP7_75t_SL g1424 ( .A1(n_472), .A2(n_697), .B1(n_1420), .B2(n_1421), .C1(n_1425), .C2(n_1426), .Y(n_1424) );
INVx1_ASAP7_75t_L g777 ( .A(n_473), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_474), .A2(n_854), .B1(n_855), .B2(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_474), .A2(n_960), .B1(n_961), .B2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_474), .A2(n_875), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .Y(n_474) );
AND2x4_ASAP7_75t_L g697 ( .A(n_475), .B(n_478), .Y(n_697) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g794 ( .A(n_477), .B(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_477), .B(n_795), .Y(n_1175) );
INVxp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g488 ( .A(n_479), .Y(n_488) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_480), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_483), .A2(n_565), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_483), .A2(n_625), .B1(n_640), .B2(n_641), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_483), .A2(n_625), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_483), .A2(n_484), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_483), .A2(n_625), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
AOI22xp33_ASAP7_75t_SL g1387 ( .A1(n_483), .A2(n_484), .B1(n_1373), .B2(n_1388), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_483), .A2(n_625), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_483), .A2(n_484), .B1(n_1459), .B2(n_1474), .Y(n_1473) );
AOI22xp33_ASAP7_75t_SL g1525 ( .A1(n_483), .A2(n_484), .B1(n_1505), .B2(n_1526), .Y(n_1525) );
AOI22xp5_ASAP7_75t_L g1798 ( .A1(n_483), .A2(n_484), .B1(n_1790), .B2(n_1799), .Y(n_1798) );
INVx5_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g625 ( .A(n_485), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_486), .B(n_631), .C(n_634), .D(n_639), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g689 ( .A(n_486), .B(n_690), .C(n_693), .D(n_698), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g1272 ( .A(n_486), .B(n_1273), .C(n_1277), .Y(n_1272) );
NAND3xp33_ASAP7_75t_L g1356 ( .A(n_486), .B(n_1357), .C(n_1359), .Y(n_1356) );
NAND3xp33_ASAP7_75t_SL g1423 ( .A(n_486), .B(n_1424), .C(n_1427), .Y(n_1423) );
CKINVDCx11_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
AOI211xp5_ASAP7_75t_SL g613 ( .A1(n_487), .A2(n_614), .B(n_616), .C(n_617), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g1100 ( .A1(n_487), .A2(n_1101), .B(n_1102), .C(n_1104), .Y(n_1100) );
AOI211xp5_ASAP7_75t_L g1380 ( .A1(n_487), .A2(n_722), .B(n_1381), .C(n_1382), .Y(n_1380) );
AOI211xp5_ASAP7_75t_L g1466 ( .A1(n_487), .A2(n_1467), .B(n_1468), .C(n_1469), .Y(n_1466) );
AOI211xp5_ASAP7_75t_L g1519 ( .A1(n_487), .A2(n_722), .B(n_1520), .C(n_1521), .Y(n_1519) );
AOI211xp5_ASAP7_75t_L g1800 ( .A1(n_487), .A2(n_614), .B(n_1801), .C(n_1802), .Y(n_1800) );
OAI31xp33_ASAP7_75t_L g864 ( .A1(n_489), .A2(n_865), .A3(n_871), .B(n_877), .Y(n_864) );
OAI31xp33_ASAP7_75t_SL g929 ( .A1(n_489), .A2(n_930), .A3(n_931), .B(n_937), .Y(n_929) );
OAI31xp33_ASAP7_75t_L g964 ( .A1(n_489), .A2(n_965), .A3(n_966), .B(n_972), .Y(n_964) );
OAI31xp33_ASAP7_75t_L g1023 ( .A1(n_489), .A2(n_1024), .A3(n_1025), .B(n_1030), .Y(n_1023) );
OAI31xp33_ASAP7_75t_SL g1208 ( .A1(n_489), .A2(n_1209), .A3(n_1210), .B(n_1212), .Y(n_1208) );
OAI31xp33_ASAP7_75t_SL g1260 ( .A1(n_489), .A2(n_1261), .A3(n_1262), .B(n_1264), .Y(n_1260) );
O2A1O1Ixp33_ASAP7_75t_L g1270 ( .A1(n_489), .A2(n_1271), .B(n_1272), .C(n_1280), .Y(n_1270) );
OAI21xp5_ASAP7_75t_L g1355 ( .A1(n_489), .A2(n_1356), .B(n_1362), .Y(n_1355) );
OAI21xp5_ASAP7_75t_L g1422 ( .A1(n_489), .A2(n_1423), .B(n_1430), .Y(n_1422) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
AOI31xp33_ASAP7_75t_L g612 ( .A1(n_490), .A2(n_613), .A3(n_620), .B(n_623), .Y(n_612) );
AOI31xp33_ASAP7_75t_L g1379 ( .A1(n_490), .A2(n_1380), .A3(n_1383), .B(n_1387), .Y(n_1379) );
AOI31xp33_ASAP7_75t_L g1797 ( .A1(n_490), .A2(n_1798), .A3(n_1800), .B(n_1803), .Y(n_1797) );
AND2x4_ASAP7_75t_L g552 ( .A(n_491), .B(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g906 ( .A(n_491), .B(n_553), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_524), .Y(n_492) );
AOI33xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .A3(n_506), .B1(n_513), .B2(n_516), .B3(n_518), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g1431 ( .A1(n_494), .A2(n_518), .B1(n_1432), .B2(n_1438), .C(n_1444), .Y(n_1431) );
BUFx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g672 ( .A(n_495), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_495), .B(n_715), .C(n_721), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_495), .B(n_880), .C(n_883), .Y(n_879) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_495), .B(n_911), .C(n_914), .Y(n_910) );
NAND3xp33_ASAP7_75t_L g1113 ( .A(n_495), .B(n_1114), .C(n_1115), .Y(n_1113) );
NAND3xp33_ASAP7_75t_L g1155 ( .A(n_495), .B(n_1156), .C(n_1157), .Y(n_1155) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_495), .B(n_1391), .C(n_1393), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1479 ( .A(n_495), .B(n_1480), .C(n_1483), .Y(n_1479) );
AOI33xp33_ASAP7_75t_L g1513 ( .A1(n_495), .A2(n_906), .A3(n_1514), .B1(n_1515), .B2(n_1516), .B3(n_1517), .Y(n_1513) );
NAND3xp33_ASAP7_75t_L g1807 ( .A(n_495), .B(n_1808), .C(n_1809), .Y(n_1807) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
OR2x6_ASAP7_75t_L g526 ( .A(n_496), .B(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g577 ( .A(n_496), .B(n_497), .Y(n_577) );
BUFx2_ASAP7_75t_L g813 ( .A(n_496), .Y(n_813) );
OR2x2_ASAP7_75t_L g900 ( .A(n_496), .B(n_901), .Y(n_900) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_496), .B(n_798), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_496), .B(n_527), .Y(n_1217) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g675 ( .A(n_500), .Y(n_675) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g807 ( .A(n_501), .B(n_767), .Y(n_807) );
INVx3_ASAP7_75t_L g885 ( .A(n_501), .Y(n_885) );
BUFx2_ASAP7_75t_L g891 ( .A(n_501), .Y(n_891) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g581 ( .A(n_502), .Y(n_581) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g517 ( .A(n_504), .Y(n_517) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_505), .Y(n_722) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g1055 ( .A(n_510), .Y(n_1055) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g790 ( .A(n_511), .Y(n_790) );
INVx2_ASAP7_75t_L g913 ( .A(n_511), .Y(n_913) );
INVx2_ASAP7_75t_L g918 ( .A(n_511), .Y(n_918) );
INVx2_ASAP7_75t_L g994 ( .A(n_511), .Y(n_994) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g678 ( .A(n_512), .Y(n_678) );
INVx3_ASAP7_75t_L g720 ( .A(n_512), .Y(n_720) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI33xp33_ASAP7_75t_L g576 ( .A1(n_518), .A2(n_577), .A3(n_578), .B1(n_582), .B2(n_587), .B3(n_589), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_518), .B(n_917), .C(n_919), .Y(n_916) );
INVx2_ASAP7_75t_L g987 ( .A(n_518), .Y(n_987) );
INVx1_ASAP7_75t_L g1067 ( .A(n_518), .Y(n_1067) );
INVx6_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g683 ( .A(n_519), .Y(n_683) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g798 ( .A(n_522), .Y(n_798) );
AOI33xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_529), .A3(n_535), .B1(n_542), .B2(n_549), .B3(n_552), .Y(n_524) );
AOI33xp33_ASAP7_75t_L g593 ( .A1(n_525), .A2(n_594), .A3(n_600), .B1(n_603), .B2(n_607), .B3(n_611), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_525), .B(n_733), .C(n_739), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g655 ( .A(n_526), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_526), .A2(n_838), .B1(n_1033), .B2(n_1038), .Y(n_1032) );
OAI22xp5_ASAP7_75t_SL g1306 ( .A1(n_526), .A2(n_669), .B1(n_1307), .B2(n_1311), .Y(n_1306) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g901 ( .A(n_528), .Y(n_901) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_538), .Y(n_661) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g1794 ( .A(n_540), .Y(n_1794) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_541), .Y(n_662) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g1411 ( .A(n_544), .Y(n_1411) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_545), .Y(n_1045) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g1037 ( .A(n_548), .Y(n_1037) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx4f_ASAP7_75t_L g611 ( .A(n_552), .Y(n_611) );
INVx4_ASAP7_75t_L g669 ( .A(n_552), .Y(n_669) );
BUFx4f_ASAP7_75t_L g839 ( .A(n_552), .Y(n_839) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AOI211xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_574), .B(n_575), .C(n_612), .Y(n_558) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI221x1_ASAP7_75t_L g751 ( .A1(n_574), .A2(n_752), .B1(n_763), .B2(n_811), .C(n_814), .Y(n_751) );
OAI31xp33_ASAP7_75t_L g953 ( .A1(n_574), .A2(n_954), .A3(n_956), .B(n_962), .Y(n_953) );
INVx1_ASAP7_75t_L g1287 ( .A(n_574), .Y(n_1287) );
AOI211xp5_ASAP7_75t_L g1367 ( .A1(n_574), .A2(n_1368), .B(n_1379), .C(n_1389), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_593), .Y(n_575) );
BUFx2_ASAP7_75t_L g1339 ( .A(n_577), .Y(n_1339) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g731 ( .A(n_581), .Y(n_731) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_581), .Y(n_1403) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
BUFx3_ASAP7_75t_L g588 ( .A(n_586), .Y(n_588) );
INVx4_ASAP7_75t_L g1337 ( .A(n_586), .Y(n_1337) );
INVx2_ASAP7_75t_SL g1434 ( .A(n_586), .Y(n_1434) );
INVx1_ASAP7_75t_L g1302 ( .A(n_588), .Y(n_1302) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g636 ( .A(n_591), .Y(n_636) );
INVx1_ASAP7_75t_L g1426 ( .A(n_591), .Y(n_1426) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g608 ( .A(n_596), .Y(n_608) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx3_ASAP7_75t_L g746 ( .A(n_597), .Y(n_746) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g610 ( .A(n_599), .Y(n_610) );
BUFx3_ASAP7_75t_L g747 ( .A(n_599), .Y(n_747) );
INVx1_ASAP7_75t_L g1222 ( .A(n_599), .Y(n_1222) );
INVx1_ASAP7_75t_L g1318 ( .A(n_599), .Y(n_1318) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_605), .Y(n_1316) );
BUFx2_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_611), .B(n_744), .C(n_745), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g1351 ( .A(n_611), .B(n_1352), .C(n_1353), .Y(n_1351) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_685), .B1(n_840), .B2(n_841), .Y(n_626) );
INVx2_ASAP7_75t_SL g840 ( .A(n_627), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g1562 ( .A1(n_628), .A2(n_1563), .B1(n_1564), .B2(n_1566), .Y(n_1562) );
INVx1_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
NAND4xp25_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .C(n_646), .D(n_649), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_670), .Y(n_653) );
AOI33xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .A3(n_659), .B1(n_663), .B2(n_664), .B3(n_668), .Y(n_654) );
INVx1_ASAP7_75t_L g827 ( .A(n_655), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g1814 ( .A(n_655), .B(n_1815), .C(n_1816), .Y(n_1814) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx3_ASAP7_75t_L g1313 ( .A(n_658), .Y(n_1313) );
INVx2_ASAP7_75t_L g1349 ( .A(n_658), .Y(n_1349) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g904 ( .A(n_667), .Y(n_904) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI22xp5_ASAP7_75t_SL g1191 ( .A1(n_669), .A2(n_900), .B1(n_1192), .B2(n_1195), .Y(n_1191) );
OAI22xp5_ASAP7_75t_SL g1444 ( .A1(n_669), .A2(n_1217), .B1(n_1445), .B2(n_1447), .Y(n_1444) );
AOI33xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .A3(n_676), .B1(n_679), .B2(n_680), .B3(n_681), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_671), .A2(n_681), .B1(n_1289), .B2(n_1299), .C(n_1306), .Y(n_1288) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g1184 ( .A(n_678), .Y(n_1184) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
CKINVDCx8_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_683), .B(n_724), .C(n_729), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_683), .B(n_888), .C(n_890), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g1340 ( .A(n_683), .B(n_1341), .C(n_1342), .Y(n_1340) );
NAND3xp33_ASAP7_75t_L g1395 ( .A(n_683), .B(n_1396), .C(n_1401), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1476 ( .A(n_683), .B(n_1477), .C(n_1478), .Y(n_1476) );
NAND3xp33_ASAP7_75t_L g1811 ( .A(n_683), .B(n_1812), .C(n_1813), .Y(n_1811) );
INVx1_ASAP7_75t_L g841 ( .A(n_685), .Y(n_841) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_750), .Y(n_686) );
INVx1_ASAP7_75t_L g749 ( .A(n_688), .Y(n_749) );
NAND4xp25_ASAP7_75t_SL g701 ( .A(n_702), .B(n_705), .C(n_707), .D(n_712), .Y(n_701) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g1257 ( .A(n_710), .Y(n_1257) );
NAND3xp33_ASAP7_75t_SL g849 ( .A(n_712), .B(n_850), .C(n_856), .Y(n_849) );
NAND3xp33_ASAP7_75t_SL g939 ( .A(n_712), .B(n_940), .C(n_945), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g1202 ( .A(n_712), .B(n_1203), .Y(n_1202) );
NAND2xp5_ASAP7_75t_SL g1255 ( .A(n_712), .B(n_1256), .Y(n_1255) );
NAND4xp25_ASAP7_75t_L g1454 ( .A(n_712), .B(n_1455), .C(n_1458), .D(n_1461), .Y(n_1454) );
NAND4xp25_ASAP7_75t_L g1496 ( .A(n_712), .B(n_1497), .C(n_1500), .D(n_1504), .Y(n_1496) );
NAND4xp25_ASAP7_75t_SL g1785 ( .A(n_712), .B(n_1786), .C(n_1789), .D(n_1792), .Y(n_1785) );
NAND4xp25_ASAP7_75t_SL g713 ( .A(n_714), .B(n_723), .C(n_732), .D(n_743), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g791 ( .A(n_717), .Y(n_791) );
INVx1_ASAP7_75t_L g1439 ( .A(n_717), .Y(n_1439) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g1392 ( .A(n_719), .Y(n_1392) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g882 ( .A(n_720), .Y(n_882) );
INVx1_ASAP7_75t_L g1181 ( .A(n_720), .Y(n_1181) );
INVx2_ASAP7_75t_L g1400 ( .A(n_720), .Y(n_1400) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g772 ( .A(n_728), .Y(n_772) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_731), .B(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g1354 ( .A(n_742), .Y(n_1354) );
AOI222xp33_ASAP7_75t_L g802 ( .A1(n_757), .A2(n_803), .B1(n_804), .B2(n_806), .C1(n_807), .C2(n_808), .Y(n_802) );
OAI21xp5_ASAP7_75t_SL g792 ( .A1(n_760), .A2(n_793), .B(n_796), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_773), .C(n_802), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_768), .B2(n_769), .Y(n_764) );
INVx2_ASAP7_75t_L g771 ( .A(n_767), .Y(n_771) );
AND2x4_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
AND2x4_ASAP7_75t_L g804 ( .A(n_770), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g1482 ( .A(n_772), .Y(n_1482) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_789), .C(n_799), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g775 ( .A(n_776), .B(n_778), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OR2x6_ASAP7_75t_L g782 ( .A(n_779), .B(n_783), .Y(n_782) );
OR2x6_ASAP7_75t_L g800 ( .A(n_779), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g810 ( .A(n_779), .Y(n_810) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_788), .Y(n_784) );
OAI221xp5_ASAP7_75t_SL g815 ( .A1(n_787), .A2(n_816), .B1(n_821), .B2(n_823), .C(n_824), .Y(n_815) );
INVx1_ASAP7_75t_L g1060 ( .A(n_790), .Y(n_1060) );
INVx1_ASAP7_75t_L g968 ( .A(n_793), .Y(n_968) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_793), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_793), .A2(n_1242), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_793), .A2(n_984), .B1(n_1442), .B2(n_1443), .Y(n_1441) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g801 ( .A(n_794), .Y(n_801) );
BUFx2_ASAP7_75t_L g873 ( .A(n_794), .Y(n_873) );
INVx2_ASAP7_75t_L g1065 ( .A(n_794), .Y(n_1065) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g933 ( .A(n_801), .Y(n_933) );
OAI221xp5_ASAP7_75t_SL g828 ( .A1(n_803), .A2(n_806), .B1(n_829), .B2(n_832), .C(n_835), .Y(n_828) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_805), .Y(n_886) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
CKINVDCx8_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_827), .B1(n_828), .B2(n_838), .Y(n_814) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g831 ( .A(n_818), .Y(n_831) );
OR2x2_ASAP7_75t_L g860 ( .A(n_818), .B(n_861), .Y(n_860) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_818), .Y(n_1039) );
INVx1_ASAP7_75t_L g1226 ( .A(n_818), .Y(n_1226) );
OR2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
AND2x2_ASAP7_75t_L g822 ( .A(n_819), .B(n_820), .Y(n_822) );
INVx1_ASAP7_75t_L g1003 ( .A(n_821), .Y(n_1003) );
BUFx3_ASAP7_75t_L g1308 ( .A(n_821), .Y(n_1308) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g834 ( .A(n_822), .Y(n_834) );
INVx1_ASAP7_75t_L g958 ( .A(n_822), .Y(n_958) );
INVx1_ASAP7_75t_L g1042 ( .A(n_822), .Y(n_1042) );
BUFx4f_ASAP7_75t_L g1229 ( .A(n_822), .Y(n_1229) );
BUFx4f_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1220 ( .A(n_826), .Y(n_1220) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g1000 ( .A(n_831), .Y(n_1000) );
INVx2_ASAP7_75t_L g1193 ( .A(n_831), .Y(n_1193) );
INVx2_ASAP7_75t_L g1196 ( .A(n_831), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g1195 ( .A1(n_833), .A2(n_1196), .B1(n_1197), .B2(n_1198), .C(n_1199), .Y(n_1195) );
INVx2_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1007 ( .A(n_837), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_838), .A2(n_989), .B1(n_997), .B2(n_999), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_839), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g1817 ( .A(n_839), .B(n_1818), .C(n_1819), .Y(n_1817) );
AO22x2_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_1267), .B1(n_1320), .B2(n_1321), .Y(n_842) );
INVx1_ASAP7_75t_L g1320 ( .A(n_843), .Y(n_1320) );
XNOR2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_1080), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_950), .B1(n_1078), .B2(n_1079), .Y(n_844) );
INVx2_ASAP7_75t_L g1078 ( .A(n_845), .Y(n_1078) );
XOR2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_907), .Y(n_845) );
NAND3x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_864), .C(n_878), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_859), .B(n_863), .Y(n_848) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g942 ( .A(n_853), .Y(n_942) );
OAI21xp5_ASAP7_75t_SL g938 ( .A1(n_863), .A2(n_939), .B(n_948), .Y(n_938) );
OAI31xp33_ASAP7_75t_SL g1068 ( .A1(n_863), .A2(n_1069), .A3(n_1070), .B(n_1074), .Y(n_1068) );
AOI211xp5_ASAP7_75t_L g1085 ( .A1(n_863), .A2(n_1086), .B(n_1099), .C(n_1112), .Y(n_1085) );
AOI211xp5_ASAP7_75t_L g1133 ( .A1(n_863), .A2(n_1134), .B(n_1145), .C(n_1154), .Y(n_1133) );
OAI31xp33_ASAP7_75t_SL g1200 ( .A1(n_863), .A2(n_1201), .A3(n_1202), .B(n_1207), .Y(n_1200) );
OAI31xp33_ASAP7_75t_L g1252 ( .A1(n_863), .A2(n_1253), .A3(n_1254), .B(n_1255), .Y(n_1252) );
OAI31xp33_ASAP7_75t_L g1326 ( .A1(n_863), .A2(n_1327), .A3(n_1328), .B(n_1329), .Y(n_1326) );
OAI31xp33_ASAP7_75t_SL g1415 ( .A1(n_863), .A2(n_1416), .A3(n_1417), .B(n_1418), .Y(n_1415) );
AOI211x1_ASAP7_75t_L g1495 ( .A1(n_863), .A2(n_1496), .B(n_1507), .C(n_1518), .Y(n_1495) );
OR2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx2_ASAP7_75t_L g991 ( .A(n_868), .Y(n_991) );
BUFx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g979 ( .A(n_869), .Y(n_979) );
INVx1_ASAP7_75t_L g1053 ( .A(n_869), .Y(n_1053) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g986 ( .A(n_873), .Y(n_986) );
INVx1_ASAP7_75t_L g1048 ( .A(n_873), .Y(n_1048) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AND4x1_ASAP7_75t_L g878 ( .A(n_879), .B(n_887), .C(n_893), .D(n_902), .Y(n_878) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx2_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g915 ( .A(n_885), .Y(n_915) );
INVx2_ASAP7_75t_L g1116 ( .A(n_885), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1467 ( .A(n_886), .Y(n_1467) );
NAND3xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_898), .C(n_899), .Y(n_893) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_895), .Y(n_1009) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g1204 ( .A(n_897), .Y(n_1204) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_899), .B(n_921), .C(n_922), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g1121 ( .A(n_899), .B(n_1122), .C(n_1126), .Y(n_1121) );
NAND3xp33_ASAP7_75t_L g1161 ( .A(n_899), .B(n_1162), .C(n_1163), .Y(n_1161) );
NAND3xp33_ASAP7_75t_L g1404 ( .A(n_899), .B(n_1405), .C(n_1406), .Y(n_1404) );
NAND3xp33_ASAP7_75t_L g1486 ( .A(n_899), .B(n_1487), .C(n_1489), .Y(n_1486) );
AOI33xp33_ASAP7_75t_L g1508 ( .A1(n_899), .A2(n_1120), .A3(n_1509), .B1(n_1510), .B2(n_1511), .B3(n_1512), .Y(n_1508) );
INVx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .C(n_906), .Y(n_902) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_906), .B(n_926), .C(n_927), .Y(n_925) );
NAND3xp33_ASAP7_75t_L g1127 ( .A(n_906), .B(n_1128), .C(n_1129), .Y(n_1127) );
NAND3xp33_ASAP7_75t_L g1164 ( .A(n_906), .B(n_1165), .C(n_1166), .Y(n_1164) );
INVx1_ASAP7_75t_L g1239 ( .A(n_906), .Y(n_1239) );
NAND3xp33_ASAP7_75t_L g1407 ( .A(n_906), .B(n_1408), .C(n_1409), .Y(n_1407) );
NAND3xp33_ASAP7_75t_L g1490 ( .A(n_906), .B(n_1491), .C(n_1492), .Y(n_1490) );
XOR2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_949), .Y(n_907) );
NAND3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_929), .C(n_938), .Y(n_908) );
AND4x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_916), .C(n_920), .D(n_925), .Y(n_909) );
INVx1_ASAP7_75t_L g981 ( .A(n_913), .Y(n_981) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g1094 ( .A(n_943), .Y(n_1094) );
INVx1_ASAP7_75t_L g1144 ( .A(n_943), .Y(n_1144) );
INVx1_ASAP7_75t_L g1079 ( .A(n_950), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_1020), .B1(n_1021), .B2(n_1077), .Y(n_950) );
INVx1_ASAP7_75t_L g1077 ( .A(n_951), .Y(n_1077) );
INVx1_ASAP7_75t_L g1018 ( .A(n_952), .Y(n_1018) );
NAND3xp33_ASAP7_75t_L g952 ( .A(n_953), .B(n_964), .C(n_973), .Y(n_952) );
HB1xp67_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
NOR3xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_988), .C(n_1008), .Y(n_973) );
NOR3xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_982), .C(n_987), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .B1(n_980), .B2(n_981), .Y(n_975) );
BUFx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx2_ASAP7_75t_L g1179 ( .A(n_979), .Y(n_1179) );
INVx1_ASAP7_75t_L g1246 ( .A(n_979), .Y(n_1246) );
OAI22xp33_ASAP7_75t_SL g982 ( .A1(n_983), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_982) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_984), .A2(n_1034), .B1(n_1035), .B2(n_1048), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1172 ( .A1(n_984), .A2(n_1173), .B1(n_1174), .B2(n_1176), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_992), .B1(n_993), .B2(n_995), .C(n_996), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI33xp33_ASAP7_75t_L g1046 ( .A1(n_997), .A2(n_1047), .A3(n_1049), .B1(n_1056), .B2(n_1061), .B3(n_1067), .Y(n_1046) );
OAI33xp33_ASAP7_75t_L g1171 ( .A1(n_997), .A2(n_1172), .A3(n_1177), .B1(n_1182), .B2(n_1186), .B3(n_1190), .Y(n_1171) );
OAI33xp33_ASAP7_75t_L g1240 ( .A1(n_997), .A2(n_1190), .A3(n_1241), .B1(n_1244), .B2(n_1245), .B3(n_1249), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1001), .B1(n_1002), .B2(n_1004), .C(n_1005), .Y(n_999) );
OAI221xp5_ASAP7_75t_L g1033 ( .A1(n_1000), .A2(n_1002), .B1(n_1034), .B2(n_1035), .C(n_1036), .Y(n_1033) );
OAI21xp33_ASAP7_75t_SL g1010 ( .A1(n_1002), .A2(n_1011), .B(n_1012), .Y(n_1010) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1022), .Y(n_1075) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1031), .C(n_1068), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1046), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1040), .B1(n_1041), .B2(n_1043), .C(n_1044), .Y(n_1038) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1042), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1051), .B1(n_1054), .B2(n_1055), .Y(n_1049) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1052), .Y(n_1058) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_SL g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1059), .B2(n_1060), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1064), .B1(n_1065), .B2(n_1066), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
OAI22xp33_ASAP7_75t_L g1186 ( .A1(n_1065), .A2(n_1187), .B1(n_1188), .B2(n_1189), .Y(n_1186) );
OAI221xp5_ASAP7_75t_L g1192 ( .A1(n_1071), .A2(n_1173), .B1(n_1176), .B2(n_1193), .C(n_1194), .Y(n_1192) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
XOR2x2_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1167), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1083), .B1(n_1131), .B2(n_1132), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
XNOR2xp5_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
AOI21xp5_ASAP7_75t_L g1090 ( .A1(n_1091), .A2(n_1092), .B(n_1093), .Y(n_1090) );
AOI21xp5_ASAP7_75t_L g1141 ( .A1(n_1091), .A2(n_1142), .B(n_1143), .Y(n_1141) );
AOI31xp33_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1106), .A3(n_1109), .B(n_1111), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
AOI31xp33_ASAP7_75t_L g1145 ( .A1(n_1111), .A2(n_1146), .A3(n_1149), .B(n_1152), .Y(n_1145) );
AOI31xp33_ASAP7_75t_L g1518 ( .A1(n_1111), .A2(n_1519), .A3(n_1522), .B(n_1525), .Y(n_1518) );
NAND4xp25_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1117), .C(n_1121), .D(n_1127), .Y(n_1112) );
NAND3xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1119), .C(n_1120), .Y(n_1117) );
NAND3xp33_ASAP7_75t_L g1158 ( .A(n_1120), .B(n_1159), .C(n_1160), .Y(n_1158) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1120), .Y(n_1190) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND4xp25_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1158), .C(n_1161), .D(n_1164), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1213), .B1(n_1265), .B2(n_1266), .Y(n_1167) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1168), .Y(n_1265) );
NAND3xp33_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1200), .C(n_1208), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1191), .Y(n_1170) );
OAI22xp33_ASAP7_75t_L g1241 ( .A1(n_1174), .A2(n_1224), .B1(n_1227), .B2(n_1242), .Y(n_1241) );
INVx2_ASAP7_75t_L g1298 ( .A(n_1174), .Y(n_1298) );
BUFx3_ASAP7_75t_L g1305 ( .A(n_1174), .Y(n_1305) );
BUFx6f_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
OAI22xp33_ASAP7_75t_SL g1177 ( .A1(n_1178), .A2(n_1179), .B1(n_1180), .B2(n_1181), .Y(n_1177) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1179), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_1179), .A2(n_1184), .B1(n_1219), .B2(n_1221), .Y(n_1244) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1181), .Y(n_1440) );
OAI22xp33_ASAP7_75t_L g1245 ( .A1(n_1184), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1307 ( .A1(n_1196), .A2(n_1293), .B1(n_1296), .B2(n_1308), .C(n_1309), .Y(n_1307) );
OAI221xp5_ASAP7_75t_L g1445 ( .A1(n_1196), .A2(n_1308), .B1(n_1442), .B2(n_1443), .C(n_1446), .Y(n_1445) );
OAI221xp5_ASAP7_75t_L g1447 ( .A1(n_1196), .A2(n_1425), .B1(n_1428), .B2(n_1448), .C(n_1449), .Y(n_1447) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1213), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1252), .C(n_1260), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1240), .Y(n_1215) );
OAI33xp33_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1218), .A3(n_1223), .B1(n_1230), .B2(n_1233), .B3(n_1239), .Y(n_1216) );
INVx1_ASAP7_75t_SL g1350 ( .A(n_1217), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1220), .B1(n_1221), .B2(n_1222), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B1(n_1227), .B2(n_1228), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_1225), .A2(n_1228), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1229), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_1234), .A2(n_1236), .B1(n_1237), .B2(n_1238), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
BUFx3_ASAP7_75t_L g1310 ( .A(n_1235), .Y(n_1310) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1267), .Y(n_1321) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1288), .Y(n_1269) );
OAI221xp5_ASAP7_75t_L g1311 ( .A1(n_1275), .A2(n_1308), .B1(n_1312), .B2(n_1314), .C(n_1315), .Y(n_1311) );
AOI21xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1284), .B(n_1287), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
OAI22xp5_ASAP7_75t_SL g1292 ( .A1(n_1293), .A2(n_1294), .B1(n_1296), .B2(n_1297), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_1294), .A2(n_1297), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
INVx3_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
OAI22xp33_ASAP7_75t_SL g1300 ( .A1(n_1301), .A2(n_1302), .B1(n_1303), .B2(n_1304), .Y(n_1300) );
BUFx3_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
NAND3x1_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1333), .C(n_1355), .Y(n_1325) );
AND4x1_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1340), .C(n_1343), .D(n_1351), .Y(n_1333) );
NAND3xp33_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1338), .C(n_1339), .Y(n_1334) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1347), .C(n_1350), .Y(n_1343) );
INVx4_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1346), .Y(n_1488) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
AO22x2_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1450), .B1(n_1451), .B2(n_1530), .Y(n_1363) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1364), .Y(n_1530) );
XNOR2xp5_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1413), .Y(n_1364) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1367), .Y(n_1412) );
NAND4xp25_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1395), .C(n_1404), .D(n_1407), .Y(n_1389) );
INVx2_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
INVx2_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
BUFx2_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1403), .Y(n_1485) );
NAND3x1_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1422), .C(n_1431), .Y(n_1414) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVxp67_ASAP7_75t_SL g1450 ( .A(n_1451), .Y(n_1450) );
AOI22xp5_ASAP7_75t_L g1451 ( .A1(n_1452), .A2(n_1493), .B1(n_1494), .B2(n_1529), .Y(n_1451) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1452), .Y(n_1529) );
NAND3xp33_ASAP7_75t_L g1465 ( .A(n_1466), .B(n_1470), .C(n_1473), .Y(n_1465) );
NAND4xp25_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1479), .C(n_1486), .D(n_1490), .Y(n_1475) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx2_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1495), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1507 ( .A(n_1508), .B(n_1513), .Y(n_1507) );
OAI221xp5_ASAP7_75t_R g1531 ( .A1(n_1532), .A2(n_1779), .B1(n_1780), .B2(n_1822), .C(n_1828), .Y(n_1531) );
NOR3xp33_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1749), .C(n_1776), .Y(n_1532) );
AOI33xp33_ASAP7_75t_L g1533 ( .A1(n_1534), .A2(n_1629), .A3(n_1674), .B1(n_1701), .B2(n_1720), .B3(n_1736), .Y(n_1533) );
AOI211xp5_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1578), .B(n_1601), .C(n_1618), .Y(n_1534) );
NOR2xp33_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1559), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_1536), .B(n_1628), .Y(n_1627) );
NOR2x1_ASAP7_75t_R g1660 ( .A(n_1536), .B(n_1661), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1536), .B(n_1616), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1741 ( .A(n_1536), .B(n_1723), .Y(n_1741) );
AOI211xp5_ASAP7_75t_SL g1752 ( .A1(n_1536), .A2(n_1600), .B(n_1753), .C(n_1754), .Y(n_1752) );
INVx2_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1537), .B(n_1609), .Y(n_1608) );
INVx2_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx4_ASAP7_75t_L g1625 ( .A(n_1538), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1631 ( .A(n_1538), .B(n_1632), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1538), .B(n_1600), .Y(n_1655) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1538), .B(n_1589), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1692 ( .A(n_1538), .B(n_1626), .Y(n_1692) );
NOR2xp33_ASAP7_75t_L g1706 ( .A(n_1538), .B(n_1600), .Y(n_1706) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1538), .B(n_1610), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1538), .B(n_1561), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1538), .B(n_1644), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1538), .B(n_1598), .Y(n_1751) );
AOI21xp5_ASAP7_75t_L g1763 ( .A1(n_1538), .A2(n_1651), .B(n_1660), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1538), .B(n_1611), .Y(n_1767) );
AND2x6_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1551), .Y(n_1538) );
AND2x4_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1546), .Y(n_1540) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
OR2x2_ASAP7_75t_L g1565 ( .A(n_1542), .B(n_1547), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1545), .Y(n_1542) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1545), .Y(n_1554) );
AND2x4_ASAP7_75t_L g1548 ( .A(n_1546), .B(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1547), .B(n_1550), .Y(n_1568) );
HB1xp67_ASAP7_75t_L g1837 ( .A(n_1549), .Y(n_1837) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1552), .Y(n_1571) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1552), .Y(n_1667) );
AND2x4_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1555), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1553), .B(n_1555), .Y(n_1577) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
AND2x4_ASAP7_75t_L g1558 ( .A(n_1554), .B(n_1555), .Y(n_1558) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g1665 ( .A1(n_1557), .A2(n_1666), .B1(n_1667), .B2(n_1668), .Y(n_1665) );
INVx2_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_SL g1573 ( .A(n_1558), .Y(n_1573) );
OAI222xp33_ASAP7_75t_L g1630 ( .A1(n_1559), .A2(n_1631), .B1(n_1635), .B2(n_1638), .C1(n_1641), .C2(n_1643), .Y(n_1630) );
OAI321xp33_ASAP7_75t_L g1766 ( .A1(n_1559), .A2(n_1694), .A3(n_1722), .B1(n_1767), .B2(n_1768), .C(n_1770), .Y(n_1766) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1560), .B(n_1610), .Y(n_1683) );
AOI221xp5_ASAP7_75t_L g1701 ( .A1(n_1560), .A2(n_1606), .B1(n_1702), .B2(n_1711), .C(n_1712), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1574), .Y(n_1560) );
INVx3_ASAP7_75t_L g1605 ( .A(n_1561), .Y(n_1605) );
OR2x2_ASAP7_75t_L g1619 ( .A(n_1561), .B(n_1620), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1569), .Y(n_1561) );
OAI22xp5_ASAP7_75t_L g1586 ( .A1(n_1564), .A2(n_1568), .B1(n_1587), .B2(n_1588), .Y(n_1586) );
OAI22xp33_ASAP7_75t_L g1613 ( .A1(n_1564), .A2(n_1568), .B1(n_1614), .B2(n_1615), .Y(n_1613) );
BUFx3_ASAP7_75t_L g1671 ( .A(n_1564), .Y(n_1671) );
BUFx6f_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
OAI22xp5_ASAP7_75t_L g1594 ( .A1(n_1565), .A2(n_1568), .B1(n_1595), .B2(n_1596), .Y(n_1594) );
HB1xp67_ASAP7_75t_L g1673 ( .A(n_1566), .Y(n_1673) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1569 ( .A1(n_1570), .A2(n_1571), .B1(n_1572), .B2(n_1573), .Y(n_1569) );
OAI22xp5_ASAP7_75t_L g1582 ( .A1(n_1573), .A2(n_1583), .B1(n_1584), .B2(n_1585), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1574), .B(n_1612), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1574), .B(n_1611), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1574), .B(n_1611), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1574), .B(n_1605), .Y(n_1653) );
INVx2_ASAP7_75t_L g1659 ( .A(n_1574), .Y(n_1659) );
OAI22xp5_ASAP7_75t_L g1726 ( .A1(n_1574), .A2(n_1699), .B1(n_1727), .B2(n_1729), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1574), .B(n_1612), .Y(n_1734) );
AOI221xp5_ASAP7_75t_L g1750 ( .A1(n_1574), .A2(n_1734), .B1(n_1751), .B2(n_1752), .C(n_1756), .Y(n_1750) );
AND2x4_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1576), .Y(n_1574) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1577), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1597), .Y(n_1578) );
OAI22xp33_ASAP7_75t_L g1732 ( .A1(n_1579), .A2(n_1703), .B1(n_1733), .B2(n_1735), .Y(n_1732) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1589), .Y(n_1580) );
CKINVDCx6p67_ASAP7_75t_R g1600 ( .A(n_1581), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1581), .B(n_1617), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1581), .B(n_1624), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1581), .B(n_1633), .Y(n_1632) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1581), .B(n_1599), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1581), .B(n_1642), .Y(n_1641) );
OR2x2_ASAP7_75t_L g1686 ( .A(n_1581), .B(n_1626), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1581), .B(n_1599), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1581), .B(n_1647), .Y(n_1769) );
OR2x6_ASAP7_75t_SL g1581 ( .A(n_1582), .B(n_1586), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1589), .B(n_1625), .Y(n_1642) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1589), .B(n_1655), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1589), .B(n_1600), .Y(n_1698) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1589), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1593), .Y(n_1589) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1590), .Y(n_1599) );
OR2x2_ASAP7_75t_L g1626 ( .A(n_1590), .B(n_1593), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1590), .B(n_1634), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1593), .B(n_1599), .Y(n_1617) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1593), .Y(n_1634) );
NOR2xp33_ASAP7_75t_L g1695 ( .A(n_1593), .B(n_1600), .Y(n_1695) );
OAI22xp5_ASAP7_75t_L g1618 ( .A1(n_1597), .A2(n_1619), .B1(n_1621), .B2(n_1627), .Y(n_1618) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1600), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1651 ( .A(n_1600), .B(n_1633), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1600), .B(n_1617), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1600), .B(n_1642), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1600), .B(n_1634), .Y(n_1737) );
OAI322xp33_ASAP7_75t_L g1740 ( .A1(n_1600), .A2(n_1686), .A3(n_1690), .B1(n_1741), .B2(n_1742), .C1(n_1744), .C2(n_1745), .Y(n_1740) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1600), .B(n_1743), .Y(n_1742) );
OR2x2_ASAP7_75t_L g1755 ( .A(n_1600), .B(n_1634), .Y(n_1755) );
NOR2xp33_ASAP7_75t_L g1765 ( .A(n_1600), .B(n_1681), .Y(n_1765) );
INVxp67_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1606), .Y(n_1602) );
O2A1O1Ixp33_ASAP7_75t_L g1693 ( .A1(n_1603), .A2(n_1627), .B(n_1694), .C(n_1696), .Y(n_1693) );
INVx1_ASAP7_75t_SL g1603 ( .A(n_1604), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1604), .B(n_1676), .Y(n_1675) );
INVx3_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1605), .B(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1605), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1605), .B(n_1611), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1605), .B(n_1610), .Y(n_1719) );
O2A1O1Ixp33_ASAP7_75t_SL g1776 ( .A1(n_1605), .A2(n_1620), .B(n_1777), .C(n_1778), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1607), .B(n_1616), .Y(n_1606) );
NOR2xp33_ASAP7_75t_L g1652 ( .A(n_1607), .B(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1610), .Y(n_1656) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1610), .Y(n_1689) );
INVx2_ASAP7_75t_SL g1610 ( .A(n_1611), .Y(n_1610) );
INVx2_ASAP7_75t_SL g1611 ( .A(n_1612), .Y(n_1611) );
HB1xp67_ASAP7_75t_L g1680 ( .A(n_1612), .Y(n_1680) );
NOR2xp33_ASAP7_75t_L g1635 ( .A(n_1616), .B(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1617), .Y(n_1661) );
OAI22xp5_ASAP7_75t_L g1762 ( .A1(n_1619), .A2(n_1739), .B1(n_1763), .B2(n_1764), .Y(n_1762) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1620), .Y(n_1640) );
INVxp67_ASAP7_75t_SL g1621 ( .A(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
AOI22xp33_ASAP7_75t_L g1716 ( .A1(n_1624), .A2(n_1688), .B1(n_1717), .B2(n_1719), .Y(n_1716) );
NOR2xp33_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1625), .B(n_1640), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1625), .B(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1625), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1625), .B(n_1725), .Y(n_1724) );
O2A1O1Ixp33_ASAP7_75t_L g1774 ( .A1(n_1625), .A2(n_1661), .B(n_1682), .C(n_1775), .Y(n_1774) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1626), .Y(n_1647) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1627), .Y(n_1648) );
AOI221xp5_ASAP7_75t_L g1720 ( .A1(n_1628), .A2(n_1721), .B1(n_1724), .B2(n_1726), .C(n_1732), .Y(n_1720) );
INVx2_ASAP7_75t_L g1723 ( .A(n_1628), .Y(n_1723) );
NOR3xp33_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1645), .C(n_1649), .Y(n_1629) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1631), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1633), .B(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1633), .Y(n_1730) );
NAND3xp33_ASAP7_75t_L g1770 ( .A(n_1636), .B(n_1723), .C(n_1743), .Y(n_1770) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
AOI211xp5_ASAP7_75t_SL g1760 ( .A1(n_1644), .A2(n_1761), .B(n_1762), .C(n_1766), .Y(n_1760) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1648), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1647), .B(n_1706), .Y(n_1705) );
NAND3xp33_ASAP7_75t_L g1713 ( .A(n_1647), .B(n_1659), .C(n_1714), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1647), .B(n_1655), .Y(n_1759) );
OAI221xp5_ASAP7_75t_L g1649 ( .A1(n_1650), .A2(n_1652), .B1(n_1654), .B2(n_1656), .C(n_1657), .Y(n_1649) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
AOI221xp5_ASAP7_75t_L g1771 ( .A1(n_1653), .A2(n_1697), .B1(n_1704), .B2(n_1772), .C(n_1774), .Y(n_1771) );
NAND2xp5_ASAP7_75t_L g1773 ( .A(n_1653), .B(n_1656), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1654), .B(n_1679), .Y(n_1678) );
A2O1A1Ixp33_ASAP7_75t_SL g1696 ( .A1(n_1656), .A2(n_1697), .B(n_1698), .C(n_1699), .Y(n_1696) );
AOI21xp5_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1660), .B(n_1662), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1687 ( .A(n_1658), .B(n_1680), .Y(n_1687) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1658), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1739 ( .A(n_1658), .B(n_1680), .Y(n_1739) );
OAI321xp33_ASAP7_75t_L g1677 ( .A1(n_1659), .A2(n_1661), .A3(n_1678), .B1(n_1681), .B2(n_1682), .C(n_1684), .Y(n_1677) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1659), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1661), .B(n_1730), .Y(n_1744) );
CKINVDCx14_ASAP7_75t_R g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
NAND3xp33_ASAP7_75t_SL g1712 ( .A(n_1664), .B(n_1713), .C(n_1716), .Y(n_1712) );
OR2x6_ASAP7_75t_SL g1664 ( .A(n_1665), .B(n_1669), .Y(n_1664) );
OAI22xp5_ASAP7_75t_L g1669 ( .A1(n_1670), .A2(n_1671), .B1(n_1672), .B2(n_1673), .Y(n_1669) );
BUFx2_ASAP7_75t_SL g1779 ( .A(n_1673), .Y(n_1779) );
NOR3xp33_ASAP7_75t_SL g1674 ( .A(n_1675), .B(n_1677), .C(n_1693), .Y(n_1674) );
INVxp67_ASAP7_75t_L g1778 ( .A(n_1675), .Y(n_1778) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1680), .Y(n_1758) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1681), .Y(n_1697) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
AOI22xp33_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1687), .B1(n_1688), .B2(n_1691), .Y(n_1684) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1690), .B(n_1723), .Y(n_1722) );
OAI211xp5_ASAP7_75t_L g1749 ( .A1(n_1690), .A2(n_1750), .B(n_1760), .C(n_1771), .Y(n_1749) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
NOR2xp33_ASAP7_75t_L g1746 ( .A(n_1694), .B(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1698), .Y(n_1777) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1707), .Y(n_1702) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1706), .Y(n_1731) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1710), .Y(n_1775) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1719), .Y(n_1745) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
OR2x2_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1731), .Y(n_1729) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
AOI211xp5_ASAP7_75t_L g1736 ( .A1(n_1737), .A2(n_1738), .B(n_1740), .C(n_1746), .Y(n_1736) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
OR2x2_ASAP7_75t_L g1757 ( .A(n_1758), .B(n_1759), .Y(n_1757) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1784), .Y(n_1831) );
NAND4xp25_ASAP7_75t_L g1806 ( .A(n_1807), .B(n_1811), .C(n_1814), .D(n_1817), .Y(n_1806) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
CKINVDCx14_ASAP7_75t_R g1822 ( .A(n_1823), .Y(n_1822) );
INVx4_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
INVxp33_ASAP7_75t_L g1829 ( .A(n_1830), .Y(n_1829) );
HB1xp67_ASAP7_75t_SL g1832 ( .A(n_1833), .Y(n_1832) );
OAI21xp5_ASAP7_75t_L g1836 ( .A1(n_1834), .A2(n_1837), .B(n_1838), .Y(n_1836) );
BUFx2_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
endmodule