module fake_ariane_1538_n_2491 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_2491);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2491;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_645;
wire n_559;
wire n_2233;
wire n_2370;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2427;
wire n_2098;
wire n_661;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1443;
wire n_1021;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_1442;
wire n_696;
wire n_482;
wire n_798;
wire n_1833;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_436;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1832;
wire n_767;
wire n_1392;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_2294;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_1592;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2122;
wire n_1611;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_1609;
wire n_600;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_439;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_2075;
wire n_1726;
wire n_699;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_536;
wire n_1162;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_501;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1733;
wire n_640;
wire n_1856;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1258;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1429;
wire n_2064;
wire n_1324;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1955;
wire n_1504;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1584;
wire n_1157;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1381;
wire n_1124;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_671;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1777;
wire n_1019;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1821;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_2052;
wire n_1091;
wire n_2485;
wire n_1063;
wire n_537;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_2239;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1870;
wire n_1299;
wire n_2063;
wire n_1925;
wire n_782;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_157),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_368),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_120),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_227),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_314),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_8),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_94),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_83),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_259),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_4),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_297),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_22),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_293),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_322),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_340),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_392),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_142),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_281),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_65),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_90),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_90),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_375),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_329),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_88),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_129),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_4),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_60),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_258),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_348),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_302),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_266),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_401),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_128),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_125),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_285),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_57),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_98),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_206),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_366),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_378),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_196),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_86),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_250),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_306),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_296),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_128),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_269),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_339),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_332),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_84),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_5),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_312),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_341),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_309),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_75),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_315),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_362),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_203),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_187),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_133),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_351),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_151),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_168),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_245),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_397),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_299),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_261),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_110),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_188),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_134),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_2),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_307),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_336),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_171),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_57),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_189),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_28),
.Y(n_491)
);

BUFx5_ASAP7_75t_L g492 ( 
.A(n_271),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_394),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_294),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_228),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_199),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_256),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_303),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_273),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_173),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_238),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_373),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_210),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_277),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_328),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_140),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_355),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_387),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_107),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_67),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_126),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_376),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_212),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_383),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_36),
.Y(n_515)
);

BUFx5_ASAP7_75t_L g516 ( 
.A(n_335),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_47),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_3),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_353),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_154),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_382),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_248),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_174),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_182),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_185),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_95),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_308),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_317),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_324),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_398),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_158),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_357),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_252),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_177),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_124),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_72),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_246),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_342),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_52),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_327),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_62),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_113),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_7),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_224),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_205),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_221),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_163),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_338),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_169),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_260),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_82),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_96),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_170),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_354),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_54),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_112),
.Y(n_556)
);

BUFx5_ASAP7_75t_L g557 ( 
.A(n_323),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_166),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_96),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_272),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_21),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_222),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_218),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_326),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_325),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_59),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_409),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_164),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_113),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_181),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_275),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_44),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_391),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_358),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_230),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_287),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_384),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_136),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_84),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_18),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_231),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_330),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_333),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_50),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_404),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_379),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_10),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_356),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_304),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_369),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_237),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_148),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_3),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_385),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_47),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_180),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_51),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_241),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_119),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_380),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_360),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_30),
.Y(n_602)
);

BUFx5_ASAP7_75t_L g603 ( 
.A(n_215),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_292),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_236),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_301),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_76),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_17),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_300),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_214),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_162),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_178),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_280),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_359),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_207),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_406),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_6),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_28),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_48),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_122),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_345),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_127),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_343),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_43),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_405),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_270),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_33),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_377),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_235),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_289),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_129),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_400),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_61),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_364),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_114),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_388),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_263),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_29),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_53),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_201),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_349),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_240),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_41),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_12),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_242),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_132),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_86),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_255),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_254),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_37),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_46),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_371),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_58),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_95),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_8),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_239),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_372),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_62),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_251),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_265),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_316),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_17),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_318),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_107),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_386),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_202),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_192),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_346),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_184),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_313),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_399),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_408),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_89),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_337),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_70),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_71),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_193),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_175),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_19),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_305),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_82),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_198),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_361),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_2),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_77),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_89),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_11),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_298),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_213),
.Y(n_689)
);

CKINVDCx16_ASAP7_75t_R g690 ( 
.A(n_390),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_58),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_268),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_0),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_146),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_370),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_147),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_64),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_45),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_229),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_41),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_319),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_290),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_363),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_71),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_253),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_321),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_25),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_396),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_367),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_75),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_365),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_320),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_115),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_1),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_347),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_141),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_40),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_51),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_61),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_191),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_311),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_217),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_68),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_195),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_334),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_352),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_121),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_101),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_389),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_33),
.Y(n_730)
);

BUFx8_ASAP7_75t_SL g731 ( 
.A(n_407),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_21),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_284),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_161),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_24),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_87),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_194),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_22),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_186),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_291),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_72),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_279),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_32),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_52),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_35),
.Y(n_745)
);

CKINVDCx12_ASAP7_75t_R g746 ( 
.A(n_310),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_165),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_344),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_59),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_350),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_232),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_395),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_16),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_149),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_44),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_283),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_381),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_731),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_412),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_412),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_480),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_480),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_622),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_654),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_654),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_731),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_717),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_717),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_419),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_419),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_595),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_419),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_579),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_419),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_602),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_419),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_419),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_595),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_419),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_416),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_428),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_437),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_446),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_443),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_442),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_607),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_509),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_429),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_510),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_511),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_535),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_442),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_429),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_541),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_555),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_607),
.Y(n_797)
);

INVxp33_ASAP7_75t_L g798 ( 
.A(n_631),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_434),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_556),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_559),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_580),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_593),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_643),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_617),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_644),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_651),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_664),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_681),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_684),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_643),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_687),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_691),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_700),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_497),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_487),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_589),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_497),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_704),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_495),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_710),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_713),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_459),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_743),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_620),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_496),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_744),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_745),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_620),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_653),
.Y(n_830)
);

CKINVDCx14_ASAP7_75t_R g831 ( 
.A(n_610),
.Y(n_831)
);

CKINVDCx16_ASAP7_75t_R g832 ( 
.A(n_641),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_733),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_690),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_653),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_635),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_415),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_673),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_673),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_517),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_655),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_686),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_507),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_417),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_421),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_736),
.Y(n_846)
);

INVxp33_ASAP7_75t_SL g847 ( 
.A(n_520),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_470),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_553),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_705),
.Y(n_850)
);

INVxp33_ASAP7_75t_SL g851 ( 
.A(n_430),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_482),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_662),
.Y(n_853)
);

BUFx2_ASAP7_75t_SL g854 ( 
.A(n_610),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_544),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_563),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_435),
.Y(n_857)
);

INVxp33_ASAP7_75t_SL g858 ( 
.A(n_436),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_444),
.Y(n_859)
);

CKINVDCx16_ASAP7_75t_R g860 ( 
.A(n_517),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_583),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_463),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_606),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_553),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_647),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_677),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_734),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_610),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_647),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_722),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_448),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_588),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_449),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_588),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_722),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_613),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_725),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_725),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_613),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_676),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_517),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_725),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_720),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_740),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_740),
.Y(n_886)
);

INVx4_ASAP7_75t_R g887 ( 
.A(n_720),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_740),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_697),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_697),
.Y(n_890)
);

INVxp33_ASAP7_75t_SL g891 ( 
.A(n_454),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_697),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_414),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_754),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_422),
.Y(n_895)
);

CKINVDCx16_ASAP7_75t_R g896 ( 
.A(n_422),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_754),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_418),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_447),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_458),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_420),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_426),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_440),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_441),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_445),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_450),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_462),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_456),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_464),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_447),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_465),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_466),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_468),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_473),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_476),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_575),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_575),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_489),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_478),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_481),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_484),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_485),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_486),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_488),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_585),
.Y(n_925)
);

INVxp33_ASAP7_75t_L g926 ( 
.A(n_529),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_503),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_529),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_519),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_585),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_524),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_467),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_530),
.Y(n_933)
);

INVxp33_ASAP7_75t_SL g934 ( 
.A(n_483),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_531),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_533),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_540),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_545),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_590),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_547),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_590),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_550),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_614),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_560),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_515),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_526),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_565),
.Y(n_947)
);

INVxp33_ASAP7_75t_L g948 ( 
.A(n_605),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_571),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_586),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_591),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_676),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_628),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_646),
.Y(n_954)
);

INVxp33_ASAP7_75t_SL g955 ( 
.A(n_536),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_648),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_663),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_670),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_680),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_688),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_701),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_708),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_512),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_539),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_737),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_757),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_746),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_542),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_605),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_543),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_755),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_551),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_552),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_561),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_566),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_572),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_584),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_597),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_629),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_629),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_640),
.Y(n_981)
);

INVxp33_ASAP7_75t_SL g982 ( 
.A(n_599),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_608),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_618),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_492),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_492),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_619),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_640),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_624),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_627),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_492),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_492),
.Y(n_992)
);

CKINVDCx14_ASAP7_75t_R g993 ( 
.A(n_614),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_633),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_638),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_650),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_658),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_569),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_675),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_679),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_685),
.Y(n_1001)
);

CKINVDCx16_ASAP7_75t_R g1002 ( 
.A(n_668),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_656),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_693),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_698),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_707),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_492),
.Y(n_1007)
);

INVxp33_ASAP7_75t_L g1008 ( 
.A(n_656),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_706),
.B(n_0),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_714),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_718),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_719),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_723),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_727),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_728),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_730),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_732),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_735),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_738),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_741),
.Y(n_1020)
);

INVxp33_ASAP7_75t_SL g1021 ( 
.A(n_749),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_753),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_706),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_410),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_742),
.Y(n_1025)
);

INVxp33_ASAP7_75t_SL g1026 ( 
.A(n_491),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_742),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_411),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_501),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_668),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_492),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_623),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_513),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_703),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_755),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_518),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_587),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_413),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_423),
.Y(n_1039)
);

INVxp67_ASAP7_75t_SL g1040 ( 
.A(n_512),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_512),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_424),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_758),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_769),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_1024),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_786),
.B(n_469),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_786),
.B(n_471),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_963),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_963),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_818),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_963),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_882),
.B(n_868),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_963),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_771),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_847),
.B(n_490),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_985),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_985),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_770),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_818),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_847),
.B(n_564),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_772),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_831),
.B(n_702),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_849),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_986),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_986),
.Y(n_1065)
);

BUFx8_ASAP7_75t_SL g1066 ( 
.A(n_771),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_849),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_793),
.B(n_425),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_969),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_766),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_979),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_979),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_793),
.B(n_427),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_815),
.B(n_431),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_831),
.B(n_678),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_774),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_981),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_815),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_991),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_854),
.B(n_678),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_776),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_870),
.B(n_432),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_777),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_864),
.B(n_433),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_882),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_763),
.Y(n_1087)
);

BUFx8_ASAP7_75t_SL g1088 ( 
.A(n_778),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_875),
.B(n_877),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_991),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_864),
.B(n_438),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_872),
.B(n_439),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_981),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_992),
.Y(n_1094)
);

BUFx8_ASAP7_75t_L g1095 ( 
.A(n_836),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_992),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_988),
.Y(n_1097)
);

CKINVDCx6p67_ASAP7_75t_R g1098 ( 
.A(n_832),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_872),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_773),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_779),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_SL g1102 ( 
.A1(n_778),
.A2(n_581),
.B1(n_452),
.B2(n_453),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_780),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_926),
.B(n_948),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_782),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_783),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_785),
.Y(n_1107)
);

BUFx8_ASAP7_75t_SL g1108 ( 
.A(n_787),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_988),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1007),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_784),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1031),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1038),
.B(n_451),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1003),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1031),
.A2(n_516),
.B(n_492),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_1003),
.Y(n_1116)
);

BUFx8_ASAP7_75t_SL g1117 ( 
.A(n_787),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_820),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_876),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_788),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_876),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_926),
.B(n_455),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_898),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_898),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_790),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_837),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_915),
.A2(n_557),
.B(n_516),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_878),
.B(n_512),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_894),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_894),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_897),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1039),
.B(n_457),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_SL g1133 ( 
.A(n_834),
.B(n_460),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_897),
.Y(n_1134)
);

BUFx8_ASAP7_75t_SL g1135 ( 
.A(n_797),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_915),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_845),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_759),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_829),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_948),
.B(n_1008),
.Y(n_1140)
);

AND2x6_ASAP7_75t_L g1141 ( 
.A(n_923),
.B(n_554),
.Y(n_1141)
);

BUFx8_ASAP7_75t_SL g1142 ( 
.A(n_797),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_781),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1009),
.A2(n_756),
.B(n_472),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_791),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_823),
.Y(n_1146)
);

BUFx8_ASAP7_75t_SL g1147 ( 
.A(n_804),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_760),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_923),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_935),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_848),
.A2(n_474),
.B1(n_475),
.B2(n_461),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_935),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_775),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_792),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_826),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_830),
.Y(n_1156)
);

BUFx8_ASAP7_75t_L g1157 ( 
.A(n_932),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_795),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_835),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_944),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_944),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_796),
.Y(n_1162)
);

OAI22x1_ASAP7_75t_SL g1163 ( 
.A1(n_804),
.A2(n_479),
.B1(n_493),
.B2(n_477),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_879),
.B(n_752),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_857),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_947),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_800),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_947),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_949),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_R g1170 ( 
.A(n_848),
.B(n_494),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_801),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_899),
.B(n_498),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_859),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_844),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_871),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_820),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_949),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_883),
.B(n_554),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_802),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_803),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_805),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_838),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1008),
.B(n_499),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_885),
.B(n_554),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_873),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_761),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_811),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_839),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_833),
.Y(n_1189)
);

AOI22x1_ASAP7_75t_SL g1190 ( 
.A1(n_925),
.A2(n_502),
.B1(n_504),
.B2(n_500),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_886),
.B(n_505),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_806),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_SL g1193 ( 
.A1(n_811),
.A2(n_508),
.B1(n_514),
.B2(n_506),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_807),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_808),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_820),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_809),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1023),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_925),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_762),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_888),
.B(n_554),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_910),
.B(n_521),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1025),
.Y(n_1203)
);

OA21x2_ASAP7_75t_L g1204 ( 
.A1(n_1027),
.A2(n_1041),
.B(n_1040),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_945),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_930),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_810),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_764),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_812),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_907),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_765),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_767),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_993),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_768),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_813),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_814),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_819),
.Y(n_1217)
);

AND2x2_ASAP7_75t_SL g1218 ( 
.A(n_1009),
.B(n_558),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_946),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_821),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_893),
.A2(n_523),
.B(n_522),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_798),
.B(n_525),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_928),
.B(n_527),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_964),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_822),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_840),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1086),
.B(n_889),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1208),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1101),
.B(n_874),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1211),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1212),
.Y(n_1231)
);

BUFx8_ASAP7_75t_L g1232 ( 
.A(n_1146),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1214),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1079),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1119),
.Y(n_1236)
);

CKINVDCx16_ASAP7_75t_R g1237 ( 
.A(n_1155),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1119),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1119),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1079),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1099),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1129),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1153),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1086),
.B(n_1042),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1099),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1215),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1101),
.B(n_880),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1129),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1129),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1071),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1216),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1131),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1138),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1044),
.B(n_884),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1067),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1138),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1148),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1131),
.Y(n_1258)
);

AND2x6_ASAP7_75t_L g1259 ( 
.A(n_1062),
.B(n_558),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1059),
.B(n_890),
.Y(n_1260)
);

OR2x6_ASAP7_75t_L g1261 ( 
.A(n_1226),
.B(n_1036),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1127),
.A2(n_902),
.B(n_901),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1148),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1200),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1067),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1107),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1058),
.B(n_980),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1061),
.B(n_903),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1131),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1071),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1071),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1072),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1182),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1077),
.B(n_904),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1072),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1200),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1121),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1130),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1136),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1072),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1189),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1153),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1087),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1073),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1104),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1182),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1115),
.A2(n_906),
.B(n_905),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1073),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1087),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1136),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1073),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1078),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_SL g1293 ( 
.A(n_1218),
.B(n_1026),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1078),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1067),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1182),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1136),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1082),
.B(n_908),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1188),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1078),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1140),
.B(n_860),
.Y(n_1301)
);

AND2x2_ASAP7_75t_SL g1302 ( 
.A(n_1218),
.B(n_895),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1149),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1084),
.B(n_909),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1093),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1093),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1188),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1172),
.B(n_1202),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1056),
.B(n_911),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1149),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1188),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1093),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1097),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1149),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1152),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1213),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1152),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1172),
.B(n_968),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1097),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1152),
.Y(n_1320)
);

BUFx8_ASAP7_75t_L g1321 ( 
.A(n_1043),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1097),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1076),
.B(n_558),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1114),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1114),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1114),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1116),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1057),
.A2(n_913),
.B(n_912),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1160),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1064),
.B(n_914),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1160),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1116),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1059),
.B(n_1063),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1116),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1063),
.B(n_1050),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1050),
.B(n_892),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1069),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1069),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1065),
.B(n_919),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1080),
.A2(n_921),
.B(n_920),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1161),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1052),
.B(n_967),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1090),
.B(n_922),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1100),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1161),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1161),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1166),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1166),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1166),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1177),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1096),
.B(n_924),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1177),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1109),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1055),
.A2(n_1032),
.B1(n_1026),
.B2(n_853),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1110),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1055),
.B(n_816),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1222),
.B(n_798),
.Y(n_1358)
);

AND2x6_ASAP7_75t_L g1359 ( 
.A(n_1112),
.B(n_558),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1060),
.A2(n_858),
.B1(n_891),
.B2(n_851),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1177),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1134),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1202),
.B(n_970),
.Y(n_1363)
);

BUFx8_ASAP7_75t_L g1364 ( 
.A(n_1070),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1134),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1103),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1105),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1106),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1204),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1066),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1068),
.A2(n_929),
.B(n_927),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1139),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1156),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1111),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1174),
.B(n_816),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1120),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1125),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1145),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1213),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1154),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1159),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1049),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1126),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1223),
.B(n_973),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1198),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1109),
.B(n_931),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1094),
.B(n_933),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1068),
.A2(n_937),
.B(n_936),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1049),
.Y(n_1389)
);

NAND2xp33_ASAP7_75t_L g1390 ( 
.A(n_1266),
.B(n_1165),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1308),
.B(n_1060),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1362),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1308),
.B(n_1122),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1293),
.A2(n_1204),
.B1(n_1102),
.B2(n_940),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1293),
.B(n_1045),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1243),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1282),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1312),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1238),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1318),
.B(n_1183),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1366),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1367),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1356),
.Y(n_1403)
);

AND2x6_ASAP7_75t_L g1404 ( 
.A(n_1369),
.B(n_1081),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1227),
.B(n_1205),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1356),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1372),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1227),
.B(n_1205),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1285),
.B(n_1384),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1358),
.B(n_1137),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1238),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1312),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1238),
.Y(n_1413)
);

AND3x2_ASAP7_75t_L g1414 ( 
.A(n_1383),
.B(n_1185),
.C(n_1133),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1368),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1234),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1360),
.B(n_1045),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1261),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1318),
.A2(n_1133),
.B1(n_1221),
.B2(n_1089),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1363),
.A2(n_1221),
.B1(n_1089),
.B2(n_1170),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1363),
.B(n_1046),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1360),
.B(n_1165),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1374),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1285),
.B(n_1083),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1173),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1232),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1373),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1381),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1302),
.B(n_1173),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1385),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1384),
.B(n_1083),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1365),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1302),
.A2(n_942),
.B1(n_950),
.B2(n_938),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1228),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1357),
.B(n_1164),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1376),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1378),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1230),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1231),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1244),
.B(n_1046),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1380),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1277),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1233),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1278),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1335),
.B(n_1175),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1328),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1266),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1333),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1361),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1357),
.B(n_1164),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1313),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1283),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1244),
.B(n_1191),
.Y(n_1454)
);

CKINVDCx6p67_ASAP7_75t_R g1455 ( 
.A(n_1237),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1338),
.B(n_1191),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1361),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1246),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1251),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1235),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1240),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1335),
.B(n_1175),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1328),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1345),
.B(n_799),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1261),
.B(n_1199),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1309),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1309),
.Y(n_1467)
);

AND2x6_ASAP7_75t_L g1468 ( 
.A(n_1369),
.B(n_1052),
.Y(n_1468)
);

BUFx10_ASAP7_75t_L g1469 ( 
.A(n_1281),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1330),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1330),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_R g1472 ( 
.A(n_1281),
.B(n_993),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1241),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1371),
.B(n_1047),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1245),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1232),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1340),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1261),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1371),
.B(n_1047),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1341),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1242),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1242),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1301),
.Y(n_1483)
);

BUFx10_ASAP7_75t_L g1484 ( 
.A(n_1370),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1340),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1229),
.B(n_1247),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1355),
.A2(n_1345),
.B1(n_1274),
.B2(n_1298),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1344),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1248),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1344),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1355),
.B(n_1219),
.Y(n_1491)
);

AND2x6_ASAP7_75t_L g1492 ( 
.A(n_1343),
.B(n_1128),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1248),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1316),
.B(n_1206),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1388),
.A2(n_1075),
.B(n_1074),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1338),
.B(n_1113),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1248),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1333),
.B(n_1219),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1229),
.B(n_1223),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1249),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1249),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1249),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1283),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1269),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1323),
.A2(n_1170),
.B1(n_1178),
.B2(n_1128),
.Y(n_1505)
);

BUFx10_ASAP7_75t_L g1506 ( 
.A(n_1370),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1247),
.B(n_1178),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1354),
.B(n_1113),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1269),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1386),
.B(n_1132),
.C(n_1075),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1289),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1379),
.B(n_1224),
.Y(n_1512)
);

CKINVDCx6p67_ASAP7_75t_R g1513 ( 
.A(n_1289),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1354),
.B(n_1132),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1321),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1269),
.Y(n_1516)
);

INVxp33_ASAP7_75t_L g1517 ( 
.A(n_1343),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1352),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1273),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1313),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1321),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1273),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1273),
.Y(n_1523)
);

AND2x6_ASAP7_75t_L g1524 ( 
.A(n_1253),
.B(n_1184),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1286),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1337),
.B(n_1260),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1286),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1286),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1352),
.Y(n_1529)
);

NAND3xp33_ASAP7_75t_L g1530 ( 
.A(n_1386),
.B(n_1085),
.C(n_1074),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1268),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1296),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1265),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1407),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1447),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1391),
.B(n_1254),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1391),
.B(n_1254),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1416),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1409),
.B(n_1267),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1398),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1533),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1463),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1533),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1526),
.B(n_1339),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1395),
.B(n_1224),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1427),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1401),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1533),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1402),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1415),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1398),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1423),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1339),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1436),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1425),
.B(n_1410),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1398),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1409),
.B(n_1267),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1437),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1431),
.A2(n_939),
.B1(n_941),
.B2(n_930),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1431),
.B(n_939),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1395),
.B(n_1337),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1438),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1396),
.B(n_941),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1396),
.B(n_896),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1397),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1453),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1454),
.B(n_1326),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1403),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1498),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1426),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1511),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1515),
.Y(n_1572)
);

INVx4_ASAP7_75t_L g1573 ( 
.A(n_1449),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1421),
.B(n_1259),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1428),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1513),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1430),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1449),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1454),
.B(n_1393),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1394),
.A2(n_943),
.B1(n_1259),
.B2(n_1323),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1406),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1464),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1442),
.Y(n_1583)
);

BUFx4f_ASAP7_75t_L g1584 ( 
.A(n_1455),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1498),
.Y(n_1585)
);

AO22x2_ASAP7_75t_L g1586 ( 
.A1(n_1487),
.A2(n_918),
.B1(n_998),
.B2(n_862),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1466),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1412),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1503),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1503),
.B(n_943),
.C(n_974),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1452),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1421),
.B(n_916),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1443),
.Y(n_1594)
);

OR2x2_ASAP7_75t_SL g1595 ( 
.A(n_1414),
.B(n_917),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1418),
.B(n_1260),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1467),
.Y(n_1597)
);

AND2x6_ASAP7_75t_L g1598 ( 
.A(n_1505),
.B(n_1256),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1448),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1439),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1440),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1517),
.B(n_1002),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1444),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1470),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1390),
.B(n_997),
.C(n_976),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1520),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1471),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1458),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1477),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1400),
.A2(n_1030),
.B1(n_1210),
.B2(n_1174),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1520),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1422),
.B(n_865),
.Y(n_1612)
);

AND2x6_ASAP7_75t_L g1613 ( 
.A(n_1505),
.B(n_1257),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1399),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1483),
.B(n_1210),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1459),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1476),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1465),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1485),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1399),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1393),
.B(n_1400),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1460),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1478),
.B(n_1255),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1394),
.A2(n_1404),
.B1(n_1491),
.B2(n_1433),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_1531),
.B(n_1323),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1488),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1465),
.B(n_1265),
.Y(n_1627)
);

INVx5_ASAP7_75t_L g1628 ( 
.A(n_1468),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1465),
.Y(n_1629)
);

AO22x2_ASAP7_75t_L g1630 ( 
.A1(n_1487),
.A2(n_869),
.B1(n_881),
.B2(n_865),
.Y(n_1630)
);

NAND3x1_ASAP7_75t_L g1631 ( 
.A(n_1435),
.B(n_1088),
.C(n_1066),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1411),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_SL g1633 ( 
.A(n_1521),
.B(n_1364),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1569),
.B(n_1494),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1566),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1560),
.B(n_1417),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1583),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1585),
.B(n_1512),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1571),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1555),
.B(n_1593),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1538),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1600),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1583),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1563),
.B(n_1054),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1579),
.A2(n_1530),
.B(n_1510),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1621),
.B(n_1441),
.Y(n_1647)
);

OR2x6_ASAP7_75t_L g1648 ( 
.A(n_1570),
.B(n_1494),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1541),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1539),
.B(n_1441),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1603),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1589),
.B(n_1424),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1557),
.B(n_1499),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1565),
.B(n_1424),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1610),
.B(n_1435),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1608),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1584),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1559),
.A2(n_1429),
.B1(n_1451),
.B2(n_817),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1587),
.B(n_1499),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1545),
.B(n_1054),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1564),
.B(n_1187),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1587),
.B(n_1433),
.Y(n_1663)
);

O2A1O1Ixp5_ASAP7_75t_L g1664 ( 
.A1(n_1567),
.A2(n_1451),
.B(n_1508),
.C(n_1496),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1572),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1597),
.B(n_1490),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1630),
.A2(n_858),
.B1(n_934),
.B2(n_891),
.C(n_851),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1597),
.B(n_1518),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1547),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1604),
.B(n_1486),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1604),
.B(n_1486),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1607),
.B(n_1529),
.Y(n_1672)
);

NOR2xp67_ASAP7_75t_L g1673 ( 
.A(n_1599),
.B(n_1510),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1607),
.B(n_1609),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1630),
.A2(n_869),
.B1(n_952),
.B2(n_881),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1609),
.B(n_1496),
.Y(n_1676)
);

BUFx5_ASAP7_75t_L g1677 ( 
.A(n_1535),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1549),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1612),
.B(n_1187),
.Y(n_1679)
);

INVx5_ASAP7_75t_L g1680 ( 
.A(n_1628),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1615),
.A2(n_817),
.B1(n_1404),
.B2(n_1446),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1624),
.A2(n_952),
.B1(n_1035),
.B2(n_971),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1582),
.B(n_1118),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1619),
.B(n_1514),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1619),
.B(n_1514),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1626),
.B(n_1414),
.Y(n_1687)
);

OAI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1590),
.A2(n_1494),
.B1(n_1419),
.B2(n_1035),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1616),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1550),
.Y(n_1690)
);

INVx8_ASAP7_75t_L g1691 ( 
.A(n_1628),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1626),
.B(n_1507),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1622),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1552),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1602),
.B(n_971),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1601),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1598),
.B(n_1507),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1534),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1635),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1680),
.Y(n_1700)
);

BUFx4f_ASAP7_75t_SL g1701 ( 
.A(n_1665),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1669),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1640),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1678),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1680),
.B(n_1628),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1650),
.B(n_1586),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1680),
.B(n_1627),
.Y(n_1707)
);

BUFx12f_ASAP7_75t_SL g1708 ( 
.A(n_1648),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1642),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1647),
.B(n_1586),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1641),
.B(n_1544),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1636),
.A2(n_1574),
.B(n_1456),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1677),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1684),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1634),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1677),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1697),
.B(n_1420),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1648),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1645),
.B(n_1088),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1648),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1691),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1697),
.B(n_1420),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1691),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1695),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1679),
.B(n_1108),
.Y(n_1726)
);

INVx6_ASAP7_75t_L g1727 ( 
.A(n_1691),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1656),
.A2(n_1561),
.B1(n_1196),
.B2(n_1176),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1649),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1690),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1649),
.Y(n_1731)
);

CKINVDCx6p67_ASAP7_75t_R g1732 ( 
.A(n_1634),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1694),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1634),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1651),
.B(n_1553),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1649),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1658),
.Y(n_1738)
);

INVx5_ASAP7_75t_L g1739 ( 
.A(n_1696),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1676),
.B(n_1419),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1654),
.B(n_1553),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1638),
.B(n_1627),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1725),
.A2(n_1662),
.B1(n_1667),
.B2(n_1661),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1702),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1720),
.B(n_1108),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1736),
.B(n_1741),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1726),
.B(n_1117),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1740),
.A2(n_1654),
.B(n_1670),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1715),
.B(n_1703),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1719),
.B(n_1687),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1713),
.B(n_1688),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1705),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1660),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_R g1755 ( 
.A(n_1701),
.B(n_1617),
.Y(n_1755)
);

AND2x2_ASAP7_75t_SL g1756 ( 
.A(n_1707),
.B(n_1633),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1704),
.Y(n_1757)
);

AOI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1740),
.A2(n_1676),
.B(n_1685),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1711),
.A2(n_1675),
.B1(n_1682),
.B2(n_1117),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1728),
.A2(n_1686),
.B1(n_1671),
.B2(n_1670),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1738),
.B(n_1605),
.C(n_1005),
.Y(n_1761)
);

NAND2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1739),
.B(n_1541),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1707),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1706),
.A2(n_1653),
.B(n_1655),
.C(n_1683),
.Y(n_1764)
);

OAI21xp33_ASAP7_75t_L g1765 ( 
.A1(n_1738),
.A2(n_955),
.B(n_934),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1714),
.A2(n_1671),
.B(n_1625),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1742),
.B(n_1644),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1709),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1718),
.A2(n_1659),
.B(n_1456),
.C(n_1580),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1730),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1742),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1714),
.A2(n_1674),
.B(n_1672),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1742),
.B(n_1672),
.Y(n_1773)
);

O2A1O1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1709),
.A2(n_1639),
.B(n_1408),
.C(n_1405),
.Y(n_1774)
);

BUFx4f_ASAP7_75t_SL g1775 ( 
.A(n_1722),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1733),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1717),
.A2(n_1692),
.B(n_1664),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1739),
.B(n_1673),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1718),
.A2(n_1462),
.B(n_982),
.C(n_1021),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1723),
.A2(n_1135),
.B1(n_1147),
.B2(n_1142),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1716),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1707),
.B(n_1663),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1735),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1717),
.A2(n_1692),
.B(n_1668),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_SL g1785 ( 
.A(n_1739),
.B(n_1584),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1735),
.B(n_1666),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1731),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1743),
.A2(n_1646),
.B1(n_1723),
.B2(n_1595),
.Y(n_1788)
);

AND2x2_ASAP7_75t_SL g1789 ( 
.A(n_1756),
.B(n_1618),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1771),
.B(n_1752),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1753),
.B(n_1721),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1748),
.B(n_1677),
.Y(n_1793)
);

INVx8_ASAP7_75t_L g1794 ( 
.A(n_1763),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1749),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1768),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_SL g1797 ( 
.A1(n_1751),
.A2(n_1646),
.B(n_1724),
.C(n_1558),
.Y(n_1797)
);

INVx2_ASAP7_75t_SL g1798 ( 
.A(n_1783),
.Y(n_1798)
);

AO22x1_ASAP7_75t_L g1799 ( 
.A1(n_1745),
.A2(n_1364),
.B1(n_1095),
.B2(n_1157),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1770),
.Y(n_1800)
);

CKINVDCx11_ASAP7_75t_R g1801 ( 
.A(n_1763),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1739),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1763),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1744),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1776),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1781),
.Y(n_1806)
);

BUFx8_ASAP7_75t_L g1807 ( 
.A(n_1755),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1775),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1750),
.B(n_1739),
.Y(n_1809)
);

INVx4_ASAP7_75t_L g1810 ( 
.A(n_1787),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1759),
.A2(n_1135),
.B1(n_1147),
.B2(n_1142),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1780),
.A2(n_1404),
.B1(n_1323),
.B2(n_1259),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1769),
.A2(n_1681),
.B(n_1193),
.C(n_1144),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1750),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1760),
.A2(n_1631),
.B1(n_1554),
.B2(n_1562),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1787),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1767),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1782),
.A2(n_1404),
.B1(n_1259),
.B2(n_1637),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1750),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1773),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1772),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1765),
.B(n_1576),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1786),
.B(n_1732),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1784),
.A2(n_1734),
.B(n_1542),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1758),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1762),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1762),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1778),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1746),
.B(n_1731),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1754),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1760),
.A2(n_1652),
.B1(n_1657),
.B2(n_1643),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_1747),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1777),
.B(n_1677),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1785),
.Y(n_1834)
);

BUFx12f_ASAP7_75t_L g1835 ( 
.A(n_1761),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1764),
.B(n_1732),
.Y(n_1836)
);

BUFx8_ASAP7_75t_L g1837 ( 
.A(n_1785),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1796),
.Y(n_1838)
);

BUFx12f_ASAP7_75t_L g1839 ( 
.A(n_1807),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_SL g1840 ( 
.A1(n_1813),
.A2(n_1779),
.B(n_955),
.C(n_1021),
.Y(n_1840)
);

NAND2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1808),
.B(n_1731),
.Y(n_1841)
);

AO31x2_ASAP7_75t_L g1842 ( 
.A1(n_1825),
.A2(n_1734),
.A3(n_1766),
.B(n_1542),
.Y(n_1842)
);

AOI31xp67_ASAP7_75t_L g1843 ( 
.A1(n_1833),
.A2(n_1271),
.A3(n_1272),
.B(n_1270),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1824),
.A2(n_1710),
.B(n_1700),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1792),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1800),
.Y(n_1846)
);

AO31x2_ASAP7_75t_L g1847 ( 
.A1(n_1788),
.A2(n_1535),
.A3(n_1479),
.B(n_1474),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1807),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1795),
.B(n_1677),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1795),
.B(n_1729),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_SL g1851 ( 
.A1(n_1815),
.A2(n_982),
.B(n_1774),
.C(n_972),
.Y(n_1851)
);

NAND2x1p5_ASAP7_75t_L g1852 ( 
.A(n_1834),
.B(n_1731),
.Y(n_1852)
);

AO32x2_ASAP7_75t_L g1853 ( 
.A1(n_1788),
.A2(n_1737),
.A3(n_1708),
.B1(n_1295),
.B2(n_1255),
.Y(n_1853)
);

O2A1O1Ixp33_ASAP7_75t_SL g1854 ( 
.A1(n_1815),
.A2(n_975),
.B(n_1015),
.C(n_900),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1804),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1811),
.A2(n_1708),
.B1(n_1613),
.B2(n_1598),
.Y(n_1856)
);

AO32x2_ASAP7_75t_L g1857 ( 
.A1(n_1810),
.A2(n_1737),
.A3(n_1295),
.B1(n_1326),
.B2(n_1578),
.Y(n_1857)
);

O2A1O1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1797),
.A2(n_850),
.B(n_843),
.C(n_852),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1824),
.A2(n_1710),
.B(n_1700),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1805),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1789),
.A2(n_1095),
.B1(n_1157),
.B2(n_1190),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1822),
.A2(n_856),
.B(n_861),
.C(n_855),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1812),
.A2(n_1724),
.B1(n_1727),
.B2(n_1729),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1803),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1833),
.A2(n_1710),
.B(n_1700),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1793),
.A2(n_1821),
.B(n_1809),
.Y(n_1866)
);

BUFx8_ASAP7_75t_L g1867 ( 
.A(n_1835),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1806),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1793),
.A2(n_1724),
.B(n_1729),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1817),
.Y(n_1870)
);

A2O1A1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1811),
.A2(n_866),
.B(n_867),
.C(n_863),
.Y(n_1871)
);

AO31x2_ASAP7_75t_L g1872 ( 
.A1(n_1830),
.A2(n_1479),
.A3(n_1474),
.B(n_1698),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1836),
.A2(n_1151),
.B(n_953),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1790),
.B(n_951),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1809),
.A2(n_1705),
.B(n_1731),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1829),
.A2(n_956),
.B(n_954),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1829),
.A2(n_1705),
.B(n_1495),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1832),
.A2(n_1823),
.B(n_1834),
.C(n_1629),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1814),
.A2(n_1598),
.B1(n_1613),
.B2(n_1226),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1828),
.B(n_1722),
.Y(n_1880)
);

AO31x2_ASAP7_75t_L g1881 ( 
.A1(n_1827),
.A2(n_1693),
.A3(n_1689),
.B(n_1594),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1798),
.A2(n_1014),
.B(n_1018),
.C(n_989),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1820),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1814),
.B(n_957),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1819),
.Y(n_1885)
);

NAND3x1_ASAP7_75t_L g1886 ( 
.A(n_1799),
.B(n_842),
.C(n_841),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1819),
.Y(n_1887)
);

AOI31xp67_ASAP7_75t_L g1888 ( 
.A1(n_1791),
.A2(n_1280),
.A3(n_1284),
.B(n_1275),
.Y(n_1888)
);

NAND2x1p5_ASAP7_75t_L g1889 ( 
.A(n_1834),
.B(n_1722),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1831),
.A2(n_1816),
.B(n_959),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1801),
.Y(n_1891)
);

O2A1O1Ixp33_ASAP7_75t_SL g1892 ( 
.A1(n_1816),
.A2(n_1020),
.B(n_978),
.C(n_983),
.Y(n_1892)
);

AOI31xp67_ASAP7_75t_L g1893 ( 
.A1(n_1791),
.A2(n_1291),
.A3(n_1292),
.B(n_1288),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_SL g1894 ( 
.A1(n_1837),
.A2(n_984),
.B(n_987),
.C(n_977),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1818),
.A2(n_960),
.B(n_961),
.C(n_958),
.Y(n_1895)
);

A2O1A1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1828),
.A2(n_965),
.B(n_966),
.C(n_962),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_SL g1897 ( 
.A1(n_1837),
.A2(n_994),
.B(n_995),
.C(n_990),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1828),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1802),
.A2(n_1810),
.B(n_1827),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1802),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1803),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1794),
.A2(n_1029),
.B(n_1028),
.Y(n_1902)
);

AO31x2_ASAP7_75t_L g1903 ( 
.A1(n_1826),
.A2(n_1480),
.A3(n_1581),
.B(n_1568),
.Y(n_1903)
);

O2A1O1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1794),
.A2(n_1034),
.B(n_1033),
.C(n_1158),
.Y(n_1904)
);

OAI222xp33_ASAP7_75t_L g1905 ( 
.A1(n_1794),
.A2(n_1037),
.B1(n_1203),
.B2(n_1581),
.C1(n_1568),
.C2(n_1143),
.Y(n_1905)
);

O2A1O1Ixp33_ASAP7_75t_SL g1906 ( 
.A1(n_1803),
.A2(n_999),
.B(n_1001),
.C(n_996),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1826),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1826),
.B(n_1722),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1885),
.B(n_1150),
.Y(n_1909)
);

CKINVDCx6p67_ASAP7_75t_R g1910 ( 
.A(n_1839),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1854),
.A2(n_1598),
.B1(n_1613),
.B2(n_1596),
.Y(n_1911)
);

OAI211xp5_ASAP7_75t_L g1912 ( 
.A1(n_1851),
.A2(n_1472),
.B(n_827),
.C(n_828),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1873),
.A2(n_1876),
.B1(n_1472),
.B2(n_1874),
.Y(n_1913)
);

OAI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1840),
.A2(n_824),
.B1(n_1226),
.B2(n_1171),
.C(n_1167),
.Y(n_1914)
);

AO21x2_ASAP7_75t_L g1915 ( 
.A1(n_1866),
.A2(n_1495),
.B(n_1274),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1855),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1883),
.A2(n_1613),
.B1(n_1445),
.B2(n_1575),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1856),
.A2(n_1546),
.B1(n_1577),
.B2(n_1468),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1878),
.A2(n_1727),
.B1(n_1098),
.B2(n_1530),
.Y(n_1919)
);

NOR2xp67_ASAP7_75t_L g1920 ( 
.A(n_1899),
.B(n_1865),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1853),
.A2(n_1163),
.B1(n_1727),
.B2(n_1469),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1845),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1861),
.A2(n_1468),
.B1(n_1349),
.B2(n_1342),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1860),
.A2(n_1100),
.B1(n_1143),
.B2(n_1000),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1877),
.A2(n_1556),
.B(n_1540),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1898),
.A2(n_1468),
.B1(n_1290),
.B2(n_1297),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_SL g1927 ( 
.A1(n_1853),
.A2(n_1469),
.B1(n_1506),
.B2(n_1484),
.Y(n_1927)
);

OAI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1879),
.A2(n_1541),
.B1(n_1548),
.B2(n_1543),
.Y(n_1928)
);

INVx3_ASAP7_75t_SL g1929 ( 
.A(n_1891),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1887),
.A2(n_1303),
.B1(n_1310),
.B2(n_1279),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1890),
.A2(n_1506),
.B1(n_1484),
.B2(n_611),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1870),
.A2(n_1315),
.B1(n_1317),
.B2(n_1314),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1900),
.A2(n_1329),
.B1(n_1331),
.B2(n_1320),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1838),
.B(n_1),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1906),
.A2(n_1596),
.B1(n_1492),
.B2(n_1524),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1907),
.A2(n_1346),
.B1(n_1347),
.B2(n_1336),
.Y(n_1936)
);

INVx4_ASAP7_75t_L g1937 ( 
.A(n_1901),
.Y(n_1937)
);

CKINVDCx8_ASAP7_75t_R g1938 ( 
.A(n_1901),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1868),
.B(n_1150),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1850),
.B(n_5),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1849),
.A2(n_1848),
.B1(n_1846),
.B2(n_1863),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1864),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1884),
.B(n_1168),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1869),
.B(n_1168),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1880),
.A2(n_1556),
.B(n_1540),
.Y(n_1945)
);

OAI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1875),
.A2(n_1548),
.B1(n_1543),
.B2(n_1620),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1881),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1881),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1842),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1842),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1902),
.A2(n_1350),
.B1(n_1351),
.B2(n_1348),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1903),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1858),
.A2(n_846),
.B1(n_1006),
.B2(n_1010),
.C(n_1004),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1903),
.Y(n_1954)
);

INVx4_ASAP7_75t_L g1955 ( 
.A(n_1841),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1867),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1886),
.A2(n_1543),
.B1(n_1548),
.B2(n_1614),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1889),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1921),
.A2(n_1871),
.B(n_1882),
.C(n_1862),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1947),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1934),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1922),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1937),
.Y(n_1963)
);

OA21x2_ASAP7_75t_L g1964 ( 
.A1(n_1950),
.A2(n_1949),
.B(n_1948),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1952),
.A2(n_1859),
.B(n_1844),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1937),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1909),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1909),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1954),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1916),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1939),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1939),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1944),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1944),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1910),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1940),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1941),
.Y(n_1977)
);

OAI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1920),
.A2(n_1852),
.B(n_1908),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1915),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1915),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1942),
.B(n_1847),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1920),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1943),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1919),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1925),
.A2(n_1904),
.B(n_1843),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1958),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1946),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1929),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1984),
.A2(n_1913),
.B1(n_1938),
.B2(n_1911),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1983),
.B(n_1847),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1983),
.A2(n_1931),
.B1(n_1957),
.B2(n_1918),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1971),
.A2(n_1917),
.B1(n_1911),
.B2(n_1924),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_SL g1993 ( 
.A1(n_1977),
.A2(n_1987),
.B1(n_1976),
.B2(n_1981),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1971),
.A2(n_1923),
.B1(n_1927),
.B2(n_1932),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1971),
.Y(n_1995)
);

NAND3xp33_ASAP7_75t_L g1996 ( 
.A(n_1977),
.B(n_1912),
.C(n_1892),
.Y(n_1996)
);

AOI221xp5_ASAP7_75t_L g1997 ( 
.A1(n_1976),
.A2(n_1897),
.B1(n_1894),
.B2(n_1914),
.C(n_1953),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1972),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1972),
.Y(n_1999)
);

OAI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1959),
.A2(n_1935),
.B1(n_1930),
.B2(n_1933),
.C(n_1951),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1975),
.Y(n_2001)
);

AOI221xp5_ASAP7_75t_L g2002 ( 
.A1(n_1982),
.A2(n_1972),
.B1(n_1980),
.B2(n_1979),
.C(n_1967),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1962),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1961),
.A2(n_1955),
.B1(n_1956),
.B2(n_1935),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_L g2005 ( 
.A1(n_1982),
.A2(n_1945),
.B(n_1936),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1962),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1967),
.A2(n_1928),
.B1(n_1926),
.B2(n_1955),
.Y(n_2007)
);

OA21x2_ASAP7_75t_L g2008 ( 
.A1(n_1969),
.A2(n_1896),
.B(n_1905),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_SL g2009 ( 
.A(n_1987),
.B(n_1895),
.C(n_1857),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1968),
.A2(n_1201),
.B1(n_1184),
.B2(n_557),
.Y(n_2010)
);

OR2x6_ASAP7_75t_L g2011 ( 
.A(n_1985),
.B(n_1888),
.Y(n_2011)
);

OAI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1978),
.A2(n_1893),
.B(n_1012),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1973),
.A2(n_1461),
.B1(n_1475),
.B2(n_1473),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_2008),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_2003),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_2001),
.B(n_1963),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2006),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_2001),
.B(n_1963),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1990),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_2008),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1995),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1998),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1999),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_2011),
.B(n_2005),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2001),
.B(n_1966),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1993),
.B(n_1966),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2010),
.Y(n_2027)
);

AND2x6_ASAP7_75t_SL g2028 ( 
.A(n_1996),
.B(n_1975),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_2011),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2004),
.B(n_1988),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2010),
.Y(n_2031)
);

BUFx3_ASAP7_75t_L g2032 ( 
.A(n_1996),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2011),
.B(n_1988),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1989),
.Y(n_2034)
);

INVxp67_ASAP7_75t_L g2035 ( 
.A(n_2009),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2002),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2012),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2000),
.B(n_1975),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1992),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2007),
.B(n_1986),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1991),
.B(n_1986),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1997),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1994),
.B(n_1973),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_2013),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_2001),
.Y(n_2045)
);

OAI31xp33_ASAP7_75t_L g2046 ( 
.A1(n_2032),
.A2(n_1980),
.A3(n_1979),
.B(n_1974),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_2029),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_2015),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_2032),
.B(n_1974),
.C(n_1969),
.Y(n_2049)
);

OAI211xp5_ASAP7_75t_L g2050 ( 
.A1(n_2032),
.A2(n_1978),
.B(n_1985),
.C(n_1969),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_L g2051 ( 
.A(n_2035),
.B(n_1965),
.C(n_1013),
.Y(n_2051)
);

OAI222xp33_ASAP7_75t_L g2052 ( 
.A1(n_2036),
.A2(n_1970),
.B1(n_1960),
.B2(n_1964),
.C1(n_1857),
.C2(n_1965),
.Y(n_2052)
);

OAI221xp5_ASAP7_75t_L g2053 ( 
.A1(n_2036),
.A2(n_1970),
.B1(n_1960),
.B2(n_1964),
.C(n_1017),
.Y(n_2053)
);

NAND4xp25_ASAP7_75t_L g2054 ( 
.A(n_2038),
.B(n_1016),
.C(n_1019),
.D(n_1011),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2038),
.B(n_1022),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_2045),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_2045),
.B(n_1162),
.Y(n_2057)
);

BUFx2_ASAP7_75t_L g2058 ( 
.A(n_2030),
.Y(n_2058)
);

AOI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_2042),
.A2(n_825),
.B1(n_794),
.B2(n_789),
.C(n_1179),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2017),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2017),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2026),
.A2(n_1964),
.B1(n_1632),
.B2(n_1614),
.Y(n_2062)
);

NAND3xp33_ASAP7_75t_L g2063 ( 
.A(n_2042),
.B(n_1964),
.C(n_611),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2027),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2027),
.Y(n_2065)
);

AO21x2_ASAP7_75t_L g2066 ( 
.A1(n_2029),
.A2(n_1181),
.B(n_1180),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2031),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_2058),
.B(n_2034),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2056),
.B(n_2033),
.Y(n_2069)
);

NAND2x1p5_ASAP7_75t_L g2070 ( 
.A(n_2057),
.B(n_2016),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2056),
.B(n_2033),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2066),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_2048),
.B(n_2034),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2060),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2064),
.B(n_2026),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_2056),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2057),
.B(n_2016),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2061),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2065),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2067),
.B(n_2030),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2062),
.B(n_2018),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_2055),
.Y(n_2082)
);

INVx4_ASAP7_75t_L g2083 ( 
.A(n_2066),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_2068),
.B(n_2024),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2077),
.B(n_2018),
.Y(n_2085)
);

OAI321xp33_ASAP7_75t_L g2086 ( 
.A1(n_2075),
.A2(n_2050),
.A3(n_2063),
.B1(n_2042),
.B2(n_2020),
.C(n_2014),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2070),
.Y(n_2087)
);

INVxp67_ASAP7_75t_L g2088 ( 
.A(n_2069),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2073),
.B(n_2029),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_2082),
.B(n_2024),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2077),
.B(n_2025),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2080),
.B(n_2037),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2088),
.B(n_2082),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2085),
.B(n_2070),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2091),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2092),
.B(n_2079),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2089),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2087),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_2086),
.B(n_2076),
.Y(n_2099)
);

NAND3x1_ASAP7_75t_L g2100 ( 
.A(n_2093),
.B(n_2076),
.C(n_2071),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2097),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2099),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2095),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2098),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2103),
.B(n_2094),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_2102),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2102),
.B(n_2096),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2105),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2106),
.B(n_2069),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2109),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2108),
.B(n_2107),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_2111),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_2110),
.B(n_2090),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2112),
.Y(n_2114)
);

XOR2xp5_ASAP7_75t_L g2115 ( 
.A(n_2113),
.B(n_2101),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2112),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2114),
.B(n_2071),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2115),
.Y(n_2118)
);

AOI211xp5_ASAP7_75t_L g2119 ( 
.A1(n_2116),
.A2(n_2104),
.B(n_2084),
.C(n_2086),
.Y(n_2119)
);

AOI21xp33_ASAP7_75t_L g2120 ( 
.A1(n_2115),
.A2(n_2100),
.B(n_2083),
.Y(n_2120)
);

NAND4xp75_ASAP7_75t_L g2121 ( 
.A(n_2118),
.B(n_2117),
.C(n_2120),
.D(n_2119),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2118),
.A2(n_2054),
.B(n_2076),
.C(n_2074),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2117),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2123),
.A2(n_2083),
.B1(n_2047),
.B2(n_2072),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2122),
.Y(n_2125)
);

AOI322xp5_ASAP7_75t_L g2126 ( 
.A1(n_2121),
.A2(n_2051),
.A3(n_2072),
.B1(n_2020),
.B2(n_2014),
.C1(n_2078),
.C2(n_2024),
.Y(n_2126)
);

CKINVDCx20_ASAP7_75t_R g2127 ( 
.A(n_2123),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_2123),
.A2(n_2083),
.B1(n_2081),
.B2(n_2024),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2123),
.A2(n_2081),
.B1(n_2020),
.B2(n_2014),
.Y(n_2129)
);

INVx2_ASAP7_75t_SL g2130 ( 
.A(n_2123),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2123),
.B(n_2025),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2123),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2123),
.Y(n_2133)
);

BUFx2_ASAP7_75t_L g2134 ( 
.A(n_2123),
.Y(n_2134)
);

NAND4xp75_ASAP7_75t_L g2135 ( 
.A(n_2121),
.B(n_2059),
.C(n_2046),
.D(n_1194),
.Y(n_2135)
);

O2A1O1Ixp5_ASAP7_75t_L g2136 ( 
.A1(n_2123),
.A2(n_2052),
.B(n_2049),
.C(n_2028),
.Y(n_2136)
);

NAND3xp33_ASAP7_75t_L g2137 ( 
.A(n_2134),
.B(n_1217),
.C(n_1195),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2131),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2130),
.B(n_2039),
.Y(n_2139)
);

NAND3xp33_ASAP7_75t_SL g2140 ( 
.A(n_2127),
.B(n_2063),
.C(n_1197),
.Y(n_2140)
);

AND4x1_ASAP7_75t_L g2141 ( 
.A(n_2132),
.B(n_1207),
.C(n_1209),
.D(n_1192),
.Y(n_2141)
);

NOR3xp33_ASAP7_75t_L g2142 ( 
.A(n_2133),
.B(n_1225),
.C(n_1220),
.Y(n_2142)
);

NOR4xp25_ASAP7_75t_L g2143 ( 
.A(n_2125),
.B(n_2039),
.C(n_2019),
.D(n_1186),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_2131),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2135),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2129),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2126),
.B(n_2041),
.Y(n_2147)
);

NAND4xp75_ASAP7_75t_L g2148 ( 
.A(n_2136),
.B(n_2037),
.C(n_2031),
.D(n_1298),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2128),
.B(n_2041),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2124),
.B(n_2019),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2134),
.B(n_2040),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2134),
.B(n_2040),
.Y(n_2152)
);

NOR2x1p5_ASAP7_75t_L g2153 ( 
.A(n_2132),
.B(n_1573),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2134),
.B(n_2043),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2134),
.Y(n_2155)
);

NOR2x1_ASAP7_75t_L g2156 ( 
.A(n_2127),
.B(n_1186),
.Y(n_2156)
);

NOR2xp67_ASAP7_75t_L g2157 ( 
.A(n_2130),
.B(n_6),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2134),
.Y(n_2158)
);

NAND4xp75_ASAP7_75t_L g2159 ( 
.A(n_2130),
.B(n_1304),
.C(n_1268),
.D(n_2043),
.Y(n_2159)
);

NOR2x1_ASAP7_75t_L g2160 ( 
.A(n_2127),
.B(n_1201),
.Y(n_2160)
);

NAND3xp33_ASAP7_75t_SL g2161 ( 
.A(n_2127),
.B(n_2053),
.C(n_1264),
.Y(n_2161)
);

NOR2x1_ASAP7_75t_L g2162 ( 
.A(n_2127),
.B(n_1217),
.Y(n_2162)
);

NOR3xp33_ASAP7_75t_SL g2163 ( 
.A(n_2132),
.B(n_7),
.C(n_9),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2134),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2134),
.B(n_2021),
.Y(n_2165)
);

NAND4xp75_ASAP7_75t_L g2166 ( 
.A(n_2130),
.B(n_1304),
.C(n_1276),
.D(n_1263),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2134),
.Y(n_2167)
);

O2A1O1Ixp33_ASAP7_75t_L g2168 ( 
.A1(n_2130),
.A2(n_1091),
.B(n_1092),
.C(n_1085),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_L g2169 ( 
.A(n_2134),
.B(n_1217),
.C(n_1092),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2134),
.Y(n_2170)
);

INVxp33_ASAP7_75t_SL g2171 ( 
.A(n_2134),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2134),
.B(n_2021),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_SL g2173 ( 
.A(n_2127),
.B(n_1091),
.C(n_1623),
.Y(n_2173)
);

NAND4xp75_ASAP7_75t_L g2174 ( 
.A(n_2130),
.B(n_2022),
.C(n_2023),
.D(n_1392),
.Y(n_2174)
);

NAND3xp33_ASAP7_75t_SL g2175 ( 
.A(n_2127),
.B(n_532),
.C(n_528),
.Y(n_2175)
);

NAND3xp33_ASAP7_75t_L g2176 ( 
.A(n_2134),
.B(n_537),
.C(n_534),
.Y(n_2176)
);

NAND3xp33_ASAP7_75t_L g2177 ( 
.A(n_2134),
.B(n_546),
.C(n_538),
.Y(n_2177)
);

NOR4xp25_ASAP7_75t_L g2178 ( 
.A(n_2130),
.B(n_2022),
.C(n_2023),
.D(n_1432),
.Y(n_2178)
);

NOR3xp33_ASAP7_75t_L g2179 ( 
.A(n_2134),
.B(n_887),
.C(n_1250),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2134),
.B(n_2044),
.Y(n_2180)
);

AOI221xp5_ASAP7_75t_L g2181 ( 
.A1(n_2171),
.A2(n_2044),
.B1(n_1578),
.B2(n_1573),
.C(n_562),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2154),
.Y(n_2182)
);

AOI221x1_ASAP7_75t_SL g2183 ( 
.A1(n_2155),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_SL g2184 ( 
.A1(n_2158),
.A2(n_2044),
.B1(n_15),
.B2(n_13),
.Y(n_2184)
);

NAND3x1_ASAP7_75t_SL g2185 ( 
.A(n_2156),
.B(n_13),
.C(n_14),
.Y(n_2185)
);

OAI211xp5_ASAP7_75t_SL g2186 ( 
.A1(n_2164),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2167),
.A2(n_549),
.B(n_548),
.Y(n_2187)
);

OAI311xp33_ASAP7_75t_L g2188 ( 
.A1(n_2151),
.A2(n_1306),
.A3(n_1322),
.B1(n_1294),
.C1(n_1250),
.Y(n_2188)
);

OAI211xp5_ASAP7_75t_L g2189 ( 
.A1(n_2170),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_2189)
);

AOI211x1_ASAP7_75t_SL g2190 ( 
.A1(n_2147),
.A2(n_24),
.B(n_20),
.C(n_23),
.Y(n_2190)
);

NAND4xp25_ASAP7_75t_L g2191 ( 
.A(n_2152),
.B(n_26),
.C(n_23),
.D(n_25),
.Y(n_2191)
);

OA22x2_ASAP7_75t_L g2192 ( 
.A1(n_2144),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_2192)
);

OAI211xp5_ASAP7_75t_SL g2193 ( 
.A1(n_2146),
.A2(n_31),
.B(n_27),
.C(n_30),
.Y(n_2193)
);

OAI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2138),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.C(n_35),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2180),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2157),
.B(n_1492),
.Y(n_2196)
);

NAND4xp25_ASAP7_75t_L g2197 ( 
.A(n_2139),
.B(n_37),
.C(n_34),
.D(n_36),
.Y(n_2197)
);

XOR2xp5_ASAP7_75t_L g2198 ( 
.A(n_2173),
.B(n_38),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2163),
.B(n_38),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_2165),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2145),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_2201)
);

AO22x2_ASAP7_75t_L g2202 ( 
.A1(n_2175),
.A2(n_43),
.B1(n_39),
.B2(n_42),
.Y(n_2202)
);

OAI21xp33_ASAP7_75t_L g2203 ( 
.A1(n_2149),
.A2(n_568),
.B(n_567),
.Y(n_2203)
);

AOI211xp5_ASAP7_75t_L g2204 ( 
.A1(n_2176),
.A2(n_48),
.B(n_45),
.C(n_46),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2165),
.B(n_49),
.Y(n_2205)
);

A2O1A1Ixp33_ASAP7_75t_L g2206 ( 
.A1(n_2150),
.A2(n_2177),
.B(n_2172),
.C(n_2168),
.Y(n_2206)
);

NAND3xp33_ASAP7_75t_SL g2207 ( 
.A(n_2179),
.B(n_574),
.C(n_573),
.Y(n_2207)
);

AOI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2148),
.A2(n_1492),
.B1(n_1524),
.B2(n_1306),
.Y(n_2208)
);

OAI321xp33_ASAP7_75t_L g2209 ( 
.A1(n_2137),
.A2(n_2140),
.A3(n_2169),
.B1(n_2141),
.B2(n_2143),
.C(n_2153),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2160),
.B(n_49),
.Y(n_2210)
);

AOI211x1_ASAP7_75t_L g2211 ( 
.A1(n_2159),
.A2(n_54),
.B(n_50),
.C(n_53),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2142),
.B(n_55),
.Y(n_2212)
);

OA22x2_ASAP7_75t_L g2213 ( 
.A1(n_2166),
.A2(n_60),
.B1(n_55),
.B2(n_56),
.Y(n_2213)
);

AO22x2_ASAP7_75t_L g2214 ( 
.A1(n_2174),
.A2(n_64),
.B1(n_56),
.B2(n_63),
.Y(n_2214)
);

CKINVDCx20_ASAP7_75t_R g2215 ( 
.A(n_2161),
.Y(n_2215)
);

OA22x2_ASAP7_75t_L g2216 ( 
.A1(n_2178),
.A2(n_66),
.B1(n_63),
.B2(n_65),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2162),
.Y(n_2217)
);

O2A1O1Ixp33_ASAP7_75t_L g2218 ( 
.A1(n_2171),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_2218)
);

AOI211x1_ASAP7_75t_L g2219 ( 
.A1(n_2155),
.A2(n_73),
.B(n_69),
.C(n_70),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2155),
.Y(n_2220)
);

NOR3xp33_ASAP7_75t_L g2221 ( 
.A(n_2155),
.B(n_1322),
.C(n_1294),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2171),
.B(n_1492),
.Y(n_2222)
);

OAI221xp5_ASAP7_75t_L g2223 ( 
.A1(n_2155),
.A2(n_74),
.B1(n_69),
.B2(n_73),
.C(n_76),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2171),
.A2(n_1524),
.B1(n_577),
.B2(n_578),
.Y(n_2224)
);

OA22x2_ASAP7_75t_L g2225 ( 
.A1(n_2155),
.A2(n_78),
.B1(n_74),
.B2(n_77),
.Y(n_2225)
);

BUFx10_ASAP7_75t_L g2226 ( 
.A(n_2155),
.Y(n_2226)
);

NAND3xp33_ASAP7_75t_SL g2227 ( 
.A(n_2155),
.B(n_582),
.C(n_576),
.Y(n_2227)
);

AOI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2171),
.A2(n_594),
.B1(n_598),
.B2(n_596),
.C(n_592),
.Y(n_2228)
);

OAI21x1_ASAP7_75t_SL g2229 ( 
.A1(n_2151),
.A2(n_78),
.B(n_79),
.Y(n_2229)
);

NOR2x1_ASAP7_75t_L g2230 ( 
.A(n_2155),
.B(n_79),
.Y(n_2230)
);

AO22x1_ASAP7_75t_L g2231 ( 
.A1(n_2171),
.A2(n_1524),
.B1(n_83),
.B2(n_80),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2154),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2171),
.A2(n_601),
.B1(n_604),
.B2(n_600),
.Y(n_2233)
);

AOI221xp5_ASAP7_75t_L g2234 ( 
.A1(n_2171),
.A2(n_616),
.B1(n_621),
.B2(n_612),
.C(n_609),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2171),
.B(n_80),
.Y(n_2235)
);

AOI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_2171),
.A2(n_626),
.B(n_625),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2171),
.B(n_81),
.Y(n_2237)
);

A2O1A1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_2155),
.A2(n_632),
.B(n_636),
.C(n_630),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2154),
.Y(n_2239)
);

OAI22xp33_ASAP7_75t_SL g2240 ( 
.A1(n_2171),
.A2(n_642),
.B1(n_645),
.B2(n_637),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_SL g2241 ( 
.A(n_2155),
.B(n_652),
.C(n_649),
.Y(n_2241)
);

A2O1A1Ixp33_ASAP7_75t_L g2242 ( 
.A1(n_2155),
.A2(n_660),
.B(n_661),
.C(n_659),
.Y(n_2242)
);

NAND4xp75_ASAP7_75t_L g2243 ( 
.A(n_2155),
.B(n_87),
.C(n_81),
.D(n_85),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2171),
.A2(n_666),
.B1(n_667),
.B2(n_665),
.Y(n_2244)
);

AOI221xp5_ASAP7_75t_L g2245 ( 
.A1(n_2171),
.A2(n_716),
.B1(n_751),
.B2(n_750),
.C(n_748),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_SL g2246 ( 
.A(n_2155),
.B(n_671),
.C(n_669),
.Y(n_2246)
);

AOI211xp5_ASAP7_75t_L g2247 ( 
.A1(n_2155),
.A2(n_91),
.B(n_85),
.C(n_88),
.Y(n_2247)
);

OAI322xp33_ASAP7_75t_L g2248 ( 
.A1(n_2155),
.A2(n_91),
.A3(n_92),
.B1(n_93),
.B2(n_94),
.C1(n_97),
.C2(n_98),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_2171),
.B(n_92),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_2200),
.B(n_2220),
.Y(n_2250)
);

NOR3xp33_ASAP7_75t_L g2251 ( 
.A(n_2182),
.B(n_674),
.C(n_672),
.Y(n_2251)
);

NOR3xp33_ASAP7_75t_L g2252 ( 
.A(n_2232),
.B(n_683),
.C(n_682),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2235),
.A2(n_692),
.B1(n_694),
.B2(n_689),
.Y(n_2253)
);

NAND3x1_ASAP7_75t_SL g2254 ( 
.A(n_2230),
.B(n_93),
.C(n_97),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2205),
.B(n_99),
.Y(n_2255)
);

NOR4xp25_ASAP7_75t_SL g2256 ( 
.A(n_2239),
.B(n_101),
.C(n_99),
.D(n_100),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2226),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2192),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2197),
.B(n_100),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2191),
.B(n_2237),
.Y(n_2260)
);

NOR2x1_ASAP7_75t_L g2261 ( 
.A(n_2195),
.B(n_2243),
.Y(n_2261)
);

NOR2x1_ASAP7_75t_L g2262 ( 
.A(n_2205),
.B(n_102),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2199),
.B(n_102),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2190),
.B(n_103),
.Y(n_2264)
);

INVxp67_ASAP7_75t_SL g2265 ( 
.A(n_2249),
.Y(n_2265)
);

OAI211xp5_ASAP7_75t_L g2266 ( 
.A1(n_2219),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_2266)
);

AND3x4_ASAP7_75t_L g2267 ( 
.A(n_2221),
.B(n_104),
.C(n_105),
.Y(n_2267)
);

INVxp67_ASAP7_75t_L g2268 ( 
.A(n_2229),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2186),
.B(n_106),
.Y(n_2269)
);

AND3x2_ASAP7_75t_L g2270 ( 
.A(n_2247),
.B(n_106),
.C(n_108),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2198),
.B(n_108),
.Y(n_2271)
);

NAND4xp75_ASAP7_75t_L g2272 ( 
.A(n_2211),
.B(n_2187),
.C(n_2236),
.D(n_2212),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_L g2273 ( 
.A(n_2228),
.B(n_611),
.C(n_570),
.Y(n_2273)
);

NAND4xp25_ASAP7_75t_L g2274 ( 
.A(n_2183),
.B(n_111),
.C(n_109),
.D(n_110),
.Y(n_2274)
);

NOR2x1p5_ASAP7_75t_L g2275 ( 
.A(n_2222),
.B(n_109),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2225),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2206),
.B(n_111),
.Y(n_2277)
);

XOR2x1_ASAP7_75t_L g2278 ( 
.A(n_2244),
.B(n_112),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2210),
.B(n_114),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2202),
.B(n_115),
.Y(n_2280)
);

NOR2x1_ASAP7_75t_L g2281 ( 
.A(n_2227),
.B(n_116),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2214),
.Y(n_2282)
);

NAND2x1p5_ASAP7_75t_L g2283 ( 
.A(n_2217),
.B(n_1523),
.Y(n_2283)
);

AND3x4_ASAP7_75t_L g2284 ( 
.A(n_2185),
.B(n_116),
.C(n_117),
.Y(n_2284)
);

NOR2xp67_ASAP7_75t_L g2285 ( 
.A(n_2189),
.B(n_117),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_2215),
.Y(n_2286)
);

AOI221xp5_ASAP7_75t_L g2287 ( 
.A1(n_2240),
.A2(n_712),
.B1(n_715),
.B2(n_711),
.C(n_709),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2193),
.B(n_118),
.Y(n_2288)
);

NOR3xp33_ASAP7_75t_L g2289 ( 
.A(n_2241),
.B(n_696),
.C(n_695),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2202),
.B(n_118),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2214),
.Y(n_2291)
);

NOR3xp33_ASAP7_75t_SL g2292 ( 
.A(n_2246),
.B(n_721),
.C(n_699),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2216),
.B(n_119),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2184),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2196),
.B(n_120),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_2203),
.Y(n_2296)
);

NAND3xp33_ASAP7_75t_L g2297 ( 
.A(n_2234),
.B(n_611),
.C(n_570),
.Y(n_2297)
);

NOR2x1_ASAP7_75t_L g2298 ( 
.A(n_2238),
.B(n_121),
.Y(n_2298)
);

XNOR2xp5_ASAP7_75t_L g2299 ( 
.A(n_2213),
.B(n_2208),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_2242),
.B(n_122),
.Y(n_2300)
);

NOR2x1_ASAP7_75t_L g2301 ( 
.A(n_2248),
.B(n_123),
.Y(n_2301)
);

NOR3xp33_ASAP7_75t_L g2302 ( 
.A(n_2207),
.B(n_726),
.C(n_724),
.Y(n_2302)
);

OAI21xp33_ASAP7_75t_L g2303 ( 
.A1(n_2181),
.A2(n_747),
.B(n_739),
.Y(n_2303)
);

OAI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2257),
.A2(n_2218),
.B(n_2204),
.C(n_2224),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2262),
.Y(n_2305)
);

NOR4xp25_ASAP7_75t_L g2306 ( 
.A(n_2282),
.B(n_2209),
.C(n_2188),
.D(n_2245),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2250),
.A2(n_2201),
.B1(n_2223),
.B2(n_2194),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2250),
.A2(n_2286),
.B1(n_2276),
.B2(n_2258),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2261),
.B(n_2233),
.Y(n_2309)
);

INVx4_ASAP7_75t_L g2310 ( 
.A(n_2277),
.Y(n_2310)
);

OAI211xp5_ASAP7_75t_L g2311 ( 
.A1(n_2263),
.A2(n_2231),
.B(n_125),
.C(n_123),
.Y(n_2311)
);

NAND3xp33_ASAP7_75t_L g2312 ( 
.A(n_2291),
.B(n_615),
.C(n_570),
.Y(n_2312)
);

OR3x2_ASAP7_75t_L g2313 ( 
.A(n_2254),
.B(n_124),
.C(n_126),
.Y(n_2313)
);

NAND5xp2_ASAP7_75t_L g2314 ( 
.A(n_2266),
.B(n_127),
.C(n_1353),
.D(n_1387),
.E(n_603),
.Y(n_2314)
);

AOI211xp5_ASAP7_75t_L g2315 ( 
.A1(n_2294),
.A2(n_729),
.B(n_570),
.C(n_615),
.Y(n_2315)
);

OA22x2_ASAP7_75t_L g2316 ( 
.A1(n_2284),
.A2(n_1325),
.B1(n_1305),
.B2(n_1334),
.Y(n_2316)
);

NOR2xp67_ASAP7_75t_L g2317 ( 
.A(n_2274),
.B(n_130),
.Y(n_2317)
);

OAI211xp5_ASAP7_75t_L g2318 ( 
.A1(n_2268),
.A2(n_729),
.B(n_657),
.C(n_634),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2265),
.B(n_516),
.Y(n_2319)
);

AOI21xp33_ASAP7_75t_SL g2320 ( 
.A1(n_2280),
.A2(n_131),
.B(n_135),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2264),
.Y(n_2321)
);

XNOR2x1_ASAP7_75t_L g2322 ( 
.A(n_2260),
.B(n_137),
.Y(n_2322)
);

NOR4xp25_ASAP7_75t_L g2323 ( 
.A(n_2290),
.B(n_1319),
.C(n_1332),
.D(n_1300),
.Y(n_2323)
);

AND3x2_ASAP7_75t_L g2324 ( 
.A(n_2251),
.B(n_1327),
.C(n_1324),
.Y(n_2324)
);

NOR2x1p5_ASAP7_75t_L g2325 ( 
.A(n_2278),
.B(n_615),
.Y(n_2325)
);

XNOR2x1_ASAP7_75t_L g2326 ( 
.A(n_2272),
.B(n_138),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2285),
.Y(n_2327)
);

OAI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2271),
.A2(n_634),
.B(n_729),
.C(n_657),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_2255),
.B(n_615),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2279),
.B(n_516),
.Y(n_2330)
);

NAND4xp25_ASAP7_75t_SL g2331 ( 
.A(n_2301),
.B(n_2281),
.C(n_2287),
.D(n_2302),
.Y(n_2331)
);

NAND4xp25_ASAP7_75t_SL g2332 ( 
.A(n_2298),
.B(n_1387),
.C(n_1528),
.D(n_1525),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2269),
.A2(n_1299),
.B1(n_1311),
.B2(n_1307),
.Y(n_2333)
);

AOI22xp33_ASAP7_75t_L g2334 ( 
.A1(n_2293),
.A2(n_516),
.B1(n_557),
.B2(n_603),
.Y(n_2334)
);

NOR4xp25_ASAP7_75t_L g2335 ( 
.A(n_2303),
.B(n_1048),
.C(n_1258),
.D(n_1252),
.Y(n_2335)
);

NAND4xp25_ASAP7_75t_L g2336 ( 
.A(n_2288),
.B(n_1527),
.C(n_1523),
.D(n_1501),
.Y(n_2336)
);

NOR4xp25_ASAP7_75t_L g2337 ( 
.A(n_2273),
.B(n_2297),
.C(n_2253),
.D(n_2259),
.Y(n_2337)
);

OAI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2292),
.A2(n_2299),
.B(n_2295),
.Y(n_2338)
);

INVxp67_ASAP7_75t_SL g2339 ( 
.A(n_2252),
.Y(n_2339)
);

AO22x2_ASAP7_75t_L g2340 ( 
.A1(n_2300),
.A2(n_2267),
.B1(n_2289),
.B2(n_2256),
.Y(n_2340)
);

AOI211x1_ASAP7_75t_L g2341 ( 
.A1(n_2270),
.A2(n_603),
.B(n_557),
.C(n_516),
.Y(n_2341)
);

INVxp67_ASAP7_75t_SL g2342 ( 
.A(n_2300),
.Y(n_2342)
);

INVx1_ASAP7_75t_SL g2343 ( 
.A(n_2296),
.Y(n_2343)
);

AO22x2_ASAP7_75t_L g2344 ( 
.A1(n_2275),
.A2(n_1527),
.B1(n_1519),
.B2(n_1522),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2283),
.Y(n_2345)
);

NOR2x2_ASAP7_75t_L g2346 ( 
.A(n_2272),
.B(n_1532),
.Y(n_2346)
);

BUFx3_ASAP7_75t_L g2347 ( 
.A(n_2250),
.Y(n_2347)
);

OAI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2257),
.A2(n_1620),
.B1(n_1588),
.B2(n_1551),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2257),
.B(n_516),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_SL g2350 ( 
.A(n_2257),
.B(n_1239),
.C(n_1236),
.Y(n_2350)
);

NOR3xp33_ASAP7_75t_L g2351 ( 
.A(n_2347),
.B(n_603),
.C(n_557),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2308),
.A2(n_557),
.B1(n_603),
.B2(n_1311),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2327),
.B(n_557),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2325),
.Y(n_2354)
);

BUFx2_ASAP7_75t_L g2355 ( 
.A(n_2305),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2342),
.B(n_2340),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2313),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2346),
.Y(n_2358)
);

NAND4xp25_ASAP7_75t_L g2359 ( 
.A(n_2317),
.B(n_603),
.C(n_1411),
.D(n_1413),
.Y(n_2359)
);

AND4x1_ASAP7_75t_L g2360 ( 
.A(n_2306),
.B(n_603),
.C(n_143),
.D(n_144),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2310),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2340),
.Y(n_2362)
);

XNOR2x1_ASAP7_75t_L g2363 ( 
.A(n_2343),
.B(n_139),
.Y(n_2363)
);

BUFx2_ASAP7_75t_L g2364 ( 
.A(n_2326),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2321),
.B(n_634),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2338),
.B(n_634),
.Y(n_2366)
);

BUFx2_ASAP7_75t_L g2367 ( 
.A(n_2344),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2316),
.B(n_657),
.Y(n_2368)
);

AOI221xp5_ASAP7_75t_L g2369 ( 
.A1(n_2331),
.A2(n_657),
.B1(n_729),
.B2(n_1296),
.C(n_1307),
.Y(n_2369)
);

HB1xp67_ASAP7_75t_L g2370 ( 
.A(n_2322),
.Y(n_2370)
);

INVx2_ASAP7_75t_SL g2371 ( 
.A(n_2344),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2329),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2309),
.B(n_145),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2341),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2330),
.B(n_150),
.Y(n_2375)
);

OAI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2307),
.A2(n_1296),
.B1(n_1311),
.B2(n_1307),
.C(n_1299),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2345),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2324),
.Y(n_2378)
);

AND2x2_ASAP7_75t_SL g2379 ( 
.A(n_2337),
.B(n_1299),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2349),
.B(n_152),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2319),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2339),
.B(n_2333),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2334),
.B(n_153),
.Y(n_2383)
);

AO22x2_ASAP7_75t_L g2384 ( 
.A1(n_2311),
.A2(n_1413),
.B1(n_1481),
.B2(n_1501),
.Y(n_2384)
);

OAI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2304),
.A2(n_1124),
.B(n_1123),
.Y(n_2385)
);

NAND4xp25_ASAP7_75t_L g2386 ( 
.A(n_2314),
.B(n_1481),
.C(n_1509),
.D(n_1504),
.Y(n_2386)
);

AOI221xp5_ASAP7_75t_L g2387 ( 
.A1(n_2323),
.A2(n_2335),
.B1(n_2348),
.B2(n_2320),
.C(n_2336),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2332),
.Y(n_2388)
);

NAND5xp2_ASAP7_75t_SL g2389 ( 
.A(n_2328),
.B(n_2318),
.C(n_2315),
.D(n_2312),
.E(n_2350),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2347),
.Y(n_2390)
);

XNOR2xp5_ASAP7_75t_L g2391 ( 
.A(n_2308),
.B(n_155),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2308),
.A2(n_1124),
.B(n_1123),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2347),
.B(n_156),
.Y(n_2393)
);

NAND4xp75_ASAP7_75t_L g2394 ( 
.A(n_2308),
.B(n_1262),
.C(n_1502),
.D(n_1500),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2308),
.A2(n_1141),
.B1(n_1620),
.B2(n_1632),
.Y(n_2395)
);

NAND3xp33_ASAP7_75t_L g2396 ( 
.A(n_2308),
.B(n_1124),
.C(n_1123),
.Y(n_2396)
);

NAND5xp2_ASAP7_75t_L g2397 ( 
.A(n_2356),
.B(n_159),
.C(n_160),
.D(n_167),
.E(n_172),
.Y(n_2397)
);

OAI211xp5_ASAP7_75t_SL g2398 ( 
.A1(n_2362),
.A2(n_176),
.B(n_179),
.C(n_183),
.Y(n_2398)
);

NOR2x2_ASAP7_75t_L g2399 ( 
.A(n_2390),
.B(n_190),
.Y(n_2399)
);

OR4x2_ASAP7_75t_L g2400 ( 
.A(n_2355),
.B(n_197),
.C(n_200),
.D(n_204),
.Y(n_2400)
);

XOR2xp5_ASAP7_75t_L g2401 ( 
.A(n_2370),
.B(n_208),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2361),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2377),
.B(n_209),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2364),
.B(n_211),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2363),
.Y(n_2405)
);

NOR3xp33_ASAP7_75t_L g2406 ( 
.A(n_2354),
.B(n_1287),
.C(n_1141),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2353),
.B(n_216),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2357),
.B(n_1591),
.Y(n_2408)
);

NOR4xp75_ASAP7_75t_L g2409 ( 
.A(n_2375),
.B(n_219),
.C(n_220),
.D(n_223),
.Y(n_2409)
);

INVxp67_ASAP7_75t_L g2410 ( 
.A(n_2367),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2391),
.Y(n_2411)
);

OAI22x1_ASAP7_75t_L g2412 ( 
.A1(n_2360),
.A2(n_2391),
.B1(n_2374),
.B2(n_2371),
.Y(n_2412)
);

OR2x6_ASAP7_75t_L g2413 ( 
.A(n_2358),
.B(n_1049),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2373),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_L g2415 ( 
.A(n_2372),
.B(n_1123),
.C(n_1124),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2380),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2378),
.B(n_225),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2365),
.Y(n_2418)
);

INVx2_ASAP7_75t_SL g2419 ( 
.A(n_2393),
.Y(n_2419)
);

OAI221xp5_ASAP7_75t_L g2420 ( 
.A1(n_2359),
.A2(n_1169),
.B1(n_1497),
.B2(n_1493),
.C(n_1457),
.Y(n_2420)
);

AOI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2382),
.A2(n_1141),
.B1(n_1611),
.B2(n_1606),
.Y(n_2421)
);

AND2x2_ASAP7_75t_SL g2422 ( 
.A(n_2379),
.B(n_2368),
.Y(n_2422)
);

NAND3x1_ASAP7_75t_L g2423 ( 
.A(n_2352),
.B(n_226),
.C(n_233),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2388),
.A2(n_1141),
.B1(n_1611),
.B2(n_1606),
.Y(n_2424)
);

NOR2x1p5_ASAP7_75t_L g2425 ( 
.A(n_2383),
.B(n_1053),
.Y(n_2425)
);

NOR3xp33_ASAP7_75t_SL g2426 ( 
.A(n_2366),
.B(n_234),
.C(n_243),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2381),
.B(n_244),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2402),
.Y(n_2428)
);

INVxp67_ASAP7_75t_L g2429 ( 
.A(n_2419),
.Y(n_2429)
);

AOI22xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2410),
.A2(n_2412),
.B1(n_2414),
.B2(n_2401),
.Y(n_2430)
);

XNOR2xp5_ASAP7_75t_L g2431 ( 
.A(n_2411),
.B(n_2384),
.Y(n_2431)
);

INVx4_ASAP7_75t_L g2432 ( 
.A(n_2422),
.Y(n_2432)
);

XNOR2xp5_ASAP7_75t_L g2433 ( 
.A(n_2416),
.B(n_2405),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2407),
.Y(n_2434)
);

AOI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_2418),
.A2(n_2387),
.B1(n_2386),
.B2(n_2395),
.Y(n_2435)
);

XNOR2xp5_ASAP7_75t_L g2436 ( 
.A(n_2409),
.B(n_2384),
.Y(n_2436)
);

NAND2xp33_ASAP7_75t_SL g2437 ( 
.A(n_2426),
.B(n_2404),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_SL g2438 ( 
.A1(n_2400),
.A2(n_2396),
.B1(n_2376),
.B2(n_2385),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_2408),
.Y(n_2439)
);

INVx4_ASAP7_75t_L g2440 ( 
.A(n_2413),
.Y(n_2440)
);

INVxp67_ASAP7_75t_L g2441 ( 
.A(n_2403),
.Y(n_2441)
);

AO22x2_ASAP7_75t_L g2442 ( 
.A1(n_2417),
.A2(n_2351),
.B1(n_2392),
.B2(n_2394),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_SL g2443 ( 
.A1(n_2413),
.A2(n_2420),
.B1(n_2399),
.B2(n_2415),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2425),
.Y(n_2444)
);

INVx1_ASAP7_75t_SL g2445 ( 
.A(n_2427),
.Y(n_2445)
);

AND3x4_ASAP7_75t_L g2446 ( 
.A(n_2397),
.B(n_2389),
.C(n_2369),
.Y(n_2446)
);

INVx3_ASAP7_75t_SL g2447 ( 
.A(n_2432),
.Y(n_2447)
);

OR2x6_ASAP7_75t_L g2448 ( 
.A(n_2428),
.B(n_2423),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2429),
.Y(n_2449)
);

OAI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2441),
.A2(n_2424),
.B1(n_2421),
.B2(n_2398),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2445),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_2437),
.B(n_2406),
.Y(n_2452)
);

AOI222xp33_ASAP7_75t_L g2453 ( 
.A1(n_2433),
.A2(n_1141),
.B1(n_1359),
.B2(n_1169),
.C1(n_1053),
.C2(n_1389),
.Y(n_2453)
);

XOR2xp5_ASAP7_75t_L g2454 ( 
.A(n_2430),
.B(n_247),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_SL g2455 ( 
.A1(n_2436),
.A2(n_1489),
.B1(n_1450),
.B2(n_1482),
.C(n_1516),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2434),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2439),
.B(n_1872),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2431),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2440),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2444),
.Y(n_2460)
);

CKINVDCx20_ASAP7_75t_R g2461 ( 
.A(n_2447),
.Y(n_2461)
);

AOI22x1_ASAP7_75t_SL g2462 ( 
.A1(n_2459),
.A2(n_2446),
.B1(n_2435),
.B2(n_2443),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2449),
.Y(n_2463)
);

AO22x2_ASAP7_75t_L g2464 ( 
.A1(n_2451),
.A2(n_2438),
.B1(n_2442),
.B2(n_262),
.Y(n_2464)
);

OAI22x1_ASAP7_75t_L g2465 ( 
.A1(n_2456),
.A2(n_1169),
.B1(n_1051),
.B2(n_264),
.Y(n_2465)
);

AND2x4_ASAP7_75t_L g2466 ( 
.A(n_2458),
.B(n_249),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2448),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2448),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2460),
.B(n_257),
.Y(n_2469)
);

AOI21x1_ASAP7_75t_L g2470 ( 
.A1(n_2454),
.A2(n_2452),
.B(n_2450),
.Y(n_2470)
);

OAI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_2461),
.A2(n_2455),
.B1(n_2457),
.B2(n_2453),
.Y(n_2471)
);

AO22x2_ASAP7_75t_L g2472 ( 
.A1(n_2463),
.A2(n_267),
.B1(n_274),
.B2(n_276),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2467),
.Y(n_2473)
);

XNOR2xp5_ASAP7_75t_L g2474 ( 
.A(n_2462),
.B(n_278),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2464),
.Y(n_2475)
);

OAI22x1_ASAP7_75t_L g2476 ( 
.A1(n_2468),
.A2(n_1169),
.B1(n_1051),
.B2(n_288),
.Y(n_2476)
);

OA21x2_ASAP7_75t_L g2477 ( 
.A1(n_2473),
.A2(n_2470),
.B(n_2466),
.Y(n_2477)
);

AOI22xp33_ASAP7_75t_L g2478 ( 
.A1(n_2475),
.A2(n_2464),
.B1(n_2474),
.B2(n_2472),
.Y(n_2478)
);

OAI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2471),
.A2(n_2469),
.B(n_2465),
.Y(n_2479)
);

OAI21xp5_ASAP7_75t_SL g2480 ( 
.A1(n_2476),
.A2(n_1053),
.B(n_1389),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2477),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2478),
.Y(n_2482)
);

XOR2xp5_ASAP7_75t_L g2483 ( 
.A(n_2479),
.B(n_282),
.Y(n_2483)
);

OR2x6_ASAP7_75t_L g2484 ( 
.A(n_2481),
.B(n_2480),
.Y(n_2484)
);

OAI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_2482),
.A2(n_1359),
.B(n_1051),
.Y(n_2485)
);

OR2x6_ASAP7_75t_L g2486 ( 
.A(n_2483),
.B(n_1382),
.Y(n_2486)
);

XNOR2xp5_ASAP7_75t_L g2487 ( 
.A(n_2484),
.B(n_2486),
.Y(n_2487)
);

XNOR2xp5_ASAP7_75t_L g2488 ( 
.A(n_2485),
.B(n_286),
.Y(n_2488)
);

OR2x6_ASAP7_75t_L g2489 ( 
.A(n_2487),
.B(n_1382),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2489),
.A2(n_2488),
.B(n_1051),
.Y(n_2490)
);

AOI211xp5_ASAP7_75t_L g2491 ( 
.A1(n_2490),
.A2(n_1389),
.B(n_1382),
.C(n_295),
.Y(n_2491)
);


endmodule