module fake_aes_3237_n_31 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
AND2x6_ASAP7_75t_L g13 ( .A(n_0), .B(n_7), .Y(n_13) );
CKINVDCx8_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_2), .B(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_1), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_15), .B(n_13), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_20), .B(n_19), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
OAI222xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_14), .B1(n_13), .B2(n_3), .C1(n_1), .C2(n_2), .Y(n_24) );
AOI211xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_21), .B(n_13), .C(n_3), .Y(n_25) );
OAI22xp33_ASAP7_75t_SL g26 ( .A1(n_24), .A2(n_21), .B1(n_5), .B2(n_8), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_28), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_27), .Y(n_30) );
AOI22xp5_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_4), .B1(n_9), .B2(n_11), .Y(n_31) );
endmodule