module fake_jpeg_9486_n_207 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_207);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_18),
.B1(n_17),
.B2(n_19),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_41),
.B1(n_14),
.B2(n_24),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_17),
.B1(n_23),
.B2(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_49),
.B(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_30),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_20),
.B(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_61),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_70),
.B(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_36),
.B1(n_40),
.B2(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_35),
.C(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.C(n_64),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_35),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_35),
.C(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_33),
.B1(n_29),
.B2(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_76),
.B(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_38),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_53),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_70),
.B1(n_64),
.B2(n_53),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_60),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_59),
.C(n_35),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_48),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_63),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_100),
.C(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_63),
.B1(n_58),
.B2(n_43),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_95),
.B1(n_106),
.B2(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_66),
.B1(n_67),
.B2(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_29),
.C(n_39),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_52),
.B1(n_65),
.B2(n_29),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_52),
.B1(n_65),
.B2(n_24),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_78),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_112),
.C(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_85),
.C(n_81),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_76),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_125),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_74),
.B(n_82),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_101),
.B(n_95),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_85),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_135),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_91),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_134),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_39),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_94),
.B1(n_73),
.B2(n_52),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_140),
.B1(n_24),
.B2(n_22),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_110),
.B(n_99),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_73),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_79),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_39),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_79),
.B1(n_65),
.B2(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_124),
.B1(n_118),
.B2(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_125),
.B1(n_112),
.B2(n_123),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_149),
.B1(n_155),
.B2(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_153),
.C(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_83),
.B1(n_51),
.B2(n_39),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_154),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_71),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_22),
.B1(n_24),
.B2(n_2),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_139),
.B(n_141),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_170),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_168),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_134),
.C(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_166),
.C(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_170),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_169),
.B1(n_153),
.B2(n_151),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_176),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_157),
.B1(n_136),
.B2(n_128),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_174),
.B1(n_10),
.B2(n_3),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_4),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_179),
.C(n_158),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_6),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_8),
.B(n_1),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_181),
.B(n_178),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_5),
.C(n_1),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_164),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_190),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_160),
.B(n_2),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_186),
.B(n_9),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_185),
.B(n_189),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_177),
.B(n_10),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_196),
.B1(n_194),
.B2(n_12),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_12),
.C(n_13),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_200),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_0),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_199),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_202),
.Y(n_207)
);


endmodule