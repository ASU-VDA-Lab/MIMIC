module fake_jpeg_21276_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_43),
.B(n_56),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_49),
.B1(n_22),
.B2(n_29),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_21),
.B(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_59),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2xp67_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_21),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_23),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_75),
.C(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_77),
.B1(n_88),
.B2(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_25),
.B1(n_18),
.B2(n_29),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_37),
.C(n_23),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_26),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_54),
.B1(n_53),
.B2(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_53),
.B1(n_26),
.B2(n_17),
.Y(n_94)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_22),
.B1(n_19),
.B2(n_28),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_37),
.Y(n_90)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_61),
.B1(n_81),
.B2(n_86),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_99),
.B1(n_106),
.B2(n_112),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_53),
.B1(n_26),
.B2(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_111),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_65),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_72),
.B1(n_78),
.B2(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_124),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_128),
.B1(n_136),
.B2(n_90),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_74),
.B1(n_69),
.B2(n_61),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_66),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_69),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_98),
.C(n_103),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_83),
.B1(n_81),
.B2(n_76),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_91),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_5),
.B(n_6),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_97),
.B(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_89),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_64),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_162),
.C(n_167),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_106),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_126),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_100),
.B1(n_102),
.B2(n_108),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_119),
.B1(n_134),
.B2(n_131),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_112),
.B1(n_90),
.B2(n_99),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_138),
.B1(n_116),
.B2(n_124),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_97),
.C(n_109),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_113),
.B(n_101),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_127),
.B(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_80),
.C(n_83),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_79),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_122),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_165),
.B1(n_166),
.B2(n_147),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_179),
.B1(n_154),
.B2(n_162),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_175),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_127),
.C(n_117),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_181),
.C(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_160),
.A3(n_151),
.B1(n_150),
.B2(n_168),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_183),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_134),
.C(n_133),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_76),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_184),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_145),
.C(n_165),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_133),
.C(n_8),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_146),
.C(n_158),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_7),
.B(n_8),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_163),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_195),
.B1(n_182),
.B2(n_174),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_159),
.B1(n_178),
.B2(n_164),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_203),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_151),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_10),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_161),
.CI(n_152),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_157),
.C(n_144),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_156),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_144),
.C(n_163),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_147),
.B1(n_156),
.B2(n_9),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_171),
.B1(n_169),
.B2(n_173),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_218),
.B1(n_199),
.B2(n_198),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_172),
.B(n_176),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_201),
.B(n_191),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_206),
.A2(n_176),
.B(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_211),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_180),
.B(n_182),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_215),
.Y(n_222)
);

NOR4xp25_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_186),
.C(n_187),
.D(n_147),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_216),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_203),
.C(n_190),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_226),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_190),
.C(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_218),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_200),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_205),
.C(n_11),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_10),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_11),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_224),
.C(n_209),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_210),
.B1(n_207),
.B2(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_236),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_16),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_223),
.C(n_229),
.Y(n_239)
);

AOI21x1_ASAP7_75t_SL g245 ( 
.A1(n_239),
.A2(n_232),
.B(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_226),
.C(n_13),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_244),
.C(n_13),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_12),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_242),
.C(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_14),
.C(n_15),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_14),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_239),
.C(n_15),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_250),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);


endmodule