module fake_aes_11237_n_30 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_0), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
AO22x1_ASAP7_75t_L g11 ( .A1(n_0), .A2(n_5), .B1(n_6), .B2(n_4), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_3), .B(n_2), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_6), .B(n_5), .Y(n_14) );
AO31x2_ASAP7_75t_L g15 ( .A1(n_8), .A2(n_1), .A3(n_3), .B(n_9), .Y(n_15) );
BUFx8_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_12), .B(n_1), .Y(n_17) );
BUFx2_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_10), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_15), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_22), .B(n_16), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_22), .B(n_16), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_16), .Y(n_25) );
AOI222xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_11), .B1(n_21), .B2(n_20), .C1(n_17), .C2(n_22), .Y(n_26) );
NAND4xp25_ASAP7_75t_L g27 ( .A(n_26), .B(n_14), .C(n_18), .D(n_20), .Y(n_27) );
OAI211xp5_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_15), .B(n_21), .C(n_26), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_27), .B(n_15), .Y(n_29) );
AOI21xp33_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_28), .B(n_11), .Y(n_30) );
endmodule