module real_jpeg_14295_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_275, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_275;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_9),
.B(n_30),
.C(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_0),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_0),
.B(n_35),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_0),
.B(n_52),
.C(n_55),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_42),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_27),
.C(n_31),
.Y(n_174)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_6),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_6),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_8),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_207)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_11),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_11),
.A2(n_24),
.B1(n_43),
.B2(n_44),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_11),
.A2(n_24),
.B1(n_54),
.B2(n_55),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_83),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_81),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_68),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_68),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_60),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_36),
.C(n_47),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_17),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_17),
.A2(n_70),
.B1(n_114),
.B2(n_124),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_17),
.B(n_124),
.C(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_17),
.A2(n_70),
.B1(n_92),
.B2(n_93),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_19),
.A2(n_29),
.B(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_21),
.B(n_174),
.Y(n_173)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_25),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_25),
.B(n_35),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_29),
.A2(n_62),
.B(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_40),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_33),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_34),
.A2(n_40),
.B(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_34),
.B(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_34),
.B(n_58),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_36),
.A2(n_47),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_36)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_44),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_75),
.C(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_47),
.A2(n_74),
.B1(n_77),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_58),
.B(n_59),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_48),
.A2(n_58),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_99),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_49),
.A2(n_53),
.B1(n_97),
.B2(n_99),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_49),
.A2(n_53),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_54),
.B(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_96),
.B(n_98),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_58),
.A2(n_98),
.B(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_59),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_67),
.B1(n_94),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_66),
.A2(n_67),
.B(n_115),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_79),
.B(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.C(n_76),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_69),
.A2(n_75),
.B1(n_176),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_69),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_70),
.B(n_93),
.C(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_75),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_75),
.A2(n_176),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_75),
.A2(n_176),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_76),
.B(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_77),
.Y(n_261)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_253),
.B(n_270),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_231),
.B(n_252),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_214),
.B(n_230),
.Y(n_86)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_183),
.A3(n_209),
.B1(n_212),
.B2(n_213),
.C(n_275),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_166),
.B(n_182),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_132),
.B(n_165),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_111),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_91),
.B(n_111),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.C(n_100),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_92),
.A2(n_93),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_93),
.B(n_176),
.C(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_95),
.A2(n_136),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_95),
.A2(n_149),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_100),
.A2(n_101),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_106),
.B(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_109),
.A2(n_110),
.B1(n_190),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_110),
.A2(n_122),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_126),
.B2(n_127),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_129),
.C(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_124),
.B2(n_125),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_117),
.C(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_124),
.A2(n_247),
.B(n_250),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_124),
.B(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_131),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_141),
.C(n_143),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_131),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_129),
.B(n_206),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_159),
.B(n_164),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_145),
.B(n_158),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_143),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_157),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_189),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_154),
.B(n_156),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_160),
.B(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_168),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_171),
.C(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_197),
.C(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_193),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_193),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_192),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_188),
.CI(n_192),
.CON(n_211),
.SN(n_211)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_208),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_203),
.B2(n_204),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_204),
.C(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_211),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_229),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_229),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_218),
.C(n_223),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_228),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_237),
.B(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_251),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_245),
.B2(n_246),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_245),
.C(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_250),
.A2(n_257),
.B1(n_258),
.B2(n_262),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_250),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_265),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_269),
.Y(n_272)
);


endmodule