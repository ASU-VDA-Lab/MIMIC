module fake_jpeg_13643_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_155;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_14),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_42),
.B(n_55),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_62),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_1),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_22),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_73),
.Y(n_99)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_15),
.B(n_5),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_79),
.Y(n_101)
);

NAND2x1_ASAP7_75t_SL g75 ( 
.A(n_33),
.B(n_5),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_26),
.C(n_40),
.Y(n_97)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_77),
.Y(n_114)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_6),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_52),
.B1(n_61),
.B2(n_65),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_81),
.A2(n_85),
.B1(n_95),
.B2(n_100),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_28),
.B1(n_40),
.B2(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_44),
.A2(n_33),
.B1(n_39),
.B2(n_34),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_12),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_41),
.B1(n_39),
.B2(n_34),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_45),
.A2(n_19),
.B1(n_18),
.B2(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_125),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_20),
.B1(n_19),
.B2(n_30),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_115),
.B1(n_80),
.B2(n_38),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_30),
.B1(n_32),
.B2(n_31),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_17),
.B1(n_31),
.B2(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_28),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_26),
.B1(n_17),
.B2(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_123),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_7),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_78),
.C(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_62),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_50),
.A2(n_38),
.B1(n_11),
.B2(n_12),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_7),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_11),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_120),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_135),
.B(n_155),
.C(n_159),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_164),
.B1(n_147),
.B2(n_168),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_14),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_14),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_38),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_99),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_87),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_107),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_160),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_98),
.B(n_117),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_163),
.C(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_119),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_128),
.B1(n_95),
.B2(n_82),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_134),
.B1(n_136),
.B2(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_108),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_165),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_96),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_103),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_125),
.B(n_111),
.C(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_199),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_90),
.B1(n_111),
.B2(n_112),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_178),
.B1(n_132),
.B2(n_143),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_130),
.B1(n_161),
.B2(n_145),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_158),
.C(n_150),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_193),
.C(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_158),
.C(n_152),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_129),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_205),
.B(n_214),
.Y(n_239)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_193),
.C(n_181),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_157),
.B1(n_169),
.B2(n_165),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_175),
.B1(n_188),
.B2(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_166),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_154),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_217),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_156),
.B(n_170),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_227),
.B(n_200),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_174),
.B1(n_196),
.B2(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_225),
.B1(n_195),
.B2(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_172),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_242),
.C(n_247),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_209),
.B1(n_222),
.B2(n_225),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_204),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_175),
.B(n_194),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_221),
.B(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_201),
.C(n_191),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_202),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_218),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_183),
.C(n_202),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

OAI322xp33_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_258),
.A3(n_239),
.B1(n_240),
.B2(n_236),
.C1(n_214),
.C2(n_234),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_259),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_245),
.B(n_203),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_241),
.B(n_237),
.C(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_217),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_263),
.B(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_260),
.B(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_243),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_269),
.B1(n_239),
.B2(n_255),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_234),
.B(n_247),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_273),
.B(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_229),
.B1(n_207),
.B2(n_228),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_242),
.B(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_213),
.C(n_212),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_257),
.C(n_261),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_280),
.Y(n_285)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_254),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_264),
.B(n_283),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_283),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_263),
.B(n_249),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_251),
.B1(n_264),
.B2(n_210),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_211),
.C(n_226),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_268),
.B1(n_251),
.B2(n_264),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_289),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_272),
.B(n_281),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_286),
.Y(n_296)
);

OAI31xp33_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_272),
.A3(n_223),
.B(n_246),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.C(n_288),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_206),
.C(n_246),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_246),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_287),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_295),
.B(n_297),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_285),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_300),
.B1(n_286),
.B2(n_294),
.Y(n_302)
);

XNOR2x2_ASAP7_75t_SL g303 ( 
.A(n_302),
.B(n_197),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_303),
.B(n_184),
.Y(n_304)
);


endmodule