module fake_jpeg_1773_n_105 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_39),
.B(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_39),
.B1(n_34),
.B2(n_32),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_34),
.B1(n_32),
.B2(n_38),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_61),
.B1(n_52),
.B2(n_2),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_50),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_29),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_72),
.B(n_3),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_22),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_60),
.C(n_15),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_84),
.C(n_67),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_52),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_85),
.B1(n_74),
.B2(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_84),
.B1(n_83),
.B2(n_86),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_17),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_77),
.C(n_69),
.Y(n_97)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_24),
.A3(n_28),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.C(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_97),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_96),
.B1(n_95),
.B2(n_90),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_94),
.B1(n_88),
.B2(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_25),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_26),
.C(n_27),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_8),
.C(n_9),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_9),
.Y(n_105)
);


endmodule