module fake_jpeg_6958_n_251 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_22),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_20),
.Y(n_42)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_37),
.B1(n_23),
.B2(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_15),
.B1(n_19),
.B2(n_18),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_14),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_51),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_18),
.B1(n_15),
.B2(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_14),
.B1(n_27),
.B2(n_21),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_30),
.A2(n_24),
.B(n_17),
.C(n_25),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_61),
.B1(n_74),
.B2(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_35),
.B1(n_33),
.B2(n_38),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_35),
.B1(n_36),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_59),
.B1(n_47),
.B2(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_79),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_68),
.Y(n_89)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_70),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_35),
.A3(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_49),
.B(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_35),
.B1(n_33),
.B2(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_32),
.B1(n_31),
.B2(n_36),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_43),
.B1(n_49),
.B2(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_29),
.B1(n_16),
.B2(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_43),
.B1(n_52),
.B2(n_51),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_90),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_54),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_104),
.B1(n_68),
.B2(n_74),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_57),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_60),
.Y(n_119)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_95),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_32),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_106),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_76),
.B1(n_66),
.B2(n_78),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_101),
.B1(n_86),
.B2(n_87),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_118),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_73),
.C(n_78),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_116),
.C(n_31),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_78),
.C(n_76),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_121),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_0),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_90),
.B(n_31),
.Y(n_140)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_123),
.A2(n_96),
.B(n_82),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_134),
.CI(n_148),
.CON(n_164),
.SN(n_164)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_101),
.B1(n_87),
.B2(n_85),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_103),
.B(n_84),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_92),
.B(n_41),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_140),
.Y(n_158)
);

OAI22x1_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_41),
.B1(n_92),
.B2(n_70),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_102),
.B1(n_64),
.B2(n_109),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_65),
.B1(n_90),
.B2(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_113),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_102),
.B1(n_100),
.B2(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_107),
.C(n_117),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_116),
.B(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_154),
.B(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_161),
.C(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_119),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_133),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_108),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_108),
.B(n_126),
.C(n_113),
.D(n_115),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_158),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_131),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_137),
.B1(n_132),
.B2(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_176),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_135),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_159),
.B1(n_153),
.B2(n_149),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_137),
.B1(n_144),
.B2(n_130),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_24),
.B1(n_2),
.B2(n_1),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_138),
.B1(n_147),
.B2(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_143),
.B(n_147),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_164),
.B1(n_24),
.B2(n_17),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_127),
.C(n_64),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.C(n_152),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_127),
.C(n_25),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_194),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_195),
.C(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_196),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_159),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_157),
.C(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_164),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_187),
.C(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_175),
.C(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_205),
.B(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_183),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_191),
.B(n_189),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_184),
.C(n_174),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_185),
.C(n_172),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_180),
.C(n_176),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_197),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_204),
.B(n_203),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_213),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_6),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_223),
.B(n_224),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_1),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_1),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_229),
.B(n_231),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_212),
.B(n_4),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_221),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_3),
.B(n_5),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_6),
.B(n_7),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_235),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_13),
.C(n_10),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_239),
.B(n_8),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_237),
.A3(n_236),
.B1(n_12),
.B2(n_13),
.C1(n_11),
.C2(n_9),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_12),
.C(n_9),
.Y(n_247)
);

OAI311xp33_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_9),
.A3(n_11),
.B1(n_244),
.C1(n_246),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_243),
.B(n_242),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_11),
.Y(n_251)
);


endmodule