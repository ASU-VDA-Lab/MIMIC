module real_aes_1127_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_691;
wire n_498;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_0), .B(n_120), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_1), .A2(n_129), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_2), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_3), .B(n_136), .Y(n_199) );
INVx1_ASAP7_75t_L g127 ( .A(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_5), .B(n_136), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_6), .B(n_140), .Y(n_492) );
INVx1_ASAP7_75t_L g526 ( .A(n_7), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_8), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_8), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_9), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_10), .Y(n_564) );
NAND2xp33_ASAP7_75t_L g137 ( .A(n_11), .B(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
AOI221x1_ASAP7_75t_L g215 ( .A1(n_13), .A2(n_25), .B1(n_120), .B2(n_129), .C(n_216), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_14), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_15), .B(n_120), .Y(n_119) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_16), .A2(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g501 ( .A(n_17), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_18), .B(n_154), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_19), .B(n_136), .Y(n_163) );
AO21x1_ASAP7_75t_L g194 ( .A1(n_20), .A2(n_120), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g445 ( .A(n_21), .Y(n_445) );
INVx1_ASAP7_75t_L g499 ( .A(n_22), .Y(n_499) );
INVx1_ASAP7_75t_SL g509 ( .A(n_23), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_24), .B(n_121), .Y(n_592) );
NAND2x1_ASAP7_75t_L g185 ( .A(n_26), .B(n_136), .Y(n_185) );
AOI33xp33_ASAP7_75t_L g538 ( .A1(n_27), .A2(n_54), .A3(n_476), .B1(n_481), .B2(n_539), .B3(n_540), .Y(n_538) );
NAND2x1_ASAP7_75t_L g173 ( .A(n_28), .B(n_138), .Y(n_173) );
INVx1_ASAP7_75t_L g558 ( .A(n_29), .Y(n_558) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_30), .A2(n_88), .B(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g141 ( .A(n_30), .B(n_88), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_31), .B(n_484), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_32), .B(n_138), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_33), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_34), .B(n_138), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_35), .A2(n_129), .B(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g126 ( .A(n_36), .B(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g130 ( .A(n_36), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g475 ( .A(n_36), .Y(n_475) );
OR2x6_ASAP7_75t_L g443 ( .A(n_37), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_38), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_39), .B(n_120), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_40), .B(n_484), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_41), .A2(n_140), .B1(n_147), .B2(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_42), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_43), .B(n_121), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_44), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_45), .B(n_138), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_46), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_46), .Y(n_798) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_47), .A2(n_104), .B1(n_450), .B2(n_455), .C1(n_811), .C2(n_816), .Y(n_103) );
XNOR2xp5_ASAP7_75t_SL g105 ( .A(n_47), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_47), .B(n_115), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_48), .B(n_121), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_49), .A2(n_129), .B(n_172), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_50), .Y(n_589) );
XOR2xp5_ASAP7_75t_L g800 ( .A(n_51), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_52), .B(n_138), .Y(n_186) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_53), .A2(n_797), .B1(n_805), .B2(n_807), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_55), .B(n_121), .Y(n_550) );
INVx1_ASAP7_75t_L g123 ( .A(n_56), .Y(n_123) );
INVx1_ASAP7_75t_L g133 ( .A(n_56), .Y(n_133) );
AND2x2_ASAP7_75t_L g551 ( .A(n_57), .B(n_154), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_58), .A2(n_75), .B1(n_473), .B2(n_484), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_59), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_60), .B(n_136), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_61), .B(n_147), .Y(n_566) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_62), .A2(n_473), .B(n_478), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_63), .A2(n_129), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g495 ( .A(n_64), .Y(n_495) );
AO21x1_ASAP7_75t_L g196 ( .A1(n_65), .A2(n_129), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_66), .B(n_120), .Y(n_149) );
INVx1_ASAP7_75t_L g549 ( .A(n_67), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_68), .B(n_120), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_69), .A2(n_473), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g209 ( .A(n_70), .B(n_155), .Y(n_209) );
INVx1_ASAP7_75t_L g125 ( .A(n_71), .Y(n_125) );
INVx1_ASAP7_75t_L g131 ( .A(n_71), .Y(n_131) );
AND2x2_ASAP7_75t_L g177 ( .A(n_72), .B(n_146), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_73), .B(n_484), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_74), .B(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g432 ( .A1(n_76), .A2(n_86), .B1(n_433), .B2(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_76), .Y(n_433) );
AND2x2_ASAP7_75t_L g511 ( .A(n_77), .B(n_146), .Y(n_511) );
INVx1_ASAP7_75t_L g496 ( .A(n_78), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_79), .A2(n_473), .B(n_508), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_80), .A2(n_473), .B(n_533), .C(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g446 ( .A(n_81), .Y(n_446) );
AND2x2_ASAP7_75t_L g145 ( .A(n_82), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_83), .B(n_120), .Y(n_165) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_84), .B(n_146), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_85), .A2(n_473), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g434 ( .A(n_86), .Y(n_434) );
AND2x2_ASAP7_75t_L g195 ( .A(n_87), .B(n_140), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_89), .B(n_138), .Y(n_164) );
AND2x2_ASAP7_75t_L g189 ( .A(n_90), .B(n_146), .Y(n_189) );
INVx1_ASAP7_75t_L g479 ( .A(n_91), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_92), .B(n_136), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_93), .A2(n_129), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_94), .B(n_138), .Y(n_217) );
AND2x2_ASAP7_75t_L g542 ( .A(n_95), .B(n_146), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_96), .A2(n_97), .B1(n_802), .B2(n_803), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_96), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_97), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_98), .B(n_136), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_99), .A2(n_556), .B(n_557), .C(n_559), .Y(n_555) );
BUFx2_ASAP7_75t_L g454 ( .A(n_100), .Y(n_454) );
BUFx2_ASAP7_75t_SL g820 ( .A(n_100), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_101), .A2(n_129), .B(n_134), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_102), .B(n_121), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_437), .B(n_447), .Y(n_104) );
OAI22x1_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_108), .B1(n_430), .B2(n_431), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_108), .A2(n_458), .B1(n_462), .B2(n_796), .Y(n_457) );
INVx2_ASAP7_75t_L g806 ( .A(n_108), .Y(n_806) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_351), .Y(n_108) );
NOR3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_263), .C(n_303), .Y(n_109) );
OAI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_178), .B1(n_227), .B2(n_242), .C(n_245), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_142), .Y(n_112) );
INVx2_ASAP7_75t_L g260 ( .A(n_113), .Y(n_260) );
AND2x2_ASAP7_75t_L g290 ( .A(n_113), .B(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g228 ( .A(n_114), .B(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g235 ( .A(n_114), .B(n_168), .Y(n_235) );
INVx2_ASAP7_75t_L g241 ( .A(n_114), .Y(n_241) );
AND2x2_ASAP7_75t_L g250 ( .A(n_114), .B(n_144), .Y(n_250) );
INVx1_ASAP7_75t_L g266 ( .A(n_114), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_114), .B(n_312), .Y(n_311) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_115), .A2(n_524), .B(n_528), .Y(n_523) );
INVx2_ASAP7_75t_SL g533 ( .A(n_115), .Y(n_533) );
BUFx4f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx3_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
AND2x4_ASAP7_75t_L g140 ( .A(n_117), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_117), .B(n_141), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_128), .B(n_140), .Y(n_118) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_126), .Y(n_120) );
INVx1_ASAP7_75t_L g497 ( .A(n_121), .Y(n_497) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
AND2x6_ASAP7_75t_L g138 ( .A(n_122), .B(n_131), .Y(n_138) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g136 ( .A(n_124), .B(n_133), .Y(n_136) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx5_ASAP7_75t_L g139 ( .A(n_126), .Y(n_139) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_126), .Y(n_559) );
AND2x2_ASAP7_75t_L g132 ( .A(n_127), .B(n_133), .Y(n_132) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_127), .Y(n_486) );
AND2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
BUFx3_ASAP7_75t_L g487 ( .A(n_130), .Y(n_487) );
INVx2_ASAP7_75t_L g477 ( .A(n_131), .Y(n_477) );
AND2x4_ASAP7_75t_L g473 ( .A(n_132), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g481 ( .A(n_133), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B(n_139), .Y(n_134) );
INVxp67_ASAP7_75t_L g502 ( .A(n_136), .Y(n_502) );
INVxp67_ASAP7_75t_L g500 ( .A(n_138), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_139), .A2(n_152), .B(n_153), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_139), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_139), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_139), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_139), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_139), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_139), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_139), .A2(n_479), .B(n_480), .C(n_482), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_139), .B(n_140), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_139), .A2(n_480), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_139), .A2(n_480), .B(n_526), .C(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g536 ( .A(n_139), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_139), .A2(n_480), .B(n_549), .C(n_550), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_139), .A2(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_SL g159 ( .A(n_140), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_140), .B(n_201), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_140), .A2(n_472), .B(n_483), .Y(n_471) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_156), .Y(n_142) );
INVx4_ASAP7_75t_L g231 ( .A(n_143), .Y(n_231) );
AND2x2_ASAP7_75t_L g262 ( .A(n_143), .B(n_169), .Y(n_262) );
AND2x2_ASAP7_75t_L g338 ( .A(n_143), .B(n_312), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_143), .B(n_168), .Y(n_380) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_144), .B(n_168), .Y(n_267) );
AND2x2_ASAP7_75t_L g291 ( .A(n_144), .B(n_169), .Y(n_291) );
BUFx2_ASAP7_75t_L g307 ( .A(n_144), .Y(n_307) );
NOR2x1_ASAP7_75t_SL g410 ( .A(n_144), .B(n_312), .Y(n_410) );
OR2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_148), .Y(n_144) );
INVx3_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_146), .A2(n_188), .B1(n_555), .B2(n_560), .Y(n_554) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_147), .B(n_563), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_154), .Y(n_176) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_154), .A2(n_215), .B(n_219), .Y(n_214) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_154), .A2(n_215), .B(n_219), .Y(n_277) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g287 ( .A(n_156), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_156), .A2(n_354), .B1(n_356), .B2(n_358), .C(n_363), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_156), .B(n_266), .Y(n_373) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_168), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
INVx1_ASAP7_75t_L g282 ( .A(n_158), .Y(n_282) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_166), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_159), .B(n_167), .Y(n_166) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_159), .A2(n_160), .B(n_166), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_165), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_168), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g251 ( .A(n_168), .B(n_239), .Y(n_251) );
INVx2_ASAP7_75t_L g293 ( .A(n_168), .Y(n_293) );
AND2x2_ASAP7_75t_L g426 ( .A(n_168), .B(n_241), .Y(n_426) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_169), .Y(n_283) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_176), .B(n_177), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_176), .A2(n_505), .B(n_511), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_210), .C(n_225), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_190), .Y(n_179) );
INVx2_ASAP7_75t_L g340 ( .A(n_180), .Y(n_340) );
AND2x2_ASAP7_75t_L g385 ( .A(n_180), .B(n_262), .Y(n_385) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g330 ( .A(n_181), .Y(n_330) );
AND2x4_ASAP7_75t_SL g345 ( .A(n_181), .B(n_257), .Y(n_345) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_188), .B(n_189), .Y(n_181) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_182), .A2(n_188), .B(n_189), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_188), .A2(n_203), .B(n_209), .Y(n_202) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_188), .A2(n_203), .B(n_209), .Y(n_222) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_188), .A2(n_545), .B(n_551), .Y(n_544) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_188), .A2(n_545), .B(n_551), .Y(n_574) );
INVx2_ASAP7_75t_L g299 ( .A(n_190), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_190), .B(n_329), .Y(n_355) );
AND2x4_ASAP7_75t_L g388 ( .A(n_190), .B(n_335), .Y(n_388) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_202), .Y(n_190) );
AND2x2_ASAP7_75t_L g226 ( .A(n_191), .B(n_221), .Y(n_226) );
OR2x2_ASAP7_75t_L g256 ( .A(n_191), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_191), .B(n_277), .Y(n_325) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g270 ( .A(n_192), .Y(n_270) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
OAI21x1_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_196), .B(n_200), .Y(n_193) );
INVx1_ASAP7_75t_L g201 ( .A(n_195), .Y(n_201) );
INVx2_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_204), .B(n_208), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_210), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_220), .Y(n_211) );
AND2x2_ASAP7_75t_L g225 ( .A(n_212), .B(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g298 ( .A(n_212), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g383 ( .A(n_212), .Y(n_383) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x4_ASAP7_75t_L g243 ( .A(n_213), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g362 ( .A(n_213), .B(n_222), .Y(n_362) );
AND2x2_ASAP7_75t_L g366 ( .A(n_213), .B(n_232), .Y(n_366) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g335 ( .A(n_214), .Y(n_335) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_214), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_220), .B(n_243), .Y(n_319) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_221), .B(n_244), .Y(n_429) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g233 ( .A(n_222), .B(n_224), .Y(n_233) );
AND2x2_ASAP7_75t_L g315 ( .A(n_222), .B(n_277), .Y(n_315) );
AND2x2_ASAP7_75t_L g334 ( .A(n_222), .B(n_223), .Y(n_334) );
BUFx2_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_223), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx3_ASAP7_75t_L g232 ( .A(n_224), .Y(n_232) );
INVxp67_ASAP7_75t_L g275 ( .A(n_224), .Y(n_275) );
INVx1_ASAP7_75t_L g248 ( .A(n_226), .Y(n_248) );
AND2x2_ASAP7_75t_L g284 ( .A(n_226), .B(n_255), .Y(n_284) );
NAND2xp33_ASAP7_75t_L g365 ( .A(n_226), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g402 ( .A(n_226), .B(n_403), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_230), .B1(n_233), .B2(n_234), .C(n_236), .Y(n_227) );
AND2x2_ASAP7_75t_L g331 ( .A(n_228), .B(n_231), .Y(n_331) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_228), .B(n_291), .Y(n_350) );
AND2x2_ASAP7_75t_L g368 ( .A(n_228), .B(n_293), .Y(n_368) );
AND2x2_ASAP7_75t_L g423 ( .A(n_228), .B(n_262), .Y(n_423) );
INVx1_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_229), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_230), .Y(n_375) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_231), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_231), .B(n_282), .Y(n_357) );
AND2x2_ASAP7_75t_L g324 ( .A(n_232), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g360 ( .A(n_232), .Y(n_360) );
AND2x2_ASAP7_75t_L g269 ( .A(n_233), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_233), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g411 ( .A(n_233), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_233), .B(n_335), .Y(n_421) );
AND2x4_ASAP7_75t_L g337 ( .A(n_234), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g408 ( .A(n_235), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
OR2x2_ASAP7_75t_L g279 ( .A(n_240), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g286 ( .A(n_241), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g317 ( .A(n_241), .B(n_291), .Y(n_317) );
AND2x2_ASAP7_75t_L g391 ( .A(n_241), .B(n_312), .Y(n_391) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g339 ( .A(n_243), .B(n_340), .Y(n_339) );
OAI32xp33_ASAP7_75t_L g404 ( .A1(n_243), .A2(n_405), .A3(n_407), .B1(n_408), .B2(n_411), .Y(n_404) );
AND2x4_ASAP7_75t_L g276 ( .A(n_244), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g374 ( .A(n_244), .B(n_277), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B1(n_252), .B2(n_258), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g363 ( .A1(n_247), .A2(n_261), .B(n_364), .C(n_365), .Y(n_363) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g347 ( .A(n_248), .B(n_275), .Y(n_347) );
INVx1_ASAP7_75t_SL g418 ( .A(n_249), .Y(n_418) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x4_ASAP7_75t_L g321 ( .A(n_251), .B(n_260), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_251), .A2(n_400), .B1(n_401), .B2(n_402), .C(n_404), .Y(n_399) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_256), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_259), .A2(n_289), .B1(n_342), .B2(n_343), .Y(n_341) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_260), .A2(n_378), .B(n_386), .C(n_399), .Y(n_377) );
INVx2_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g297 ( .A(n_262), .B(n_266), .Y(n_297) );
OAI211xp5_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_268), .B(n_271), .C(n_300), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g414 ( .A(n_266), .B(n_410), .Y(n_414) );
OAI32xp33_ASAP7_75t_L g371 ( .A1(n_267), .A2(n_372), .A3(n_374), .B1(n_375), .B2(n_376), .Y(n_371) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_270), .B(n_362), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_278), .B1(n_284), .B2(n_285), .C(n_288), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g428 ( .A(n_275), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_276), .B(n_340), .Y(n_342) );
A2O1A1O1Ixp25_ASAP7_75t_L g413 ( .A1(n_276), .A2(n_345), .B(n_361), .C(n_407), .D(n_414), .Y(n_413) );
AOI31xp33_ASAP7_75t_L g415 ( .A1(n_276), .A2(n_297), .A3(n_407), .B(n_414), .Y(n_415) );
AND2x2_ASAP7_75t_L g329 ( .A(n_277), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_279), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx2_ASAP7_75t_L g406 ( .A(n_281), .Y(n_406) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g401 ( .A(n_282), .B(n_293), .Y(n_401) );
INVx1_ASAP7_75t_L g316 ( .A(n_284), .Y(n_316) );
AND2x2_ASAP7_75t_L g301 ( .A(n_285), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AOI31xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .A3(n_296), .B(n_298), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_291), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g424 ( .A(n_291), .B(n_370), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g369 ( .A(n_293), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g395 ( .A(n_293), .Y(n_395) );
INVxp67_ASAP7_75t_L g364 ( .A(n_294), .Y(n_364) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g302 ( .A(n_298), .Y(n_302) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND3xp33_ASAP7_75t_SL g303 ( .A(n_304), .B(n_320), .C(n_336), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_313), .B1(n_317), .B2(n_318), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g390 ( .A(n_307), .Y(n_390) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_311), .Y(n_370) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_311), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_311), .B(n_380), .Y(n_397) );
NAND2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_331), .B2(n_332), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_329), .A2(n_334), .B1(n_368), .B2(n_369), .C(n_371), .Y(n_367) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
AND2x2_ASAP7_75t_L g344 ( .A(n_335), .B(n_345), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_SL g392 ( .A1(n_335), .A2(n_393), .B(n_397), .C(n_398), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B(n_341), .C(n_346), .Y(n_336) );
AND2x2_ASAP7_75t_L g387 ( .A(n_340), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g398 ( .A(n_345), .Y(n_398) );
AOI21xp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_348), .B(n_349), .Y(n_346) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_377), .C(n_412), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_367), .Y(n_352) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g376 ( .A(n_361), .Y(n_376) );
INVxp67_ASAP7_75t_L g400 ( .A(n_365), .Y(n_400) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g384 ( .A(n_374), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_384), .B2(n_385), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_392), .Y(n_386) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g425 ( .A(n_410), .B(n_426), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_416), .B2(n_419), .C(n_422), .Y(n_412) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI31xp33_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .A3(n_425), .B(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g436 ( .A(n_432), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g821 ( .A(n_439), .Y(n_821) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x6_ASAP7_75t_SL g461 ( .A(n_441), .B(n_443), .Y(n_461) );
OR2x6_ASAP7_75t_SL g796 ( .A(n_441), .B(n_442), .Y(n_796) );
OR2x2_ASAP7_75t_L g810 ( .A(n_441), .B(n_443), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g812 ( .A(n_449), .B(n_813), .Y(n_812) );
CKINVDCx9p33_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx2_ASAP7_75t_L g815 ( .A(n_452), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_452), .A2(n_818), .B(n_821), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g814 ( .A(n_454), .B(n_815), .Y(n_814) );
OAI21xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_797), .B(n_804), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx4_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_460), .A2(n_463), .B1(n_796), .B2(n_806), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND3x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_683), .C(n_760), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_635), .Y(n_464) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_466), .B(n_575), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_512), .B1(n_519), .B2(n_568), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_488), .Y(n_467) );
NOR2xp67_ASAP7_75t_SL g618 ( .A(n_468), .B(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g633 ( .A(n_468), .B(n_634), .Y(n_633) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_468), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_SL g690 ( .A(n_468), .B(n_691), .Y(n_690) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_469), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_469), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g625 ( .A(n_469), .Y(n_625) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_469), .Y(n_630) );
AND2x2_ASAP7_75t_L g659 ( .A(n_469), .B(n_599), .Y(n_659) );
OR2x2_ASAP7_75t_L g663 ( .A(n_469), .B(n_504), .Y(n_663) );
AND2x4_ASAP7_75t_L g676 ( .A(n_469), .B(n_634), .Y(n_676) );
NOR2x1_ASAP7_75t_SL g678 ( .A(n_469), .B(n_491), .Y(n_678) );
AND2x2_ASAP7_75t_L g706 ( .A(n_469), .B(n_584), .Y(n_706) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVxp67_ASAP7_75t_L g565 ( .A(n_473), .Y(n_565) );
NOR2x1p5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g540 ( .A(n_476), .Y(n_540) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x6_ASAP7_75t_L g480 ( .A(n_477), .B(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_480), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
INVxp67_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVx2_ASAP7_75t_L g594 ( .A(n_480), .Y(n_594) );
AND2x2_ASAP7_75t_L g485 ( .A(n_481), .B(n_486), .Y(n_485) );
INVxp33_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
INVx1_ASAP7_75t_L g567 ( .A(n_484), .Y(n_567) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g587 ( .A(n_485), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_487), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_488), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_489), .A2(n_764), .B1(n_766), .B2(n_769), .Y(n_763) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_504), .Y(n_489) );
INVx1_ASAP7_75t_L g518 ( .A(n_490), .Y(n_518) );
AND2x2_ASAP7_75t_L g621 ( .A(n_490), .B(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g626 ( .A(n_490), .B(n_584), .Y(n_626) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g583 ( .A(n_491), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g599 ( .A(n_491), .Y(n_599) );
AND2x2_ASAP7_75t_L g632 ( .A(n_491), .B(n_504), .Y(n_632) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .B(n_503), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_497), .B(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_498) );
INVx2_ASAP7_75t_L g516 ( .A(n_504), .Y(n_516) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_504), .Y(n_601) );
INVx1_ASAP7_75t_L g620 ( .A(n_504), .Y(n_620) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_504), .Y(n_689) );
INVx1_ASAP7_75t_L g701 ( .A(n_504), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI31xp33_ASAP7_75t_SL g755 ( .A1(n_513), .A2(n_756), .A3(n_757), .B(n_758), .Y(n_755) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g680 ( .A(n_515), .B(n_582), .Y(n_680) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g596 ( .A(n_516), .Y(n_596) );
AND2x4_ASAP7_75t_SL g716 ( .A(n_518), .B(n_620), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_519), .A2(n_637), .B(n_640), .Y(n_636) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
INVx2_ASAP7_75t_L g609 ( .A(n_520), .Y(n_609) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g736 ( .A(n_521), .B(n_644), .Y(n_736) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g646 ( .A(n_522), .B(n_552), .Y(n_646) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_523), .B(n_532), .Y(n_606) );
AND2x4_ASAP7_75t_L g616 ( .A(n_523), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g661 ( .A(n_523), .B(n_553), .Y(n_661) );
INVx2_ASAP7_75t_L g669 ( .A(n_523), .Y(n_669) );
INVx1_ASAP7_75t_L g768 ( .A(n_523), .Y(n_768) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_523), .Y(n_777) );
INVx1_ASAP7_75t_L g714 ( .A(n_529), .Y(n_714) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_530), .B(n_543), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g570 ( .A(n_531), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g709 ( .A(n_531), .B(n_644), .Y(n_709) );
AND2x2_ASAP7_75t_L g726 ( .A(n_531), .B(n_544), .Y(n_726) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_532), .B(n_574), .Y(n_749) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_542), .Y(n_532) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_533), .A2(n_534), .B(n_542), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_535), .B(n_541), .Y(n_534) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g672 ( .A(n_543), .B(n_570), .Y(n_672) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_552), .Y(n_543) );
INVx2_ASAP7_75t_L g578 ( .A(n_544), .Y(n_578) );
NOR2xp67_ASAP7_75t_L g759 ( .A(n_544), .B(n_552), .Y(n_759) );
NOR2x1_ASAP7_75t_L g767 ( .A(n_544), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x2_ASAP7_75t_L g675 ( .A(n_552), .B(n_579), .Y(n_675) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_553), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g604 ( .A(n_553), .Y(n_604) );
AND2x4_ASAP7_75t_L g668 ( .A(n_553), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g698 ( .A(n_553), .Y(n_698) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_561), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_569), .A2(n_582), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g696 ( .A(n_570), .B(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g739 ( .A(n_570), .Y(n_739) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g682 ( .A(n_573), .B(n_606), .Y(n_682) );
INVx3_ASAP7_75t_L g644 ( .A(n_574), .Y(n_644) );
AND2x2_ASAP7_75t_L g776 ( .A(n_574), .B(n_777), .Y(n_776) );
NAND3xp33_ASAP7_75t_SL g575 ( .A(n_576), .B(n_607), .C(n_623), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B1(n_597), .B2(n_602), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_577), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g707 ( .A(n_577), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g718 ( .A(n_577), .B(n_613), .Y(n_718) );
AND2x2_ASAP7_75t_L g788 ( .A(n_577), .B(n_661), .Y(n_788) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g617 ( .A(n_579), .Y(n_617) );
INVx1_ASAP7_75t_L g666 ( .A(n_579), .Y(n_666) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI222xp33_ASAP7_75t_L g733 ( .A1(n_581), .A2(n_734), .B1(n_735), .B2(n_737), .C1(n_738), .C2(n_740), .Y(n_733) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_595), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_582), .B(n_609), .Y(n_608) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_582), .B(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g700 ( .A(n_583), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g756 ( .A(n_583), .B(n_630), .Y(n_756) );
INVx2_ASAP7_75t_L g622 ( .A(n_584), .Y(n_622) );
INVx1_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_584), .Y(n_691) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .C(n_589), .Y(n_586) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_596), .Y(n_639) );
INVx3_ASAP7_75t_L g658 ( .A(n_596), .Y(n_658) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g724 ( .A(n_598), .Y(n_724) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g711 ( .A(n_600), .Y(n_711) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g712 ( .A(n_603), .Y(n_712) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g613 ( .A(n_604), .Y(n_613) );
AND2x2_ASAP7_75t_L g731 ( .A(n_604), .B(n_616), .Y(n_731) );
AND2x2_ASAP7_75t_L g794 ( .A(n_604), .B(n_726), .Y(n_794) );
AND2x2_ASAP7_75t_L g723 ( .A(n_605), .B(n_643), .Y(n_723) );
INVx1_ASAP7_75t_L g734 ( .A(n_605), .Y(n_734) );
AND2x2_ASAP7_75t_L g751 ( .A(n_605), .B(n_698), .Y(n_751) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_614), .B2(n_618), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_610), .A2(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g655 ( .A(n_613), .B(n_616), .Y(n_655) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g758 ( .A(n_616), .B(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g721 ( .A(n_619), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_620), .Y(n_649) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_621), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g694 ( .A(n_621), .Y(n_694) );
AND2x2_ASAP7_75t_L g792 ( .A(n_621), .B(n_689), .Y(n_792) );
INVx1_ASAP7_75t_L g747 ( .A(n_622), .Y(n_747) );
INVx1_ASAP7_75t_L g653 ( .A(n_624), .Y(n_653) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g742 ( .A(n_625), .Y(n_742) );
INVx4_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI32xp33_ASAP7_75t_L g722 ( .A1(n_629), .A2(n_723), .A3(n_724), .B1(n_725), .B2(n_726), .Y(n_722) );
AND2x2_ASAP7_75t_L g717 ( .A(n_630), .B(n_632), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_SL g780 ( .A1(n_630), .A2(n_781), .B(n_782), .C(n_784), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_632), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g784 ( .A(n_632), .Y(n_784) );
AND2x2_ASAP7_75t_L g638 ( .A(n_633), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g765 ( .A(n_633), .Y(n_765) );
AND2x2_ASAP7_75t_L g771 ( .A(n_633), .B(n_658), .Y(n_771) );
NOR3x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_652), .C(n_670), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_647), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
AND2x2_ASAP7_75t_L g660 ( .A(n_643), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g703 ( .A(n_643), .B(n_668), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_643), .B(n_689), .Y(n_730) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_651), .B(n_658), .Y(n_757) );
INVx2_ASAP7_75t_L g779 ( .A(n_651), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_656), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_653), .A2(n_744), .B1(n_748), .B2(n_750), .C(n_755), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_654), .A2(n_774), .B1(n_775), .B2(n_778), .Y(n_773) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B1(n_662), .B2(n_664), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x2_ASAP7_75t_L g702 ( .A(n_658), .B(n_678), .Y(n_702) );
INVx1_ASAP7_75t_L g708 ( .A(n_658), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_658), .B(n_676), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_661), .B(n_729), .Y(n_795) );
NAND2x1_ASAP7_75t_L g778 ( .A(n_662), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_663), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2x1_ASAP7_75t_SL g781 ( .A(n_666), .B(n_668), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_666), .B(n_766), .Y(n_787) );
OR2x2_ASAP7_75t_L g748 ( .A(n_667), .B(n_749), .Y(n_748) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g783 ( .A(n_668), .B(n_709), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_677), .Y(n_670) );
OAI21xp33_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_673), .B(n_676), .Y(n_671) );
OR2x2_ASAP7_75t_L g735 ( .A(n_674), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g769 ( .A(n_675), .B(n_767), .Y(n_769) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_676), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g725 ( .A(n_676), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_681), .Y(n_677) );
AND2x2_ASAP7_75t_L g710 ( .A(n_678), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_727), .Y(n_684) );
NOR3xp33_ASAP7_75t_SL g685 ( .A(n_686), .B(n_704), .C(n_719), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_692), .B(n_695), .C(n_699), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g753 ( .A(n_698), .Y(n_753) );
AND2x2_ASAP7_75t_L g766 ( .A(n_698), .B(n_767), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g774 ( .A(n_700), .Y(n_774) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_712), .B(n_713), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_709), .B2(n_710), .Y(n_705) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_706), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_717), .B2(n_718), .Y(n_713) );
INVx1_ASAP7_75t_SL g720 ( .A(n_718), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_724), .B(n_765), .Y(n_764) );
OAI22xp33_ASAP7_75t_SL g790 ( .A1(n_725), .A2(n_791), .B1(n_793), .B2(n_795), .Y(n_790) );
AOI211x1_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_732), .B(n_733), .C(n_743), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_745), .A2(n_786), .B(n_788), .Y(n_785) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g754 ( .A(n_749), .Y(n_754) );
NOR2xp67_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_752), .B(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND4xp25_ASAP7_75t_L g761 ( .A(n_762), .B(n_772), .C(n_785), .D(n_789), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_770), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_780), .Y(n_772) );
INVxp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVxp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
CKINVDCx11_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
CKINVDCx8_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
endmodule