module fake_jpeg_6463_n_245 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_30),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_20),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_47),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_20),
.C(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_21),
.B1(n_17),
.B2(n_29),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_21),
.B1(n_17),
.B2(n_29),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_35),
.B1(n_34),
.B2(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_65),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_71),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_58),
.B1(n_60),
.B2(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_80),
.Y(n_88)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_50),
.B1(n_45),
.B2(n_44),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_33),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_90),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_76),
.B1(n_79),
.B2(n_59),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_85),
.B(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_41),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_94),
.C(n_88),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_61),
.B(n_62),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_94),
.B(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_106),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_14),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_59),
.C(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_79),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_75),
.B1(n_72),
.B2(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_109),
.A2(n_112),
.B1(n_100),
.B2(n_87),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_39),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_75),
.B1(n_72),
.B2(n_77),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_120),
.B1(n_74),
.B2(n_52),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_127),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_118),
.B(n_121),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_33),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_45),
.B1(n_44),
.B2(n_42),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_14),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_49),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_124),
.B(n_25),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_65),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_87),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_92),
.C(n_90),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.C(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_41),
.C(n_48),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_52),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_45),
.B(n_66),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_149),
.B(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_121),
.B(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_57),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_33),
.B(n_39),
.C(n_64),
.D(n_15),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_153),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_15),
.B(n_25),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_33),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_106),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_150),
.C(n_133),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_163),
.C(n_175),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_115),
.B(n_111),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_147),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_109),
.C(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_176),
.B(n_166),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_126),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_152),
.C(n_141),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_131),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_135),
.B1(n_139),
.B2(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_190),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_185),
.B(n_184),
.CI(n_197),
.CON(n_210),
.SN(n_210)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_122),
.B1(n_121),
.B2(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_137),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_148),
.B(n_138),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_162),
.B(n_164),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_138),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_193),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_129),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_198),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_39),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_128),
.C(n_95),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_187),
.B(n_185),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_15),
.B(n_25),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_194),
.B1(n_182),
.B2(n_173),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_181),
.B1(n_191),
.B2(n_178),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_182),
.B1(n_170),
.B2(n_168),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_162),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_180),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_214),
.B(n_10),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_160),
.B(n_68),
.C(n_11),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_160),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_25),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_220),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_219),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_25),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_204),
.Y(n_228)
);

OA21x2_ASAP7_75t_SL g222 ( 
.A1(n_218),
.A2(n_207),
.B(n_209),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_223),
.B(n_226),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_203),
.B1(n_216),
.B2(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_9),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_225),
.B(n_228),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_0),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.CI(n_12),
.CON(n_242),
.SN(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_13),
.B(n_12),
.C(n_11),
.D(n_3),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_242),
.B(n_1),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_3),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_244),
.Y(n_245)
);


endmodule