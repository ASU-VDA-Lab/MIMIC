module fake_jpeg_5634_n_97 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_97);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_97;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_25),
.B(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_2),
.Y(n_38)
);

CKINVDCx12_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_2),
.Y(n_56)
);

XNOR2x1_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_16),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_39),
.C(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_15),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_14),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_53),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B1(n_19),
.B2(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_60),
.B1(n_65),
.B2(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_36),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_70),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_35),
.C(n_44),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_71),
.C(n_76),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_38),
.B(n_50),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_75),
.B(n_64),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_52),
.B(n_45),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_51),
.C(n_43),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_66),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_47),
.C(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_66),
.A3(n_54),
.B1(n_62),
.B2(n_60),
.C1(n_56),
.C2(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_69),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_71),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_34),
.B1(n_40),
.B2(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_78),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_89),
.A3(n_86),
.B1(n_83),
.B2(n_78),
.C1(n_79),
.C2(n_77),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_92),
.B(n_88),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_94),
.A3(n_88),
.B1(n_76),
.B2(n_40),
.C1(n_7),
.C2(n_9),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);


endmodule