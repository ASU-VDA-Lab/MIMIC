module fake_jpeg_9517_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_1),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_20),
.B1(n_29),
.B2(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_64),
.B1(n_70),
.B2(n_34),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_63),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_33),
.B1(n_44),
.B2(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_32),
.B1(n_20),
.B2(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_34),
.B1(n_25),
.B2(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_22),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_32),
.B1(n_20),
.B2(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_35),
.B1(n_21),
.B2(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_78),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_18),
.B1(n_36),
.B2(n_37),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_46),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_6),
.Y(n_124)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_101),
.B1(n_33),
.B2(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_41),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_46),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_2),
.C(n_6),
.Y(n_122)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_91),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_88),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_46),
.CI(n_40),
.CON(n_89),
.SN(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_17),
.B1(n_35),
.B2(n_21),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_31),
.B(n_27),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_46),
.B(n_44),
.C(n_17),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_36),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_37),
.Y(n_104)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_109),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_113),
.B1(n_85),
.B2(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_37),
.B1(n_31),
.B2(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_27),
.B(n_4),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_124),
.B(n_94),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_27),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_82),
.C(n_74),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_128),
.B(n_110),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_80),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_123),
.B(n_14),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_102),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_128),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_89),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_147),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_135),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_132),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_140),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_81),
.B(n_79),
.C(n_92),
.Y(n_139)
);

XOR2x1_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_154),
.Y(n_174)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_73),
.B1(n_71),
.B2(n_86),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_100),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_155),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_112),
.B(n_125),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_13),
.C(n_15),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_116),
.B(n_106),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_72),
.C(n_87),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_127),
.B1(n_124),
.B2(n_103),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_139),
.B1(n_164),
.B2(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_15),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_176),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_115),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_168),
.B(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_116),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_173),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_149),
.B(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_170),
.B(n_167),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_188),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_183),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_147),
.B1(n_166),
.B2(n_137),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_185),
.B1(n_194),
.B2(n_195),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_142),
.B1(n_143),
.B2(n_137),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_187),
.C(n_193),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_131),
.C(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_132),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_141),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_94),
.B1(n_83),
.B2(n_88),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_83),
.B1(n_7),
.B2(n_8),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_6),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_7),
.B(n_8),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_173),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_203),
.B1(n_184),
.B2(n_189),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_157),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_212),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_172),
.B1(n_167),
.B2(n_178),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_168),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_163),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVxp33_ASAP7_75t_SL g211 ( 
.A(n_181),
.Y(n_211)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_156),
.B(n_161),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_196),
.B1(n_189),
.B2(n_179),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_217),
.B1(n_223),
.B2(n_215),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_199),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_204),
.C(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_229),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_206),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_231),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_213),
.B1(n_218),
.B2(n_216),
.Y(n_227)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_195),
.B1(n_198),
.B2(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

NAND4xp25_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_156),
.C(n_190),
.D(n_209),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_204),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_232),
.A2(n_217),
.B1(n_223),
.B2(n_10),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_7),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_231),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_228),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_224),
.B1(n_232),
.B2(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_225),
.C(n_238),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_246),
.B(n_9),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_242),
.B(n_236),
.C(n_12),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.C(n_245),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_12),
.Y(n_251)
);


endmodule