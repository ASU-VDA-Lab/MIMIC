module fake_jpeg_24118_n_317 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_39),
.B(n_8),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_40),
.B(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_38),
.B1(n_42),
.B2(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_8),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_36),
.B1(n_15),
.B2(n_19),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_35),
.C(n_26),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_26),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_38),
.B1(n_53),
.B2(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_81),
.B1(n_44),
.B2(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_88),
.B(n_91),
.Y(n_130)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_82),
.B1(n_74),
.B2(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_45),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_38),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_99),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_66),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_103),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_16),
.C(n_26),
.Y(n_116)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_16),
.B1(n_14),
.B2(n_26),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_109),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_64),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_111),
.Y(n_134)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_116),
.B1(n_67),
.B2(n_85),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_99),
.B(n_93),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_97),
.B(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_113),
.Y(n_141)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_124),
.B1(n_127),
.B2(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_92),
.Y(n_143)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_16),
.B1(n_14),
.B2(n_26),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_95),
.B1(n_105),
.B2(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_47),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_144),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_112),
.B(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_146),
.B1(n_148),
.B2(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_147),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_149),
.C(n_85),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_91),
.B1(n_88),
.B2(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_63),
.B1(n_76),
.B2(n_65),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_35),
.C(n_50),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_49),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_63),
.B1(n_65),
.B2(n_100),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_14),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_41),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_70),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_108),
.B1(n_115),
.B2(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_171),
.B1(n_184),
.B2(n_145),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_168),
.B(n_170),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_127),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_125),
.B(n_19),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_128),
.B1(n_83),
.B2(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_120),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_181),
.C(n_183),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_120),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_146),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_139),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_107),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_113),
.C(n_109),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_69),
.B1(n_109),
.B2(n_34),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_191),
.Y(n_224)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_208),
.C(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_132),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_152),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_199),
.B(n_205),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_199),
.B1(n_189),
.B2(n_206),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_145),
.B(n_153),
.Y(n_199)
);

NOR4xp25_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_153),
.C(n_147),
.D(n_148),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_69),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_1),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_171),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_34),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_174),
.B1(n_177),
.B2(n_166),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_215),
.B1(n_227),
.B2(n_22),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_220),
.C(n_221),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_175),
.B1(n_159),
.B2(n_167),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_68),
.C(n_32),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_68),
.C(n_32),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_1),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_24),
.B1(n_15),
.B2(n_22),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_190),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_233),
.Y(n_258)
);

AO21x2_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_194),
.B(n_197),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_215),
.B1(n_219),
.B2(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_208),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_189),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_250),
.C(n_231),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_196),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_249),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_194),
.B1(n_200),
.B2(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_23),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_248),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_211),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_28),
.C(n_25),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_264),
.Y(n_272)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_228),
.C(n_214),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_216),
.B1(n_225),
.B2(n_227),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_225),
.C(n_27),
.Y(n_263)
);

OAI221xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_28),
.B1(n_11),
.B2(n_12),
.C(n_6),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_23),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_240),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_234),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_232),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_241),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_236),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_11),
.C(n_13),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_281),
.B(n_12),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_253),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_12),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_252),
.B1(n_257),
.B2(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_291),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_265),
.B1(n_259),
.B2(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_290),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_280),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_10),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_13),
.B(n_6),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_8),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_13),
.CI(n_7),
.CON(n_294),
.SN(n_294)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_27),
.B1(n_18),
.B2(n_25),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_300),
.C(n_9),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_28),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_9),
.B(n_4),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_283),
.C(n_292),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_307),
.B(n_308),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_305),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_18),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_18),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_18),
.B(n_25),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_298),
.C(n_301),
.Y(n_311)
);

O2A1O1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_302),
.B(n_294),
.C(n_23),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_310),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_3),
.C(n_4),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_3),
.C(n_4),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_3),
.B(n_4),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_3),
.B(n_23),
.Y(n_317)
);


endmodule