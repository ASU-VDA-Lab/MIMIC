module fake_jpeg_20762_n_19 (n_0, n_3, n_2, n_1, n_19);

input n_0;
input n_3;
input n_2;
input n_1;

output n_19;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_18;
wire n_4;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

AOI22xp33_ASAP7_75t_SL g4 ( 
.A1(n_2),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_0),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_9),
.B(n_10),
.Y(n_12)
);

O2A1O1Ixp33_ASAP7_75t_L g10 ( 
.A1(n_6),
.A2(n_1),
.B(n_3),
.C(n_0),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_13)
);

XNOR2x1_ASAP7_75t_SL g14 ( 
.A(n_13),
.B(n_3),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_15),
.C(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

AOI221xp5_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_12),
.B1(n_5),
.B2(n_11),
.C(n_15),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_0),
.B(n_8),
.Y(n_18)
);

BUFx24_ASAP7_75t_SL g19 ( 
.A(n_18),
.Y(n_19)
);


endmodule