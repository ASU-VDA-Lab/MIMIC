module real_jpeg_18280_n_21 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_21);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_21;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_66),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_SL g79 ( 
.A(n_2),
.B(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_5),
.C(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_15),
.C(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_6),
.B(n_55),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_22),
.B1(n_42),
.B2(n_46),
.C(n_48),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_14),
.C(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_9),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_35),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_17),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_17),
.B(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_31),
.C(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

AOI31xp33_ASAP7_75t_L g74 ( 
.A1(n_20),
.A2(n_36),
.A3(n_58),
.B(n_72),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.C(n_39),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_36),
.C(n_37),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.C(n_35),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.C(n_33),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_57),
.B(n_71),
.C(n_74),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_49),
.B(n_78),
.C(n_80),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_76),
.B(n_77),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B(n_75),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_70),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B(n_69),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);


endmodule