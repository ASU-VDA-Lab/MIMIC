module fake_jpeg_11206_n_595 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_595);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_595;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_71),
.Y(n_125)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_62),
.B(n_69),
.Y(n_204)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_14),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_81),
.Y(n_188)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_84),
.Y(n_162)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_85),
.Y(n_150)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g202 ( 
.A(n_89),
.Y(n_202)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_102),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_114),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_19),
.B(n_15),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_20),
.Y(n_120)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_124),
.Y(n_157)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_54),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_29),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_169),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_69),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_128),
.B(n_136),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_29),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g215 ( 
.A(n_142),
.Y(n_215)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_102),
.Y(n_144)
);

CKINVDCx12_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_145),
.B(n_194),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_101),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_148),
.B(n_174),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_75),
.A2(n_55),
.B1(n_54),
.B2(n_52),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_149),
.A2(n_107),
.B1(n_89),
.B2(n_84),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_110),
.A2(n_27),
.B1(n_49),
.B2(n_34),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_44),
.B1(n_33),
.B2(n_52),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_61),
.B(n_27),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_111),
.B(n_30),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_176),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_77),
.B(n_49),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_65),
.B(n_25),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_113),
.B(n_25),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_191),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_115),
.B(n_34),
.Y(n_191)
);

BUFx4f_ASAP7_75t_SL g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_66),
.B(n_30),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_59),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_197),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_95),
.B(n_59),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_15),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_14),
.Y(n_265)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_146),
.A2(n_35),
.B(n_24),
.C(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_208),
.B(n_246),
.Y(n_279)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_212),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_145),
.A2(n_83),
.B1(n_94),
.B2(n_79),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_213),
.A2(n_223),
.B1(n_236),
.B2(n_202),
.Y(n_290)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_214),
.Y(n_325)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_216),
.Y(n_303)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_217),
.Y(n_307)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_220),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_186),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_221),
.B(n_249),
.Y(n_282)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_222),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_80),
.B1(n_44),
.B2(n_37),
.Y(n_223)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_226),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_204),
.B1(n_197),
.B2(n_146),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_228),
.A2(n_232),
.B1(n_244),
.B2(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_230),
.A2(n_199),
.B1(n_184),
.B2(n_151),
.Y(n_324)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_149),
.A2(n_46),
.B1(n_37),
.B2(n_35),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_143),
.Y(n_233)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_233),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_127),
.A2(n_46),
.B1(n_32),
.B2(n_55),
.Y(n_236)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

CKINVDCx12_ASAP7_75t_R g238 ( 
.A(n_135),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_238),
.Y(n_297)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_167),
.A2(n_55),
.B1(n_54),
.B2(n_3),
.Y(n_244)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_137),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_247),
.Y(n_310)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_131),
.B(n_55),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_157),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_154),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_268),
.B1(n_202),
.B2(n_162),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_186),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_125),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_259),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_262),
.Y(n_289)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_204),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_264),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_265),
.B(n_266),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_142),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_195),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_267),
.A2(n_276),
.B1(n_244),
.B2(n_232),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_134),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_275),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_140),
.B(n_7),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_150),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_272),
.B(n_273),
.Y(n_326)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_274),
.B(n_201),
.Y(n_327)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_165),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_159),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_213),
.A2(n_171),
.B1(n_175),
.B2(n_178),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_227),
.A2(n_234),
.B(n_235),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_288),
.B(n_322),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_290),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_220),
.A2(n_162),
.B1(n_138),
.B2(n_132),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_285),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_209),
.B(n_158),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_299),
.B(n_304),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_224),
.B(n_153),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_306),
.B(n_313),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_243),
.A2(n_138),
.B1(n_132),
.B2(n_168),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_312),
.A2(n_324),
.B1(n_262),
.B2(n_206),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_229),
.B(n_188),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_249),
.C(n_242),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_255),
.C(n_251),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_190),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_316),
.A2(n_317),
.B(n_329),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_215),
.B(n_129),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_208),
.B(n_164),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_319),
.B(n_330),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_231),
.A2(n_171),
.B1(n_179),
.B2(n_196),
.Y(n_322)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g329 ( 
.A(n_221),
.B(n_193),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_210),
.B(n_8),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_256),
.B(n_201),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_253),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_237),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_341),
.Y(n_383)
);

INVx6_ASAP7_75t_SL g336 ( 
.A(n_297),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_336),
.Y(n_407)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_337),
.Y(n_412)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_318),
.A2(n_215),
.B(n_216),
.C(n_236),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_338),
.A2(n_349),
.B(n_286),
.Y(n_391)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_340),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_326),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_342),
.B(n_365),
.C(n_371),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_282),
.A2(n_223),
.B(n_268),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_343),
.A2(n_360),
.B(n_286),
.Y(n_402)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_308),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_350),
.Y(n_398)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_318),
.A2(n_240),
.B(n_225),
.Y(n_349)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

OAI22x1_ASAP7_75t_SL g353 ( 
.A1(n_284),
.A2(n_259),
.B1(n_253),
.B2(n_219),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_353),
.A2(n_359),
.B1(n_290),
.B2(n_317),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_359),
.B1(n_368),
.B2(n_348),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_217),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_358),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_284),
.A2(n_245),
.B1(n_257),
.B2(n_9),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_282),
.A2(n_9),
.B(n_319),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_301),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_363),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_314),
.C(n_282),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_367),
.A2(n_372),
.B1(n_302),
.B2(n_277),
.Y(n_404)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_369),
.Y(n_396)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_316),
.B(n_293),
.C(n_300),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_374),
.Y(n_397)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_287),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_292),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_376),
.Y(n_401)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_296),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_316),
.B(n_306),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_333),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_312),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_379),
.B(n_385),
.C(n_405),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_380),
.A2(n_382),
.B1(n_395),
.B2(n_404),
.Y(n_428)
);

OAI32xp33_ASAP7_75t_L g381 ( 
.A1(n_378),
.A2(n_303),
.A3(n_285),
.B1(n_324),
.B2(n_283),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_388),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_323),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_317),
.Y(n_385)
);

AOI32xp33_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_329),
.A3(n_334),
.B1(n_303),
.B2(n_310),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_387),
.B(n_339),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_377),
.A2(n_285),
.B1(n_309),
.B2(n_325),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_402),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_377),
.A2(n_291),
.B1(n_331),
.B2(n_333),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_399),
.Y(n_421)
);

OAI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_370),
.A2(n_302),
.B1(n_277),
.B2(n_296),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_370),
.A2(n_321),
.B1(n_331),
.B2(n_298),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_367),
.A2(n_298),
.B1(n_321),
.B2(n_328),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_414),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_375),
.C(n_344),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_344),
.B(n_286),
.C(n_328),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_357),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_409),
.B(n_339),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_340),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_397),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_380),
.A2(n_355),
.B1(n_361),
.B2(n_353),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_422),
.A2(n_434),
.B1(n_431),
.B2(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_410),
.Y(n_425)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_427),
.Y(n_453)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_349),
.B(n_355),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_432),
.A2(n_436),
.B(n_382),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_356),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_433),
.B(n_446),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_409),
.A2(n_361),
.B1(n_335),
.B2(n_343),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_364),
.Y(n_435)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

INVx13_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_438),
.Y(n_456)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_379),
.C(n_385),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_398),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_442),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_414),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_376),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_447),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_336),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_372),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_449),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_401),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_405),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_450),
.A2(n_455),
.B1(n_458),
.B2(n_424),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_428),
.A2(n_388),
.B1(n_402),
.B2(n_406),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_437),
.B(n_384),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_444),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_384),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_463),
.C(n_472),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_432),
.A2(n_401),
.B(n_381),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_468),
.B(n_475),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_420),
.A2(n_390),
.B1(n_411),
.B2(n_413),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_470),
.A2(n_445),
.B1(n_431),
.B2(n_424),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_430),
.B(n_390),
.C(n_393),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_393),
.C(n_412),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_435),
.C(n_447),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_433),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_373),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_476),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_430),
.B(n_338),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_478),
.Y(n_482)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_467),
.Y(n_480)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_477),
.Y(n_483)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_477),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_488),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_442),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_485),
.Y(n_526)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_486),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_451),
.B(n_416),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_455),
.A2(n_420),
.B1(n_418),
.B2(n_423),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_489),
.A2(n_470),
.B1(n_454),
.B2(n_460),
.Y(n_508)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_492),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_425),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_471),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_497),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_431),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_494),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_453),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_452),
.B(n_429),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_457),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_468),
.A2(n_417),
.B(n_422),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_505),
.Y(n_512)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_466),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_499),
.A2(n_504),
.B1(n_457),
.B2(n_456),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_473),
.C(n_463),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_503),
.A2(n_479),
.B1(n_460),
.B2(n_454),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_462),
.B(n_354),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_521),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_508),
.A2(n_503),
.B1(n_497),
.B2(n_482),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_461),
.C(n_458),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_510),
.B(n_518),
.C(n_522),
.Y(n_538)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_513),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_480),
.A2(n_479),
.B1(n_450),
.B2(n_421),
.Y(n_517)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_517),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_500),
.B(n_465),
.C(n_478),
.Y(n_518)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_519),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_478),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_443),
.C(n_439),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_419),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_481),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_525),
.Y(n_529)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_529),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_524),
.Y(n_554)
);

AOI321xp33_ASAP7_75t_L g533 ( 
.A1(n_514),
.A2(n_486),
.A3(n_487),
.B1(n_485),
.B2(n_483),
.C(n_490),
.Y(n_533)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_518),
.A2(n_487),
.B(n_493),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_543),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_501),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_536),
.B(n_542),
.Y(n_553)
);

OAI321xp33_ASAP7_75t_L g537 ( 
.A1(n_520),
.A2(n_488),
.A3(n_496),
.B1(n_495),
.B2(n_484),
.C(n_491),
.Y(n_537)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_537),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_508),
.A2(n_509),
.B1(n_506),
.B2(n_515),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_540),
.A2(n_541),
.B1(n_526),
.B2(n_516),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_411),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_507),
.B(n_482),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_510),
.B(n_499),
.C(n_469),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_519),
.Y(n_556)
);

BUFx12_ASAP7_75t_L g545 ( 
.A(n_516),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_545),
.B(n_469),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_534),
.A2(n_531),
.B1(n_530),
.B2(n_527),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_546),
.A2(n_550),
.B1(n_539),
.B2(n_554),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_512),
.C(n_517),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_547),
.A2(n_549),
.B(n_555),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_512),
.C(n_521),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_541),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_551),
.B(n_554),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_538),
.B(n_527),
.C(n_519),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_556),
.B(n_558),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_511),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_560),
.Y(n_566)
);

OAI21xp33_ASAP7_75t_L g561 ( 
.A1(n_559),
.A2(n_557),
.B(n_533),
.Y(n_561)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_561),
.Y(n_573)
);

FAx1_ASAP7_75t_SL g562 ( 
.A(n_555),
.B(n_545),
.CI(n_532),
.CON(n_562),
.SN(n_562)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_567),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_528),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_565),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_558),
.B(n_528),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_529),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_569),
.B(n_552),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_549),
.A2(n_545),
.B(n_419),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_570),
.A2(n_421),
.B(n_352),
.Y(n_578)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_574),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_561),
.A2(n_550),
.B1(n_548),
.B2(n_459),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_575),
.B(n_577),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_413),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_564),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_568),
.B(n_337),
.C(n_399),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_579),
.B(n_571),
.Y(n_583)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_580),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_572),
.B(n_573),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_582),
.A2(n_585),
.B(n_563),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_583),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_579),
.A2(n_562),
.B1(n_564),
.B2(n_571),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_581),
.Y(n_589)
);

OAI321xp33_ASAP7_75t_L g591 ( 
.A1(n_589),
.A2(n_590),
.A3(n_587),
.B1(n_580),
.B2(n_576),
.C(n_565),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_586),
.B(n_584),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_576),
.C(n_427),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_SL g593 ( 
.A1(n_592),
.A2(n_427),
.B(n_438),
.C(n_374),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_593),
.A2(n_438),
.B1(n_351),
.B2(n_369),
.Y(n_594)
);

BUFx24_ASAP7_75t_SL g595 ( 
.A(n_594),
.Y(n_595)
);


endmodule