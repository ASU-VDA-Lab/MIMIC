module real_aes_15675_n_361 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_361);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_361;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1802;
wire n_727;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1323;
wire n_1280;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g760 ( .A(n_0), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g1150 ( .A1(n_1), .A2(n_321), .B1(n_588), .B2(n_878), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g1172 ( .A(n_1), .Y(n_1172) );
INVx1_ASAP7_75t_L g1327 ( .A(n_2), .Y(n_1327) );
AO22x1_ASAP7_75t_L g1361 ( .A1(n_2), .A2(n_236), .B1(n_643), .B2(n_1267), .Y(n_1361) );
INVx1_ASAP7_75t_L g377 ( .A(n_3), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_3), .B(n_387), .Y(n_410) );
AND2x2_ASAP7_75t_L g627 ( .A(n_3), .B(n_255), .Y(n_627) );
AND2x2_ASAP7_75t_L g645 ( .A(n_3), .B(n_531), .Y(n_645) );
INVx1_ASAP7_75t_L g1337 ( .A(n_4), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_4), .A2(n_123), .B1(n_547), .B2(n_798), .Y(n_1360) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_5), .A2(n_325), .B1(n_762), .B2(n_878), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g938 ( .A1(n_5), .A2(n_7), .B1(n_648), .B2(n_655), .C(n_939), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_6), .A2(n_42), .B1(n_588), .B2(n_592), .Y(n_587) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_6), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g928 ( .A1(n_7), .A2(n_13), .B1(n_604), .B2(n_709), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_8), .A2(n_319), .B1(n_876), .B2(n_878), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_8), .A2(n_264), .B1(n_783), .B2(n_831), .C(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_9), .A2(n_201), .B1(n_597), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_9), .A2(n_181), .B1(n_786), .B2(n_787), .Y(n_785) );
XOR2x2_ASAP7_75t_L g392 ( .A(n_10), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g969 ( .A(n_11), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_11), .A2(n_352), .B1(n_632), .B2(n_636), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g1769 ( .A(n_12), .Y(n_1769) );
A2O1A1Ixp33_ASAP7_75t_L g948 ( .A1(n_13), .A2(n_729), .B(n_949), .C(n_955), .Y(n_948) );
INVx1_ASAP7_75t_L g1530 ( .A(n_14), .Y(n_1530) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_14), .A2(n_221), .B1(n_1541), .B2(n_1555), .Y(n_1554) );
AOI22xp33_ASAP7_75t_SL g1459 ( .A1(n_15), .A2(n_230), .B1(n_767), .B2(n_1460), .Y(n_1459) );
INVxp67_ASAP7_75t_SL g1483 ( .A(n_15), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_16), .A2(n_312), .B1(n_799), .B2(n_821), .C(n_823), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_16), .A2(n_336), .B1(n_596), .B2(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_17), .A2(n_92), .B1(n_1541), .B2(n_1545), .Y(n_1575) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_18), .A2(n_338), .B1(n_833), .B2(n_942), .Y(n_1224) );
INVx1_ASAP7_75t_L g1243 ( .A(n_18), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1638 ( .A1(n_19), .A2(n_345), .B1(n_1548), .B2(n_1551), .Y(n_1638) );
INVx2_ASAP7_75t_L g445 ( .A(n_20), .Y(n_445) );
OAI22xp5_ASAP7_75t_SL g1043 ( .A1(n_21), .A2(n_285), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_21), .A2(n_285), .B1(n_673), .B2(n_675), .C(n_1057), .Y(n_1056) );
XNOR2x1_ASAP7_75t_L g1015 ( .A(n_22), .B(n_1016), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1779 ( .A1(n_23), .A2(n_119), .B1(n_711), .B2(n_1116), .Y(n_1779) );
AOI22xp33_ASAP7_75t_L g1793 ( .A1(n_23), .A2(n_167), .B1(n_827), .B2(n_904), .Y(n_1793) );
INVx1_ASAP7_75t_L g1494 ( .A(n_24), .Y(n_1494) );
OAI222xp33_ASAP7_75t_L g1515 ( .A1(n_24), .A2(n_170), .B1(n_725), .B2(n_1170), .C1(n_1516), .C2(n_1521), .Y(n_1515) );
INVx1_ASAP7_75t_L g1436 ( .A(n_25), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_26), .A2(n_270), .B1(n_657), .B2(n_660), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_26), .A2(n_265), .B1(n_588), .B2(n_858), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_27), .A2(n_263), .B1(n_606), .B2(n_613), .Y(n_1154) );
INVx1_ASAP7_75t_L g1167 ( .A(n_27), .Y(n_1167) );
AOI22xp5_ASAP7_75t_L g1547 ( .A1(n_28), .A2(n_226), .B1(n_1548), .B2(n_1551), .Y(n_1547) );
INVx1_ASAP7_75t_L g1108 ( .A(n_29), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_30), .A2(n_127), .B1(n_597), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_30), .A2(n_295), .B1(n_737), .B2(n_738), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g1788 ( .A1(n_31), .A2(n_219), .B1(n_613), .B2(n_719), .Y(n_1788) );
INVx1_ASAP7_75t_L g1795 ( .A(n_31), .Y(n_1795) );
AOI22xp33_ASAP7_75t_SL g1783 ( .A1(n_32), .A2(n_84), .B1(n_709), .B2(n_1778), .Y(n_1783) );
AOI22xp33_ASAP7_75t_SL g1801 ( .A1(n_32), .A2(n_247), .B1(n_1802), .B2(n_1803), .Y(n_1801) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_33), .Y(n_372) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_33), .B(n_370), .Y(n_1542) );
INVx1_ASAP7_75t_L g1055 ( .A(n_34), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1636 ( .A1(n_35), .A2(n_195), .B1(n_1541), .B2(n_1637), .Y(n_1636) );
OAI22xp5_ASAP7_75t_SL g1411 ( .A1(n_36), .A2(n_296), .B1(n_398), .B2(n_419), .Y(n_1411) );
INVxp67_ASAP7_75t_SL g1440 ( .A(n_36), .Y(n_1440) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_37), .Y(n_1445) );
INVxp67_ASAP7_75t_L g869 ( .A(n_38), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_38), .A2(n_218), .B1(n_1541), .B2(n_1545), .Y(n_1589) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_39), .A2(n_336), .B1(n_657), .B2(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_39), .A2(n_312), .B1(n_853), .B2(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g1512 ( .A(n_40), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_41), .A2(n_91), .B1(n_771), .B2(n_773), .Y(n_924) );
AOI221xp5_ASAP7_75t_L g950 ( .A1(n_41), .A2(n_206), .B1(n_898), .B2(n_951), .C(n_952), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_42), .A2(n_97), .B1(n_648), .B2(n_650), .C(n_654), .Y(n_647) );
INVx1_ASAP7_75t_L g1227 ( .A(n_43), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_44), .A2(n_284), .B1(n_882), .B2(n_1079), .Y(n_1457) );
INVx1_ASAP7_75t_L g1476 ( .A(n_44), .Y(n_1476) );
OAI21xp5_ASAP7_75t_L g837 ( .A1(n_45), .A2(n_838), .B(n_839), .Y(n_837) );
NAND5xp2_ASAP7_75t_L g1259 ( .A(n_46), .B(n_1260), .C(n_1283), .D(n_1292), .E(n_1300), .Y(n_1259) );
INVx1_ASAP7_75t_L g1308 ( .A(n_46), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_47), .A2(n_146), .B1(n_632), .B2(n_636), .Y(n_1157) );
OAI211xp5_ASAP7_75t_SL g1159 ( .A1(n_47), .A2(n_936), .B(n_1160), .C(n_1165), .Y(n_1159) );
INVx1_ASAP7_75t_L g1226 ( .A(n_48), .Y(n_1226) );
INVx1_ASAP7_75t_L g1511 ( .A(n_49), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_50), .A2(n_187), .B1(n_900), .B2(n_904), .Y(n_974) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_50), .A2(n_330), .B1(n_588), .B2(n_999), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_51), .A2(n_165), .B1(n_1541), .B2(n_1545), .Y(n_1562) );
INVxp67_ASAP7_75t_L g1767 ( .A(n_51), .Y(n_1767) );
AOI22xp5_ASAP7_75t_L g1808 ( .A1(n_51), .A2(n_1809), .B1(n_1812), .B2(n_1817), .Y(n_1808) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_52), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_53), .A2(n_54), .B1(n_588), .B2(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g794 ( .A(n_53), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_54), .A2(n_137), .B1(n_781), .B2(n_783), .C(n_784), .Y(n_780) );
XOR2x2_ASAP7_75t_L g961 ( .A(n_55), .B(n_962), .Y(n_961) );
XOR2xp5_ASAP7_75t_L g1142 ( .A(n_56), .B(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1453 ( .A(n_57), .Y(n_1453) );
AOI22xp33_ASAP7_75t_SL g1151 ( .A1(n_58), .A2(n_292), .B1(n_711), .B2(n_882), .Y(n_1151) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_58), .A2(n_257), .B1(n_745), .B2(n_952), .C(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1054 ( .A(n_59), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_60), .A2(n_266), .B1(n_594), .B2(n_597), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_60), .A2(n_140), .B1(n_657), .B2(n_659), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_61), .A2(n_171), .B1(n_547), .B2(n_798), .C(n_799), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_61), .A2(n_243), .B1(n_473), .B2(n_853), .Y(n_1287) );
INVx1_ASAP7_75t_L g1123 ( .A(n_62), .Y(n_1123) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_63), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_64), .A2(n_243), .B1(n_833), .B2(n_1267), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_64), .A2(n_171), .B1(n_853), .B2(n_1079), .Y(n_1286) );
INVx1_ASAP7_75t_L g416 ( .A(n_65), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_66), .A2(n_155), .B1(n_770), .B2(n_882), .Y(n_881) );
AOI21xp33_ASAP7_75t_L g907 ( .A1(n_66), .A2(n_693), .B(n_781), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_67), .A2(n_805), .B1(n_806), .B2(n_863), .Y(n_804) );
INVxp67_ASAP7_75t_SL g863 ( .A(n_67), .Y(n_863) );
INVx1_ASAP7_75t_L g920 ( .A(n_68), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g1112 ( .A1(n_69), .A2(n_291), .B1(n_588), .B2(n_709), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_69), .A2(n_309), .B1(n_657), .B2(n_659), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g1455 ( .A1(n_70), .A2(n_175), .B1(n_876), .B2(n_1042), .Y(n_1455) );
INVxp67_ASAP7_75t_SL g1482 ( .A(n_70), .Y(n_1482) );
INVx1_ASAP7_75t_L g817 ( .A(n_71), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_72), .A2(n_254), .B1(n_490), .B2(n_494), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_72), .A2(n_254), .B1(n_535), .B2(n_537), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_73), .Y(n_886) );
OAI21xp5_ASAP7_75t_SL g911 ( .A1(n_74), .A2(n_632), .B(n_912), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_75), .Y(n_1274) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_76), .A2(n_264), .B1(n_604), .B2(n_767), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_76), .A2(n_319), .B1(n_787), .B2(n_904), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_77), .A2(n_97), .B1(n_592), .B2(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_77), .Y(n_686) );
INVx1_ASAP7_75t_L g819 ( .A(n_78), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_79), .A2(n_214), .B1(n_853), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_79), .A2(n_88), .B1(n_660), .B2(n_942), .Y(n_1091) );
OAI21xp5_ASAP7_75t_L g1139 ( .A1(n_80), .A2(n_632), .B(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1019 ( .A(n_81), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1414 ( .A1(n_82), .A2(n_158), .B1(n_643), .B2(n_1094), .Y(n_1414) );
INVxp67_ASAP7_75t_SL g1433 ( .A(n_82), .Y(n_1433) );
AOI22xp33_ASAP7_75t_SL g1028 ( .A1(n_83), .A2(n_287), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_83), .A2(n_90), .B1(n_746), .B2(n_831), .C(n_1050), .Y(n_1049) );
AOI221xp5_ASAP7_75t_L g1792 ( .A1(n_84), .A2(n_327), .B1(n_655), .B2(n_798), .C(n_984), .Y(n_1792) );
INVx1_ASAP7_75t_L g1484 ( .A(n_85), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_86), .A2(n_276), .B1(n_588), .B2(n_1030), .Y(n_1198) );
AOI221xp5_ASAP7_75t_L g1203 ( .A1(n_86), .A2(n_273), .B1(n_649), .B2(n_655), .C(n_823), .Y(n_1203) );
INVx1_ASAP7_75t_L g1021 ( .A(n_87), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_88), .A2(n_293), .B1(n_853), .B2(n_1079), .Y(n_1082) );
INVx1_ASAP7_75t_L g1191 ( .A(n_89), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_89), .A2(n_302), .B1(n_660), .B2(n_904), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_90), .A2(n_193), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_91), .A2(n_134), .B1(n_659), .B2(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g412 ( .A(n_93), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g1501 ( .A1(n_94), .A2(n_334), .B1(n_588), .B2(n_1030), .Y(n_1501) );
INVxp67_ASAP7_75t_SL g1506 ( .A(n_94), .Y(n_1506) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_95), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_96), .Y(n_1074) );
XNOR2xp5_ASAP7_75t_L g1216 ( .A(n_98), .B(n_1217), .Y(n_1216) );
AOI22xp5_ASAP7_75t_L g1566 ( .A1(n_99), .A2(n_225), .B1(n_1548), .B2(n_1551), .Y(n_1566) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_100), .A2(n_322), .B1(n_1114), .B2(n_1116), .Y(n_1113) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_100), .A2(n_346), .B1(n_741), .B2(n_939), .C(n_1137), .Y(n_1136) );
OAI211xp5_ASAP7_75t_L g1270 ( .A1(n_101), .A2(n_1271), .B(n_1272), .C(n_1273), .Y(n_1270) );
INVx1_ASAP7_75t_L g1304 ( .A(n_101), .Y(n_1304) );
INVx1_ASAP7_75t_L g758 ( .A(n_102), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_102), .A2(n_139), .B1(n_671), .B2(n_675), .C(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_103), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_103), .A2(n_121), .B1(n_909), .B2(n_910), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_104), .A2(n_242), .B1(n_643), .B2(n_906), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_104), .A2(n_259), .B1(n_592), .B2(n_604), .Y(n_1430) );
INVx1_ASAP7_75t_L g438 ( .A(n_105), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g1234 ( .A1(n_106), .A2(n_823), .B(n_1137), .Y(n_1234) );
INVx1_ASAP7_75t_L g1242 ( .A(n_106), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_107), .A2(n_309), .B1(n_588), .B2(n_592), .Y(n_1120) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_107), .A2(n_291), .B1(n_655), .B2(n_1050), .C(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1182 ( .A(n_108), .Y(n_1182) );
INVx1_ASAP7_75t_L g1403 ( .A(n_109), .Y(n_1403) );
INVx1_ASAP7_75t_L g763 ( .A(n_110), .Y(n_763) );
INVx1_ASAP7_75t_L g370 ( .A(n_111), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_112), .A2(n_256), .B1(n_655), .B2(n_830), .C(n_1222), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_112), .A2(n_178), .B1(n_588), .B2(n_619), .Y(n_1244) );
INVx1_ASAP7_75t_L g1070 ( .A(n_113), .Y(n_1070) );
INVx1_ASAP7_75t_L g1069 ( .A(n_114), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g1153 ( .A1(n_115), .A2(n_290), .B1(n_588), .B2(n_709), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g1174 ( .A(n_115), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_116), .A2(n_289), .B1(n_709), .B2(n_1041), .C(n_1077), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_116), .A2(n_237), .B1(n_649), .B2(n_651), .C(n_831), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_117), .A2(n_184), .B1(n_1032), .B2(n_1079), .Y(n_1456) );
INVx1_ASAP7_75t_L g1480 ( .A(n_117), .Y(n_1480) );
OAI222xp33_ASAP7_75t_L g1347 ( .A1(n_118), .A2(n_340), .B1(n_1348), .B2(n_1350), .C1(n_1352), .C2(n_1354), .Y(n_1347) );
INVx1_ASAP7_75t_L g1365 ( .A(n_118), .Y(n_1365) );
AOI21xp33_ASAP7_75t_L g1800 ( .A1(n_119), .A2(n_691), .B(n_799), .Y(n_1800) );
INVx1_ASAP7_75t_L g578 ( .A(n_120), .Y(n_578) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_120), .A2(n_122), .B1(n_671), .B2(n_675), .C(n_679), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_121), .Y(n_888) );
INVx1_ASAP7_75t_L g569 ( .A(n_122), .Y(n_569) );
INVx1_ASAP7_75t_L g1334 ( .A(n_123), .Y(n_1334) );
OAI211xp5_ASAP7_75t_L g1405 ( .A1(n_124), .A2(n_1406), .B(n_1407), .C(n_1408), .Y(n_1405) );
INVxp33_ASAP7_75t_SL g1423 ( .A(n_124), .Y(n_1423) );
CKINVDCx5p33_ASAP7_75t_R g1195 ( .A(n_125), .Y(n_1195) );
AOI22xp5_ASAP7_75t_L g1571 ( .A1(n_126), .A2(n_328), .B1(n_1548), .B2(n_1551), .Y(n_1571) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_127), .A2(n_246), .B1(n_688), .B2(n_693), .C(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_SL g977 ( .A(n_128), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_128), .A2(n_261), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
INVx1_ASAP7_75t_L g828 ( .A(n_129), .Y(n_828) );
INVx1_ASAP7_75t_L g1187 ( .A(n_130), .Y(n_1187) );
AOI21xp33_ASAP7_75t_L g1212 ( .A1(n_130), .A2(n_693), .B(n_823), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_131), .A2(n_166), .B1(n_636), .B2(n_838), .Y(n_1183) );
OAI211xp5_ASAP7_75t_L g1201 ( .A1(n_131), .A2(n_641), .B(n_1202), .C(n_1205), .Y(n_1201) );
INVx1_ASAP7_75t_L g968 ( .A(n_132), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g1009 ( .A1(n_132), .A2(n_176), .B1(n_719), .B2(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1449 ( .A(n_133), .Y(n_1449) );
OAI222xp33_ASAP7_75t_L g1472 ( .A1(n_133), .A2(n_216), .B1(n_1169), .B2(n_1473), .C1(n_1474), .C2(n_1481), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_134), .A2(n_206), .B1(n_771), .B2(n_926), .Y(n_925) );
XOR2x2_ASAP7_75t_L g700 ( .A(n_135), .B(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1540 ( .A1(n_135), .A2(n_229), .B1(n_1541), .B2(n_1545), .Y(n_1540) );
INVxp67_ASAP7_75t_SL g972 ( .A(n_136), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_136), .A2(n_205), .B1(n_597), .B2(n_1005), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_137), .A2(n_141), .B1(n_709), .B2(n_776), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_138), .A2(n_265), .B1(n_651), .B2(n_830), .C(n_831), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_138), .A2(n_270), .B1(n_588), .B2(n_619), .Y(n_851) );
INVx1_ASAP7_75t_L g757 ( .A(n_139), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_140), .A2(n_174), .B1(n_594), .B2(n_597), .Y(n_599) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_141), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g1556 ( .A1(n_142), .A2(n_241), .B1(n_1548), .B2(n_1551), .Y(n_1556) );
OA21x2_ASAP7_75t_L g1017 ( .A1(n_143), .A2(n_622), .B(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_144), .A2(n_168), .B1(n_602), .B2(n_709), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_144), .A2(n_194), .B1(n_655), .B2(n_741), .C(n_745), .Y(n_740) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_145), .A2(n_304), .B1(n_613), .B2(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g748 ( .A(n_145), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_147), .A2(n_283), .B1(n_606), .B2(n_613), .Y(n_605) );
INVx1_ASAP7_75t_L g667 ( .A(n_147), .Y(n_667) );
INVx1_ASAP7_75t_L g808 ( .A(n_148), .Y(n_808) );
INVx1_ASAP7_75t_L g1464 ( .A(n_149), .Y(n_1464) );
INVx1_ASAP7_75t_L g1772 ( .A(n_150), .Y(n_1772) );
OAI221xp5_ASAP7_75t_SL g1797 ( .A1(n_150), .A2(n_262), .B1(n_671), .B2(n_1169), .C(n_1798), .Y(n_1797) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_151), .A2(n_160), .B1(n_515), .B2(n_518), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g526 ( .A1(n_151), .A2(n_160), .B1(n_527), .B2(n_528), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_152), .A2(n_349), .B1(n_725), .B2(n_1170), .C(n_1229), .Y(n_1228) );
OAI22xp33_ASAP7_75t_L g1248 ( .A1(n_152), .A2(n_349), .B1(n_571), .B2(n_1045), .Y(n_1248) );
AO22x1_ASAP7_75t_L g873 ( .A1(n_153), .A2(n_203), .B1(n_770), .B2(n_771), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_153), .B(n_732), .Y(n_902) );
INVx1_ASAP7_75t_L g1299 ( .A(n_154), .Y(n_1299) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_155), .A2(n_203), .B1(n_657), .B2(n_900), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_156), .Y(n_721) );
INVx1_ASAP7_75t_L g504 ( .A(n_157), .Y(n_504) );
INVx1_ASAP7_75t_L g1429 ( .A(n_158), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g1156 ( .A(n_159), .Y(n_1156) );
INVx1_ASAP7_75t_L g426 ( .A(n_161), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_162), .A2(n_347), .B1(n_632), .B2(n_636), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_163), .A2(n_294), .B1(n_632), .B2(n_636), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_164), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1780 ( .A1(n_167), .A2(n_315), .B1(n_1116), .B2(n_1781), .Y(n_1780) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_168), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_169), .A2(n_191), .B1(n_632), .B2(n_636), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_169), .A2(n_641), .B(n_646), .C(n_662), .Y(n_640) );
INVx1_ASAP7_75t_L g1493 ( .A(n_170), .Y(n_1493) );
INVx1_ASAP7_75t_L g1329 ( .A(n_172), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_172), .A2(n_267), .B1(n_833), .B2(n_1267), .Y(n_1381) );
INVx1_ASAP7_75t_L g1141 ( .A(n_173), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_174), .A2(n_266), .B1(n_688), .B2(n_689), .C(n_693), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g1469 ( .A1(n_175), .A2(n_230), .B1(n_745), .B2(n_784), .C(n_1176), .Y(n_1469) );
INVx1_ASAP7_75t_L g966 ( .A(n_176), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g1409 ( .A(n_177), .Y(n_1409) );
AOI22xp33_ASAP7_75t_SL g1235 ( .A1(n_178), .A2(n_320), .B1(n_643), .B2(n_657), .Y(n_1235) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_179), .A2(n_641), .B(n_1220), .C(n_1225), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1251 ( .A1(n_179), .A2(n_343), .B1(n_636), .B2(n_838), .Y(n_1251) );
INVx1_ASAP7_75t_L g1417 ( .A(n_180), .Y(n_1417) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_181), .A2(n_278), .B1(n_770), .B2(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g1026 ( .A(n_182), .Y(n_1026) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_182), .A2(n_233), .B1(n_651), .B2(n_741), .C(n_952), .Y(n_1063) );
OAI211xp5_ASAP7_75t_L g1261 ( .A1(n_183), .A2(n_1262), .B(n_1263), .C(n_1269), .Y(n_1261) );
NOR2xp33_ASAP7_75t_L g1282 ( .A(n_183), .B(n_845), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_184), .A2(n_284), .B1(n_738), .B2(n_786), .Y(n_1470) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_185), .A2(n_237), .B1(n_1041), .B2(n_1042), .C(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_185), .A2(n_289), .B1(n_660), .B2(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g706 ( .A(n_186), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_186), .A2(n_324), .B1(n_675), .B2(n_725), .C(n_726), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_187), .A2(n_356), .B1(n_588), .B2(n_1008), .Y(n_1007) );
INVx2_ASAP7_75t_L g1544 ( .A(n_188), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_188), .B(n_303), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_188), .B(n_1550), .Y(n_1552) );
AOI22xp33_ASAP7_75t_L g1499 ( .A1(n_189), .A2(n_354), .B1(n_855), .B2(n_1002), .Y(n_1499) );
INVx1_ASAP7_75t_L g1519 ( .A(n_189), .Y(n_1519) );
AOI22xp5_ASAP7_75t_L g1561 ( .A1(n_190), .A2(n_277), .B1(n_1548), .B2(n_1551), .Y(n_1561) );
INVx1_ASAP7_75t_L g1207 ( .A(n_192), .Y(n_1207) );
INVx1_ASAP7_75t_L g1062 ( .A(n_193), .Y(n_1062) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_194), .A2(n_298), .B1(n_592), .B2(n_604), .Y(n_717) );
INVx1_ASAP7_75t_L g1129 ( .A(n_196), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_197), .A2(n_286), .B1(n_632), .B2(n_845), .Y(n_933) );
OAI211xp5_ASAP7_75t_L g935 ( .A1(n_197), .A2(n_936), .B(n_937), .C(n_943), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_198), .Y(n_894) );
XOR2x2_ASAP7_75t_L g564 ( .A(n_199), .B(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_200), .A2(n_346), .B1(n_597), .B2(n_1114), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_200), .A2(n_322), .B1(n_659), .B2(n_942), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_201), .A2(n_278), .B1(n_797), .B2(n_798), .C(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g1787 ( .A(n_202), .Y(n_1787) );
AOI22xp5_ASAP7_75t_L g1572 ( .A1(n_204), .A2(n_311), .B1(n_1541), .B2(n_1555), .Y(n_1572) );
INVxp67_ASAP7_75t_SL g980 ( .A(n_205), .Y(n_980) );
INVx1_ASAP7_75t_L g1392 ( .A(n_207), .Y(n_1392) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_208), .B(n_725), .Y(n_985) );
INVx1_ASAP7_75t_L g996 ( .A(n_208), .Y(n_996) );
INVx1_ASAP7_75t_L g1463 ( .A(n_209), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_210), .A2(n_281), .B1(n_833), .B2(n_906), .Y(n_1264) );
AOI22xp33_ASAP7_75t_SL g1288 ( .A1(n_210), .A2(n_301), .B1(n_588), .B2(n_858), .Y(n_1288) );
AOI22xp33_ASAP7_75t_SL g1192 ( .A1(n_211), .A2(n_273), .B1(n_588), .B2(n_1030), .Y(n_1192) );
AOI22xp33_ASAP7_75t_SL g1213 ( .A1(n_211), .A2(n_276), .B1(n_657), .B2(n_787), .Y(n_1213) );
INVx1_ASAP7_75t_L g1529 ( .A(n_212), .Y(n_1529) );
XNOR2xp5_ASAP7_75t_L g1810 ( .A(n_213), .B(n_1811), .Y(n_1810) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_214), .A2(n_293), .B1(n_651), .B2(n_693), .C(n_830), .Y(n_1095) );
INVx1_ASAP7_75t_L g1039 ( .A(n_215), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_215), .A2(n_275), .B1(n_833), .B2(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1450 ( .A(n_216), .Y(n_1450) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_217), .A2(n_474), .B(n_499), .C(n_503), .Y(n_498) );
INVx1_ASAP7_75t_L g553 ( .A(n_217), .Y(n_553) );
INVx1_ASAP7_75t_L g1796 ( .A(n_219), .Y(n_1796) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_220), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_222), .Y(n_1230) );
CKINVDCx5p33_ASAP7_75t_R g1277 ( .A(n_223), .Y(n_1277) );
INVx2_ASAP7_75t_L g444 ( .A(n_224), .Y(n_444) );
INVx1_ASAP7_75t_L g483 ( .A(n_224), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_224), .B(n_445), .Y(n_612) );
INVx1_ASAP7_75t_L g1342 ( .A(n_227), .Y(n_1342) );
NAND2xp33_ASAP7_75t_SL g1382 ( .A(n_227), .B(n_547), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_228), .A2(n_323), .B1(n_463), .B2(n_1032), .Y(n_1500) );
INVx1_ASAP7_75t_L g1517 ( .A(n_228), .Y(n_1517) );
AOI22xp33_ASAP7_75t_SL g1498 ( .A1(n_231), .A2(n_252), .B1(n_588), .B2(n_1008), .Y(n_1498) );
INVxp67_ASAP7_75t_SL g1522 ( .A(n_231), .Y(n_1522) );
INVx1_ASAP7_75t_L g437 ( .A(n_232), .Y(n_437) );
INVx1_ASAP7_75t_L g1037 ( .A(n_233), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_234), .A2(n_318), .B1(n_1548), .B2(n_1551), .Y(n_1574) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_235), .A2(n_308), .B1(n_1271), .B2(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1302 ( .A(n_235), .Y(n_1302) );
AOI21xp5_ASAP7_75t_L g1343 ( .A1(n_236), .A2(n_862), .B(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1386 ( .A(n_238), .Y(n_1386) );
OAI21xp5_ASAP7_75t_L g1526 ( .A1(n_239), .A2(n_838), .B(n_1527), .Y(n_1526) );
BUFx3_ASAP7_75t_L g450 ( .A(n_240), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_242), .A2(n_279), .B1(n_592), .B2(n_1029), .Y(n_1434) );
INVx1_ASAP7_75t_L g1088 ( .A(n_244), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_245), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_246), .A2(n_295), .B1(n_597), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g1777 ( .A1(n_247), .A2(n_327), .B1(n_767), .B2(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1319 ( .A(n_248), .Y(n_1319) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_248), .B(n_1322), .Y(n_1321) );
AOI21xp33_ASAP7_75t_L g1418 ( .A1(n_249), .A2(n_799), .B(n_823), .Y(n_1418) );
INVx1_ASAP7_75t_L g1428 ( .A(n_249), .Y(n_1428) );
INVx1_ASAP7_75t_L g1127 ( .A(n_250), .Y(n_1127) );
XOR2x2_ASAP7_75t_L g1398 ( .A(n_251), .B(n_1399), .Y(n_1398) );
AOI22xp5_ASAP7_75t_L g1567 ( .A1(n_251), .A2(n_268), .B1(n_1541), .B2(n_1545), .Y(n_1567) );
AOI21xp33_ASAP7_75t_L g1508 ( .A1(n_252), .A2(n_746), .B(n_831), .Y(n_1508) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_253), .A2(n_272), .B1(n_606), .B2(n_613), .Y(n_929) );
INVx1_ASAP7_75t_L g944 ( .A(n_253), .Y(n_944) );
BUFx3_ASAP7_75t_L g387 ( .A(n_255), .Y(n_387) );
INVx1_ASAP7_75t_L g531 ( .A(n_255), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_256), .A2(n_320), .B1(n_588), .B2(n_1042), .Y(n_1247) );
AOI22xp33_ASAP7_75t_SL g1152 ( .A1(n_257), .A2(n_313), .B1(n_711), .B2(n_882), .Y(n_1152) );
XNOR2x1_ASAP7_75t_L g1066 ( .A(n_258), .B(n_1067), .Y(n_1066) );
NAND2xp5_ASAP7_75t_SL g1413 ( .A(n_259), .B(n_823), .Y(n_1413) );
INVxp67_ASAP7_75t_SL g1775 ( .A(n_260), .Y(n_1775) );
OAI211xp5_ASAP7_75t_SL g1790 ( .A1(n_260), .A2(n_936), .B(n_1791), .C(n_1794), .Y(n_1790) );
AOI21xp5_ASAP7_75t_L g975 ( .A1(n_261), .A2(n_783), .B(n_799), .Y(n_975) );
INVx1_ASAP7_75t_L g1773 ( .A(n_262), .Y(n_1773) );
INVx1_ASAP7_75t_L g1166 ( .A(n_263), .Y(n_1166) );
INVx1_ASAP7_75t_L g1338 ( .A(n_267), .Y(n_1338) );
INVx1_ASAP7_75t_L g1087 ( .A(n_269), .Y(n_1087) );
INVx1_ASAP7_75t_L g921 ( .A(n_271), .Y(n_921) );
INVx1_ASAP7_75t_L g945 ( .A(n_272), .Y(n_945) );
INVx1_ASAP7_75t_L g1206 ( .A(n_274), .Y(n_1206) );
NAND2xp33_ASAP7_75t_SL g1031 ( .A(n_275), .B(n_1032), .Y(n_1031) );
NAND2xp5_ASAP7_75t_SL g1415 ( .A(n_279), .B(n_1050), .Y(n_1415) );
XNOR2x2_ASAP7_75t_L g915 ( .A(n_280), .B(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g1285 ( .A1(n_281), .A2(n_359), .B1(n_588), .B2(n_1030), .Y(n_1285) );
INVx1_ASAP7_75t_L g452 ( .A(n_282), .Y(n_452) );
INVx1_ASAP7_75t_L g459 ( .A(n_282), .Y(n_459) );
INVx1_ASAP7_75t_L g663 ( .A(n_283), .Y(n_663) );
INVx1_ASAP7_75t_L g1059 ( .A(n_287), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_288), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_290), .A2(n_321), .B1(n_784), .B2(n_1132), .C(n_1162), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_292), .A2(n_313), .B1(n_659), .B2(n_942), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g778 ( .A1(n_294), .A2(n_641), .B(n_779), .C(n_789), .Y(n_778) );
OAI21xp33_ASAP7_75t_L g1421 ( .A1(n_296), .A2(n_1294), .B(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1496 ( .A(n_297), .Y(n_1496) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_298), .Y(n_730) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_299), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_300), .Y(n_1073) );
AOI221xp5_ASAP7_75t_SL g1268 ( .A1(n_301), .A2(n_359), .B1(n_547), .B2(n_691), .C(n_831), .Y(n_1268) );
INVx1_ASAP7_75t_L g1197 ( .A(n_302), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_303), .B(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1550 ( .A(n_303), .Y(n_1550) );
INVx1_ASAP7_75t_L g749 ( .A(n_304), .Y(n_749) );
INVx1_ASAP7_75t_L g510 ( .A(n_305), .Y(n_510) );
OAI211xp5_ASAP7_75t_L g543 ( .A1(n_305), .A2(n_403), .B(n_544), .C(n_549), .Y(n_543) );
OAI211xp5_ASAP7_75t_SL g970 ( .A1(n_306), .A2(n_675), .B(n_971), .C(n_976), .Y(n_970) );
INVx1_ASAP7_75t_L g994 ( .A(n_306), .Y(n_994) );
INVx1_ASAP7_75t_L g836 ( .A(n_307), .Y(n_836) );
INVx1_ASAP7_75t_L g1291 ( .A(n_308), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1590 ( .A1(n_310), .A2(n_350), .B1(n_1548), .B2(n_1551), .Y(n_1590) );
INVx1_ASAP7_75t_L g397 ( .A(n_314), .Y(n_397) );
INVx1_ASAP7_75t_L g1799 ( .A(n_315), .Y(n_1799) );
INVx1_ASAP7_75t_L g835 ( .A(n_316), .Y(n_835) );
CKINVDCx16_ASAP7_75t_R g1349 ( .A(n_317), .Y(n_1349) );
AOI22xp5_ASAP7_75t_L g1509 ( .A1(n_323), .A2(n_354), .B1(n_660), .B2(n_1094), .Y(n_1509) );
INVx1_ASAP7_75t_L g705 ( .A(n_324), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_325), .B(n_954), .Y(n_953) );
OAI21xp33_ASAP7_75t_L g1461 ( .A1(n_326), .A2(n_632), .B(n_1462), .Y(n_1461) );
OAI21xp5_ASAP7_75t_SL g1096 ( .A1(n_329), .A2(n_838), .B(n_1097), .Y(n_1096) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_330), .A2(n_356), .B1(n_655), .B2(n_982), .C(n_984), .Y(n_981) );
INVx1_ASAP7_75t_L g425 ( .A(n_331), .Y(n_425) );
INVx1_ASAP7_75t_L g401 ( .A(n_332), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_333), .Y(n_914) );
INVxp67_ASAP7_75t_SL g1524 ( .A(n_334), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g1109 ( .A(n_335), .Y(n_1109) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_337), .Y(n_383) );
INVx1_ASAP7_75t_L g1246 ( .A(n_338), .Y(n_1246) );
INVx1_ASAP7_75t_L g989 ( .A(n_339), .Y(n_989) );
NOR2xp33_ASAP7_75t_R g1372 ( .A(n_340), .B(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1313 ( .A(n_341), .Y(n_1313) );
INVx1_ASAP7_75t_L g1147 ( .A(n_342), .Y(n_1147) );
OAI221xp5_ASAP7_75t_SL g1168 ( .A1(n_342), .A2(n_360), .B1(n_671), .B2(n_1169), .C(n_1171), .Y(n_1168) );
INVx1_ASAP7_75t_L g1250 ( .A(n_344), .Y(n_1250) );
OAI211xp5_ASAP7_75t_L g734 ( .A1(n_347), .A2(n_641), .B(n_735), .C(n_747), .Y(n_734) );
XOR2x2_ASAP7_75t_L g750 ( .A(n_348), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
INVx1_ASAP7_75t_L g434 ( .A(n_351), .Y(n_434) );
INVx1_ASAP7_75t_L g482 ( .A(n_351), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_353), .Y(n_630) );
OAI22xp33_ASAP7_75t_SL g1199 ( .A1(n_355), .A2(n_358), .B1(n_571), .B2(n_1045), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1208 ( .A1(n_355), .A2(n_358), .B1(n_671), .B2(n_1170), .C(n_1209), .Y(n_1208) );
XNOR2xp5_ASAP7_75t_L g1179 ( .A(n_357), .B(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1148 ( .A(n_360), .Y(n_1148) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_388), .B(n_1532), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx4f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_373), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g1807 ( .A(n_367), .B(n_376), .Y(n_1807) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g1816 ( .A(n_369), .B(n_372), .Y(n_1816) );
INVx1_ASAP7_75t_L g1819 ( .A(n_369), .Y(n_1819) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g1821 ( .A(n_372), .B(n_1819), .Y(n_1821) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g560 ( .A(n_376), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g435 ( .A(n_377), .B(n_387), .Y(n_435) );
AND2x4_ASAP7_75t_L g694 ( .A(n_377), .B(n_386), .Y(n_694) );
INVx1_ASAP7_75t_L g527 ( .A(n_378), .Y(n_527) );
AND2x4_ASAP7_75t_SL g1806 ( .A(n_378), .B(n_1807), .Y(n_1806) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x6_ASAP7_75t_L g379 ( .A(n_380), .B(n_385), .Y(n_379) );
OR2x6_ASAP7_75t_L g536 ( .A(n_380), .B(n_530), .Y(n_536) );
INVxp67_ASAP7_75t_L g954 ( .A(n_380), .Y(n_954) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
BUFx4f_ASAP7_75t_L g682 ( .A(n_381), .Y(n_682) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx2_ASAP7_75t_L g400 ( .A(n_383), .Y(n_400) );
NAND2x1_ASAP7_75t_L g405 ( .A(n_383), .B(n_384), .Y(n_405) );
INVx2_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
AND2x2_ASAP7_75t_L g532 ( .A(n_383), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g548 ( .A(n_383), .B(n_384), .Y(n_548) );
INVx1_ASAP7_75t_L g558 ( .A(n_383), .Y(n_558) );
OR2x2_ASAP7_75t_L g399 ( .A(n_384), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_384), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g533 ( .A(n_384), .Y(n_533) );
BUFx2_ASAP7_75t_L g552 ( .A(n_384), .Y(n_552) );
INVx1_ASAP7_75t_L g629 ( .A(n_384), .Y(n_629) );
AND2x2_ASAP7_75t_L g644 ( .A(n_384), .B(n_423), .Y(n_644) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g546 ( .A(n_386), .Y(n_546) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g542 ( .A(n_387), .Y(n_542) );
AND2x4_ASAP7_75t_L g556 ( .A(n_387), .B(n_557), .Y(n_556) );
XNOR2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_1100), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_864), .B1(n_1098), .B2(n_1099), .Y(n_389) );
INVx1_ASAP7_75t_L g1099 ( .A(n_390), .Y(n_1099) );
XNOR2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_697), .Y(n_390) );
OA22x2_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_563), .B1(n_564), .B2(n_696), .Y(n_391) );
INVx1_ASAP7_75t_L g696 ( .A(n_392), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_488), .C(n_525), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_439), .Y(n_394) );
OAI33xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_406), .A3(n_411), .B1(n_424), .B2(n_427), .B3(n_436), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_401), .B2(n_402), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_397), .A2(n_425), .B1(n_462), .B2(n_467), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_398), .A2(n_417), .B1(n_437), .B2(n_438), .Y(n_436) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g1380 ( .A(n_399), .Y(n_1380) );
BUFx2_ASAP7_75t_L g1479 ( .A(n_399), .Y(n_1479) );
BUFx3_ASAP7_75t_L g1518 ( .A(n_399), .Y(n_1518) );
AND2x2_ASAP7_75t_L g628 ( .A(n_400), .B(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g1276 ( .A(n_400), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_401), .A2(n_426), .B1(n_472), .B2(n_474), .Y(n_471) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_403), .A2(n_413), .B1(n_425), .B2(n_426), .Y(n_424) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx4f_ASAP7_75t_L g973 ( .A(n_404), .Y(n_973) );
INVx4_ASAP7_75t_L g1211 ( .A(n_404), .Y(n_1211) );
BUFx4f_ASAP7_75t_L g1281 ( .A(n_404), .Y(n_1281) );
OR2x6_ASAP7_75t_L g1383 ( .A(n_404), .B(n_1384), .Y(n_1383) );
BUFx4f_ASAP7_75t_L g1475 ( .A(n_404), .Y(n_1475) );
BUFx4f_ASAP7_75t_L g1507 ( .A(n_404), .Y(n_1507) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g1233 ( .A(n_405), .Y(n_1233) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_407), .B(n_1360), .Y(n_1359) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g812 ( .A(n_408), .Y(n_812) );
OR2x6_ASAP7_75t_L g861 ( .A(n_408), .B(n_862), .Y(n_861) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_408), .B(n_862), .Y(n_1077) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g586 ( .A(n_409), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_409), .B(n_627), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_416), .B2(n_417), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_412), .A2(n_437), .B1(n_447), .B2(n_453), .Y(n_446) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_415), .Y(n_793) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_415), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_416), .A2(n_438), .B1(n_485), .B2(n_487), .Y(n_484) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g685 ( .A(n_420), .Y(n_685) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_420), .Y(n_729) );
INVx2_ASAP7_75t_SL g979 ( .A(n_420), .Y(n_979) );
INVx1_ASAP7_75t_L g1061 ( .A(n_420), .Y(n_1061) );
INVx1_ASAP7_75t_L g1173 ( .A(n_420), .Y(n_1173) );
INVx2_ASAP7_75t_L g1525 ( .A(n_420), .Y(n_1525) );
INVx8_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g541 ( .A(n_421), .B(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_435), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g442 ( .A(n_432), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_432), .Y(n_524) );
OR2x2_ASAP7_75t_L g611 ( .A(n_432), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_SL g1377 ( .A(n_432), .B(n_435), .Y(n_1377) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g562 ( .A(n_433), .Y(n_562) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx4_ASAP7_75t_L g655 ( .A(n_435), .Y(n_655) );
INVx1_ASAP7_75t_SL g784 ( .A(n_435), .Y(n_784) );
INVx4_ASAP7_75t_L g831 ( .A(n_435), .Y(n_831) );
NAND4xp25_ASAP7_75t_L g1412 ( .A(n_435), .B(n_1413), .C(n_1414), .D(n_1415), .Y(n_1412) );
OAI33xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_446), .A3(n_461), .B1(n_471), .B2(n_476), .B3(n_484), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g1185 ( .A1(n_441), .A2(n_1186), .B1(n_1193), .B2(n_1194), .Y(n_1185) );
BUFx4f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx4f_ASAP7_75t_L g1024 ( .A(n_442), .Y(n_1024) );
BUFx8_ASAP7_75t_L g1239 ( .A(n_442), .Y(n_1239) );
BUFx2_ASAP7_75t_L g1426 ( .A(n_442), .Y(n_1426) );
NAND2xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_445), .Y(n_443) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_444), .Y(n_522) );
INVx1_ASAP7_75t_L g577 ( .A(n_444), .Y(n_577) );
AND3x4_ASAP7_75t_L g585 ( .A(n_444), .B(n_508), .C(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_444), .B(n_508), .Y(n_1335) );
INVx3_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
BUFx3_ASAP7_75t_L g508 ( .A(n_445), .Y(n_508) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g486 ( .A(n_448), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g1326 ( .A1(n_448), .A2(n_1327), .B1(n_1328), .B2(n_1329), .Y(n_1326) );
BUFx4f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x4_ASAP7_75t_L g492 ( .A(n_449), .B(n_493), .Y(n_492) );
OR2x4_ASAP7_75t_L g517 ( .A(n_449), .B(n_480), .Y(n_517) );
INVx2_ASAP7_75t_L g608 ( .A(n_449), .Y(n_608) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_450), .Y(n_460) );
INVx2_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_450), .B(n_459), .Y(n_470) );
AND2x4_ASAP7_75t_L g501 ( .A(n_450), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g591 ( .A(n_451), .Y(n_591) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
INVx2_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g635 ( .A(n_456), .B(n_611), .Y(n_635) );
INVx3_ASAP7_75t_L g1341 ( .A(n_456), .Y(n_1341) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g475 ( .A(n_457), .Y(n_475) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_457), .Y(n_1331) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
BUFx2_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
BUFx2_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
INVx2_ASAP7_75t_L g573 ( .A(n_460), .Y(n_573) );
AND2x4_ASAP7_75t_L g598 ( .A(n_460), .B(n_583), .Y(n_598) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_463), .Y(n_473) );
AND2x4_ASAP7_75t_L g519 ( .A(n_463), .B(n_493), .Y(n_519) );
INVx2_ASAP7_75t_L g856 ( .A(n_463), .Y(n_856) );
BUFx6f_ASAP7_75t_L g1079 ( .A(n_463), .Y(n_1079) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx8_ASAP7_75t_L g596 ( .A(n_464), .Y(n_596) );
INVx2_ASAP7_75t_L g713 ( .A(n_464), .Y(n_713) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_464), .Y(n_715) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AND2x4_ASAP7_75t_L g590 ( .A(n_466), .B(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g1336 ( .A1(n_467), .A2(n_1027), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g487 ( .A(n_468), .Y(n_487) );
CKINVDCx8_ASAP7_75t_R g1196 ( .A(n_468), .Y(n_1196) );
INVx3_ASAP7_75t_L g1328 ( .A(n_468), .Y(n_1328) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g624 ( .A(n_469), .Y(n_624) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g497 ( .A(n_470), .Y(n_497) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_477), .B(n_880), .C(n_881), .Y(n_879) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g600 ( .A(n_478), .Y(n_600) );
BUFx2_ASAP7_75t_L g716 ( .A(n_478), .Y(n_716) );
BUFx2_ASAP7_75t_L g1458 ( .A(n_478), .Y(n_1458) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g1034 ( .A(n_479), .Y(n_1034) );
NAND3x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .C(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g493 ( .A(n_480), .Y(n_493) );
OR2x6_ASAP7_75t_L g496 ( .A(n_480), .B(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g500 ( .A(n_480), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g576 ( .A(n_480), .B(n_577), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g862 ( .A(n_480), .B(n_483), .Y(n_862) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g575 ( .A(n_482), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_482), .B(n_645), .Y(n_1374) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g1427 ( .A1(n_487), .A2(n_1027), .B1(n_1428), .B2(n_1429), .C(n_1430), .Y(n_1427) );
OAI31xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_498), .A3(n_514), .B(n_520), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_497), .Y(n_1038) );
INVx1_ASAP7_75t_L g1190 ( .A(n_497), .Y(n_1190) );
CKINVDCx8_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
BUFx3_ASAP7_75t_L g592 ( .A(n_501), .Y(n_592) );
BUFx2_ASAP7_75t_L g619 ( .A(n_501), .Y(n_619) );
BUFx2_ASAP7_75t_L g709 ( .A(n_501), .Y(n_709) );
INVx2_ASAP7_75t_L g859 ( .A(n_501), .Y(n_859) );
BUFx2_ASAP7_75t_L g999 ( .A(n_501), .Y(n_999) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_501), .Y(n_1030) );
INVx1_ASAP7_75t_L g583 ( .A(n_502), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_510), .B2(n_511), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_504), .A2(n_550), .B1(n_553), .B2(n_554), .Y(n_549) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
AND2x4_ASAP7_75t_L g512 ( .A(n_507), .B(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI31xp33_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_534), .A3(n_543), .B(n_559), .Y(n_525) );
INVx3_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_532), .Y(n_653) );
INVx2_ASAP7_75t_L g692 ( .A(n_532), .Y(n_692) );
BUFx3_ASAP7_75t_L g823 ( .A(n_532), .Y(n_823) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g551 ( .A(n_542), .B(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_547), .Y(n_649) );
AND2x6_ASAP7_75t_L g661 ( .A(n_547), .B(n_627), .Y(n_661) );
AND2x4_ASAP7_75t_SL g674 ( .A(n_547), .B(n_645), .Y(n_674) );
BUFx3_ASAP7_75t_L g688 ( .A(n_547), .Y(n_688) );
INVx1_ASAP7_75t_L g782 ( .A(n_547), .Y(n_782) );
BUFx3_ASAP7_75t_L g830 ( .A(n_547), .Y(n_830) );
BUFx3_ASAP7_75t_L g984 ( .A(n_547), .Y(n_984) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_547), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g744 ( .A(n_548), .Y(n_744) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g677 ( .A(n_552), .Y(n_677) );
BUFx2_ASAP7_75t_L g816 ( .A(n_552), .Y(n_816) );
INVx1_ASAP7_75t_L g1371 ( .A(n_552), .Y(n_1371) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_557), .B(n_627), .Y(n_634) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g633 ( .A(n_562), .B(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_L g638 ( .A(n_562), .Y(n_638) );
INVx1_ASAP7_75t_L g1297 ( .A(n_562), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_562), .B(n_634), .Y(n_1364) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_620), .C(n_639), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_605), .C(n_616), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_584), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_578), .B2(n_579), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_570), .A2(n_579), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_570), .A2(n_579), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_570), .A2(n_579), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
AOI221x1_ASAP7_75t_L g1424 ( .A1(n_570), .A2(n_579), .B1(n_1403), .B2(n_1409), .C(n_1425), .Y(n_1424) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x4_ASAP7_75t_SL g848 ( .A(n_572), .B(n_574), .Y(n_848) );
AND2x2_ASAP7_75t_L g889 ( .A(n_572), .B(n_574), .Y(n_889) );
AND2x2_ASAP7_75t_L g995 ( .A(n_572), .B(n_574), .Y(n_995) );
AND2x6_ASAP7_75t_L g1353 ( .A(n_572), .B(n_576), .Y(n_1353) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g618 ( .A(n_574), .B(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_SL g849 ( .A(n_574), .B(n_580), .Y(n_849) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
OR2x2_ASAP7_75t_L g625 ( .A(n_575), .B(n_626), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_576), .B(n_590), .Y(n_637) );
INVx1_ASAP7_75t_L g1346 ( .A(n_576), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_576), .B(n_582), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_579), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_579), .A2(n_889), .B1(n_920), .B2(n_921), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_579), .A2(n_994), .B1(n_995), .B2(n_996), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_579), .A2(n_889), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
AO22x1_ASAP7_75t_L g1448 ( .A1(n_579), .A2(n_889), .B1(n_1449), .B2(n_1450), .Y(n_1448) );
AOI22xp5_ASAP7_75t_L g1771 ( .A1(n_579), .A2(n_995), .B1(n_1772), .B2(n_1773), .Y(n_1771) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI33xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .A3(n_593), .B1(n_599), .B2(n_600), .B3(n_601), .Y(n_584) );
AOI33xp33_ASAP7_75t_L g707 ( .A1(n_585), .A2(n_708), .A3(n_710), .B1(n_714), .B2(n_716), .B3(n_717), .Y(n_707) );
BUFx3_ASAP7_75t_L g765 ( .A(n_585), .Y(n_765) );
AOI33xp33_ASAP7_75t_L g850 ( .A1(n_585), .A2(n_851), .A3(n_852), .B1(n_854), .B2(n_857), .B3(n_860), .Y(n_850) );
AOI33xp33_ASAP7_75t_L g997 ( .A1(n_585), .A2(n_600), .A3(n_998), .B1(n_1000), .B2(n_1004), .B3(n_1007), .Y(n_997) );
INVx1_ASAP7_75t_L g1081 ( .A(n_585), .Y(n_1081) );
AOI33xp33_ASAP7_75t_L g1284 ( .A1(n_585), .A2(n_1285), .A3(n_1286), .B1(n_1287), .B2(n_1288), .B3(n_1289), .Y(n_1284) );
AOI33xp33_ASAP7_75t_L g1497 ( .A1(n_585), .A2(n_1498), .A3(n_1499), .B1(n_1500), .B2(n_1501), .B3(n_1502), .Y(n_1497) );
INVx2_ASAP7_75t_SL g695 ( .A(n_586), .Y(n_695) );
INVx1_ASAP7_75t_L g801 ( .A(n_586), .Y(n_801) );
OAI31xp33_ASAP7_75t_L g1320 ( .A1(n_586), .A2(n_1321), .A3(n_1325), .B(n_1347), .Y(n_1320) );
BUFx2_ASAP7_75t_L g1778 ( .A(n_588), .Y(n_1778) );
INVx8_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g762 ( .A(n_589), .Y(n_762) );
INVx2_ASAP7_75t_L g1041 ( .A(n_589), .Y(n_1041) );
INVx3_ASAP7_75t_L g1460 ( .A(n_589), .Y(n_1460) );
INVx8_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx3_ASAP7_75t_L g604 ( .A(n_590), .Y(n_604) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_590), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1344 ( .A(n_590), .Y(n_1344) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g614 ( .A(n_596), .B(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_596), .Y(n_770) );
INVx2_ASAP7_75t_SL g1115 ( .A(n_596), .Y(n_1115) );
INVx2_ASAP7_75t_SL g1241 ( .A(n_596), .Y(n_1241) );
INVx3_ASAP7_75t_L g1782 ( .A(n_596), .Y(n_1782) );
BUFx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g771 ( .A(n_598), .Y(n_771) );
BUFx12f_ASAP7_75t_L g853 ( .A(n_598), .Y(n_853) );
INVx5_ASAP7_75t_L g1003 ( .A(n_598), .Y(n_1003) );
AND2x4_ASAP7_75t_L g1395 ( .A(n_598), .B(n_1324), .Y(n_1395) );
AOI33xp33_ASAP7_75t_L g922 ( .A1(n_600), .A2(n_765), .A3(n_923), .B1(n_924), .B2(n_925), .B3(n_928), .Y(n_922) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx3_ASAP7_75t_L g776 ( .A(n_604), .Y(n_776) );
INVx2_ASAP7_75t_SL g877 ( .A(n_604), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_606), .B(n_1438), .Y(n_1437) );
OR2x6_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
OR2x2_ASAP7_75t_L g719 ( .A(n_607), .B(n_609), .Y(n_719) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g841 ( .A(n_610), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g615 ( .A(n_611), .Y(n_615) );
OR2x2_ASAP7_75t_L g623 ( .A(n_611), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g1324 ( .A(n_612), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1065 ( .A(n_613), .Y(n_1065) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_614), .A2(n_760), .B1(n_761), .B2(n_763), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_614), .A2(n_840), .B1(n_894), .B2(n_895), .Y(n_912) );
INVx2_ASAP7_75t_L g1010 ( .A(n_614), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_614), .A2(n_840), .B1(n_1127), .B2(n_1129), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_614), .A2(n_840), .B1(n_1206), .B2(n_1207), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_614), .A2(n_840), .B1(n_1226), .B2(n_1227), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_614), .A2(n_840), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
AND2x4_ASAP7_75t_L g761 ( .A(n_615), .B(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g840 ( .A(n_615), .B(n_762), .Y(n_840) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_616), .B(n_703), .C(n_718), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g1144 ( .A(n_616), .B(n_1145), .C(n_1154), .Y(n_1144) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND4xp75_ASAP7_75t_L g751 ( .A(n_617), .B(n_752), .C(n_755), .D(n_777), .Y(n_751) );
NAND3xp33_ASAP7_75t_SL g1071 ( .A(n_617), .B(n_1072), .C(n_1075), .Y(n_1071) );
NAND3xp33_ASAP7_75t_SL g1110 ( .A(n_617), .B(n_1111), .C(n_1121), .Y(n_1110) );
AND5x1_ASAP7_75t_L g1399 ( .A(n_617), .B(n_1400), .C(n_1424), .D(n_1435), .E(n_1439), .Y(n_1399) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g843 ( .A1(n_618), .A2(n_828), .B(n_844), .C(n_846), .Y(n_843) );
INVx3_ASAP7_75t_L g884 ( .A(n_618), .Y(n_884) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_618), .Y(n_930) );
NOR3xp33_ASAP7_75t_SL g1022 ( .A(n_618), .B(n_1023), .C(n_1043), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1237 ( .A(n_618), .B(n_1238), .C(n_1248), .Y(n_1237) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_618), .A2(n_848), .B1(n_849), .B2(n_1274), .C(n_1291), .Y(n_1290) );
BUFx2_ASAP7_75t_L g878 ( .A(n_619), .Y(n_878) );
AOI21xp33_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_630), .B(n_631), .Y(n_620) );
AOI21xp33_ASAP7_75t_SL g720 ( .A1(n_621), .A2(n_721), .B(n_722), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_621), .A2(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_621), .B(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_621), .B(n_914), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g931 ( .A1(n_621), .A2(n_932), .B(n_933), .Y(n_931) );
AOI21xp33_ASAP7_75t_SL g988 ( .A1(n_621), .A2(n_989), .B(n_990), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_621), .A2(n_844), .B1(n_1069), .B2(n_1070), .C(n_1071), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_621), .A2(n_844), .B1(n_1108), .B2(n_1109), .C(n_1110), .Y(n_1107) );
AOI21xp5_ASAP7_75t_L g1155 ( .A1(n_621), .A2(n_1156), .B(n_1157), .Y(n_1155) );
AOI21xp5_ASAP7_75t_L g1181 ( .A1(n_621), .A2(n_1182), .B(n_1183), .Y(n_1181) );
AOI21xp5_ASAP7_75t_L g1249 ( .A1(n_621), .A2(n_1250), .B(n_1251), .Y(n_1249) );
AOI211x1_ASAP7_75t_L g1444 ( .A1(n_621), .A2(n_1445), .B(n_1446), .C(n_1461), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_621), .B(n_1529), .Y(n_1528) );
AOI211x1_ASAP7_75t_L g1768 ( .A1(n_621), .A2(n_1769), .B(n_1770), .C(n_1784), .Y(n_1768) );
INVx8_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g1303 ( .A(n_623), .Y(n_1303) );
BUFx3_ASAP7_75t_L g1432 ( .A(n_624), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_625), .B(n_1394), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g678 ( .A(n_627), .Y(n_678) );
AND2x2_ASAP7_75t_L g815 ( .A(n_627), .B(n_816), .Y(n_815) );
INVx3_ASAP7_75t_L g658 ( .A(n_628), .Y(n_658) );
AND2x2_ASAP7_75t_L g666 ( .A(n_628), .B(n_645), .Y(n_666) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_628), .Y(n_906) );
INVx2_ASAP7_75t_L g1786 ( .A(n_632), .Y(n_1786) );
AND2x4_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
AND2x4_ASAP7_75t_L g838 ( .A(n_633), .B(n_635), .Y(n_838) );
INVx2_ASAP7_75t_L g1301 ( .A(n_635), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_636), .B(n_1388), .Y(n_1387) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OR2x6_ASAP7_75t_L g845 ( .A(n_637), .B(n_638), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_670), .B(n_695), .Y(n_639) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_SL g896 ( .A1(n_642), .A2(n_661), .B1(n_886), .B2(n_897), .C(n_899), .Y(n_896) );
INVx3_ASAP7_75t_L g936 ( .A(n_642), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_642), .A2(n_790), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_642), .A2(n_661), .B1(n_1108), .B2(n_1131), .C(n_1133), .Y(n_1130) );
NAND2xp5_ASAP7_75t_R g1471 ( .A(n_642), .B(n_1453), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_642), .B(n_1496), .Y(n_1513) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
BUFx2_ASAP7_75t_L g900 ( .A(n_643), .Y(n_900) );
INVx1_ASAP7_75t_L g1804 ( .A(n_643), .Y(n_1804) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx3_ASAP7_75t_L g660 ( .A(n_644), .Y(n_660) );
INVx2_ASAP7_75t_L g788 ( .A(n_644), .Y(n_788) );
BUFx3_ASAP7_75t_L g833 ( .A(n_644), .Y(n_833) );
AND2x4_ASAP7_75t_L g669 ( .A(n_645), .B(n_653), .Y(n_669) );
AND2x2_ASAP7_75t_L g826 ( .A(n_645), .B(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_L g1279 ( .A(n_645), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_645), .B(n_653), .Y(n_1298) );
AOI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_656), .B(n_661), .Y(n_646) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g1163 ( .A(n_649), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g940 ( .A(n_651), .Y(n_940) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g733 ( .A(n_652), .Y(n_733) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_653), .Y(n_746) );
INVx1_ASAP7_75t_L g1223 ( .A(n_653), .Y(n_1223) );
HB1xp67_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g737 ( .A(n_658), .Y(n_737) );
INVx2_ASAP7_75t_L g786 ( .A(n_658), .Y(n_786) );
INVx2_ASAP7_75t_L g942 ( .A(n_658), .Y(n_942) );
INVx1_ASAP7_75t_L g1094 ( .A(n_658), .Y(n_1094) );
INVx2_ASAP7_75t_L g1267 ( .A(n_658), .Y(n_1267) );
BUFx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g739 ( .A(n_660), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_661), .A2(n_736), .B(n_740), .Y(n_735) );
AOI21xp5_ASAP7_75t_SL g779 ( .A1(n_661), .A2(n_780), .B(n_785), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g825 ( .A1(n_661), .A2(n_826), .B1(n_828), .B2(n_829), .C(n_832), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g937 ( .A1(n_661), .A2(n_938), .B(n_941), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_661), .A2(n_668), .B(n_966), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_661), .A2(n_826), .B1(n_1021), .B2(n_1049), .C(n_1051), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1089 ( .A1(n_661), .A2(n_826), .B1(n_1069), .B2(n_1090), .C(n_1091), .Y(n_1089) );
AOI21xp5_ASAP7_75t_L g1160 ( .A1(n_661), .A2(n_1161), .B(n_1164), .Y(n_1160) );
AOI21xp5_ASAP7_75t_L g1202 ( .A1(n_661), .A2(n_1203), .B(n_1204), .Y(n_1202) );
AOI21xp5_ASAP7_75t_L g1220 ( .A1(n_661), .A2(n_1221), .B(n_1224), .Y(n_1220) );
AOI21xp5_ASAP7_75t_L g1468 ( .A1(n_661), .A2(n_1469), .B(n_1470), .Y(n_1468) );
INVx1_ASAP7_75t_L g1514 ( .A(n_661), .Y(n_1514) );
AOI21xp5_ASAP7_75t_L g1791 ( .A1(n_661), .A2(n_1792), .B(n_1793), .Y(n_1791) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_667), .B2(n_668), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_664), .A2(n_668), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_664), .A2(n_944), .B1(n_945), .B2(n_946), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_664), .A2(n_669), .B1(n_1463), .B2(n_1464), .Y(n_1467) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_666), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_666), .A2(n_669), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AND2x4_ASAP7_75t_L g1318 ( .A(n_666), .B(n_1297), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_668), .A2(n_1127), .B1(n_1128), .B2(n_1129), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_668), .A2(n_790), .B1(n_1795), .B2(n_1796), .Y(n_1794) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_669), .A2(n_760), .B1(n_763), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_669), .A2(n_790), .B1(n_835), .B2(n_836), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_669), .A2(n_790), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g947 ( .A(n_669), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1053 ( .A1(n_669), .A2(n_790), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
AOI22xp5_ASAP7_75t_L g1086 ( .A1(n_669), .A2(n_790), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_669), .A2(n_790), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
AOI22xp5_ASAP7_75t_L g1510 ( .A1(n_669), .A2(n_790), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g725 ( .A(n_672), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_672), .A2(n_676), .B1(n_920), .B2(n_921), .Y(n_955) );
INVx1_ASAP7_75t_L g1473 ( .A(n_672), .Y(n_1473) );
INVx4_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx3_ASAP7_75t_L g818 ( .A(n_674), .Y(n_818) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g1170 ( .A(n_676), .Y(n_1170) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g1278 ( .A(n_678), .Y(n_1278) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B1(n_684), .B2(n_686), .C(n_687), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_680), .A2(n_727), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g1171 ( .A1(n_680), .A2(n_1172), .B1(n_1173), .B2(n_1174), .C(n_1175), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_680), .A2(n_728), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx3_ASAP7_75t_L g1271 ( .A(n_682), .Y(n_1271) );
INVx4_ASAP7_75t_L g1406 ( .A(n_682), .Y(n_1406) );
OAI221xp5_ASAP7_75t_L g792 ( .A1(n_684), .A2(n_793), .B1(n_794), .B2(n_795), .C(n_796), .Y(n_792) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g783 ( .A(n_690), .Y(n_783) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_691), .Y(n_951) );
INVx1_ASAP7_75t_L g983 ( .A(n_691), .Y(n_983) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g798 ( .A(n_692), .Y(n_798) );
INVx1_ASAP7_75t_L g1520 ( .A(n_693), .Y(n_1520) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g799 ( .A(n_694), .Y(n_799) );
INVx2_ASAP7_75t_L g952 ( .A(n_694), .Y(n_952) );
INVx1_ASAP7_75t_L g1137 ( .A(n_694), .Y(n_1137) );
OAI221xp5_ASAP7_75t_L g1474 ( .A1(n_694), .A2(n_1475), .B1(n_1476), .B2(n_1477), .C(n_1480), .Y(n_1474) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_695), .A2(n_724), .B(n_734), .Y(n_723) );
AOI21xp5_ASAP7_75t_SL g891 ( .A1(n_695), .A2(n_892), .B(n_911), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_802), .B2(n_803), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
XNOR2x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_750), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_720), .C(n_723), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g768 ( .A(n_709), .Y(n_768) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx2_ASAP7_75t_L g774 ( .A(n_713), .Y(n_774) );
INVx3_ASAP7_75t_L g842 ( .A(n_713), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_713), .A2(n_1187), .B1(n_1188), .B2(n_1191), .C(n_1192), .Y(n_1186) );
OR2x6_ASAP7_75t_SL g1322 ( .A(n_713), .B(n_1323), .Y(n_1322) );
INVx5_ASAP7_75t_L g927 ( .A(n_715), .Y(n_927) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_715), .Y(n_1001) );
INVx2_ASAP7_75t_SL g1006 ( .A(n_715), .Y(n_1006) );
INVx2_ASAP7_75t_SL g1027 ( .A(n_715), .Y(n_1027) );
INVx3_ASAP7_75t_L g1333 ( .A(n_715), .Y(n_1333) );
AOI33xp33_ASAP7_75t_L g764 ( .A1(n_716), .A2(n_765), .A3(n_766), .B1(n_769), .B2(n_772), .B3(n_775), .Y(n_764) );
INVx5_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
BUFx2_ASAP7_75t_L g822 ( .A(n_744), .Y(n_822) );
BUFx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AND3x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .C(n_764), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_761), .A2(n_841), .B1(n_1087), .B2(n_1088), .Y(n_1097) );
AOI222xp33_ASAP7_75t_L g1300 ( .A1(n_761), .A2(n_1277), .B1(n_1301), .B2(n_1302), .C1(n_1303), .C2(n_1304), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_761), .A2(n_841), .B1(n_1511), .B2(n_1512), .Y(n_1527) );
AOI22xp5_ASAP7_75t_L g1348 ( .A1(n_762), .A2(n_858), .B1(n_1317), .B2(n_1349), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_765), .B(n_875), .Y(n_874) );
AOI33xp33_ASAP7_75t_L g1111 ( .A1(n_765), .A2(n_1112), .A3(n_1113), .B1(n_1117), .B2(n_1118), .B3(n_1120), .Y(n_1111) );
AOI33xp33_ASAP7_75t_L g1149 ( .A1(n_765), .A2(n_1118), .A3(n_1150), .B1(n_1151), .B2(n_1152), .B3(n_1153), .Y(n_1149) );
AOI33xp33_ASAP7_75t_L g1454 ( .A1(n_765), .A2(n_1455), .A3(n_1456), .B1(n_1457), .B2(n_1458), .B3(n_1459), .Y(n_1454) );
AOI33xp33_ASAP7_75t_L g1776 ( .A1(n_765), .A2(n_1034), .A3(n_1777), .B1(n_1779), .B2(n_1780), .B3(n_1783), .Y(n_1776) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_791), .B(n_800), .Y(n_777) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g797 ( .A(n_782), .Y(n_797) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g827 ( .A(n_788), .Y(n_827) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_790), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_793), .A2(n_977), .B1(n_978), .B2(n_980), .C(n_981), .Y(n_976) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx2_ASAP7_75t_L g958 ( .A(n_801), .Y(n_958) );
BUFx2_ASAP7_75t_L g1236 ( .A(n_801), .Y(n_1236) );
AOI21x1_ASAP7_75t_L g1260 ( .A1(n_801), .A2(n_1261), .B(n_1282), .Y(n_1260) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .C(n_843), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_813), .B(n_837), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g1046 ( .A1(n_810), .A2(n_1047), .B(n_1056), .Y(n_1046) );
OAI21xp33_ASAP7_75t_L g1789 ( .A1(n_810), .A2(n_1790), .B(n_1797), .Y(n_1789) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g1084 ( .A(n_811), .Y(n_1084) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_812), .B(n_1395), .Y(n_1394) );
NAND3xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_825), .C(n_834), .Y(n_813) );
AOI222xp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_817), .B1(n_818), .B2(n_819), .C1(n_820), .C2(n_824), .Y(n_814) );
INVx1_ASAP7_75t_L g910 ( .A(n_815), .Y(n_910) );
AOI222xp33_ASAP7_75t_L g1092 ( .A1(n_815), .A2(n_818), .B1(n_1073), .B2(n_1074), .C1(n_1093), .C2(n_1095), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g1273 ( .A1(n_816), .A2(n_1274), .B1(n_1275), .B2(n_1277), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_816), .A2(n_1275), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_817), .A2(n_819), .B1(n_848), .B2(n_849), .Y(n_847) );
INVx1_ASAP7_75t_L g909 ( .A(n_818), .Y(n_909) );
AOI222xp33_ASAP7_75t_L g1134 ( .A1(n_818), .A2(n_1122), .B1(n_1123), .B2(n_1135), .C1(n_1136), .C2(n_1138), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_818), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g898 ( .A(n_822), .Y(n_898) );
INVx1_ASAP7_75t_L g1176 ( .A(n_822), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_823), .Y(n_1132) );
INVx2_ASAP7_75t_L g1262 ( .A(n_826), .Y(n_1262) );
AND2x4_ASAP7_75t_L g1389 ( .A(n_827), .B(n_1390), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_835), .A2(n_836), .B1(n_840), .B2(n_841), .Y(n_839) );
INVx1_ASAP7_75t_SL g1020 ( .A(n_838), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g1064 ( .A1(n_840), .A2(n_1054), .B1(n_1055), .B2(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_841), .Y(n_1294) );
INVx2_ASAP7_75t_L g1036 ( .A(n_842), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_844), .B(n_886), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_844), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1018) );
INVx3_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx5_ASAP7_75t_L g1441 ( .A(n_845), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_850), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g1072 ( .A1(n_848), .A2(n_849), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
AOI22xp5_ASAP7_75t_L g1492 ( .A1(n_848), .A2(n_849), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
INVx1_ASAP7_75t_L g1045 ( .A(n_849), .Y(n_1045) );
BUFx2_ASAP7_75t_L g882 ( .A(n_853), .Y(n_882) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_856), .A2(n_1195), .B1(n_1196), .B2(n_1197), .C(n_1198), .Y(n_1194) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g1008 ( .A(n_859), .Y(n_1008) );
INVx2_ASAP7_75t_L g1042 ( .A(n_859), .Y(n_1042) );
INVx1_ASAP7_75t_SL g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1289 ( .A(n_861), .Y(n_1289) );
INVx1_ASAP7_75t_L g1502 ( .A(n_861), .Y(n_1502) );
INVx1_ASAP7_75t_L g1098 ( .A(n_864), .Y(n_1098) );
XOR2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_960), .Y(n_864) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
OAI22x1_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B1(n_915), .B2(n_959), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
XNOR2x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
AND3x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_891), .C(n_913), .Y(n_870) );
NOR2xp33_ASAP7_75t_SL g871 ( .A(n_872), .B(n_883), .Y(n_871) );
OAI21xp5_ASAP7_75t_SL g872 ( .A1(n_873), .A2(n_874), .B(n_879), .Y(n_872) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .C(n_887), .Y(n_883) );
INVx1_ASAP7_75t_L g1011 ( .A(n_884), .Y(n_1011) );
NAND2xp5_ASAP7_75t_SL g1451 ( .A(n_884), .B(n_1452), .Y(n_1451) );
AND4x1_ASAP7_75t_L g1491 ( .A(n_884), .B(n_1492), .C(n_1495), .D(n_1497), .Y(n_1491) );
NAND4xp25_ASAP7_75t_SL g1770 ( .A(n_884), .B(n_1771), .C(n_1774), .D(n_1776), .Y(n_1770) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .C(n_901), .Y(n_892) );
AOI31xp33_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .A3(n_907), .B(n_908), .Y(n_901) );
INVx2_ASAP7_75t_SL g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g1052 ( .A(n_905), .Y(n_1052) );
INVx3_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
BUFx6f_ASAP7_75t_L g1802 ( .A(n_906), .Y(n_1802) );
INVx1_ASAP7_75t_L g1138 ( .A(n_910), .Y(n_1138) );
INVx1_ASAP7_75t_L g959 ( .A(n_915), .Y(n_959) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_931), .C(n_934), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_929), .C(n_930), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_922), .Y(n_918) );
INVx8_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g1431 ( .A1(n_927), .A2(n_1417), .B1(n_1432), .B2(n_1433), .C(n_1434), .Y(n_1431) );
NOR3xp33_ASAP7_75t_L g1184 ( .A(n_930), .B(n_1185), .C(n_1199), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_948), .B(n_956), .Y(n_934) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_946), .A2(n_1128), .B1(n_1166), .B2(n_1167), .Y(n_1165) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_950), .B(n_953), .Y(n_949) );
INVx1_ASAP7_75t_L g1523 ( .A(n_954), .Y(n_1523) );
OAI21xp5_ASAP7_75t_L g1158 ( .A1(n_956), .A2(n_1159), .B(n_1168), .Y(n_1158) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g987 ( .A(n_958), .Y(n_987) );
HB1xp67_ASAP7_75t_L g1420 ( .A(n_958), .Y(n_1420) );
XNOR2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_1012), .Y(n_960) );
NAND3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_988), .C(n_991), .Y(n_962) );
OAI31xp33_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_970), .A3(n_985), .B(n_986), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_967), .Y(n_964) );
OAI211xp5_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B(n_974), .C(n_975), .Y(n_971) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
NOR3xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_1009), .C(n_1011), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_997), .Y(n_992) );
INVx1_ASAP7_75t_L g1044 ( .A(n_995), .Y(n_1044) );
INVx2_ASAP7_75t_R g1002 ( .A(n_1003), .Y(n_1002) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1003), .Y(n_1032) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1003), .Y(n_1116) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
XNOR2x1_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1066), .Y(n_1014) );
NAND4xp75_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1022), .C(n_1046), .D(n_1064), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1025), .B1(n_1033), .B2(n_1035), .Y(n_1023) );
OAI211xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .B(n_1028), .C(n_1031), .Y(n_1025) );
OAI22xp5_ASAP7_75t_SL g1425 ( .A1(n_1033), .A2(n_1426), .B1(n_1427), .B2(n_1431), .Y(n_1425) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g1119 ( .A(n_1034), .Y(n_1119) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1034), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1037), .B1(n_1038), .B2(n_1039), .C(n_1040), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1053), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1059), .B1(n_1060), .B2(n_1062), .C(n_1063), .Y(n_1057) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1083), .Y(n_1067) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1078), .B1(n_1080), .B2(n_1082), .Y(n_1075) );
AOI21xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1085), .B(n_1096), .Y(n_1083) );
AOI21xp5_ASAP7_75t_L g1124 ( .A1(n_1084), .A2(n_1125), .B(n_1139), .Y(n_1124) );
OAI21xp5_ASAP7_75t_L g1200 ( .A1(n_1084), .A2(n_1201), .B(n_1208), .Y(n_1200) );
OAI21xp5_ASAP7_75t_L g1465 ( .A1(n_1084), .A2(n_1466), .B(n_1472), .Y(n_1465) );
NAND3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1089), .C(n_1092), .Y(n_1085) );
AO22x2_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B1(n_1488), .B2(n_1531), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
AO22x2_ASAP7_75t_L g1102 ( .A1(n_1103), .A2(n_1254), .B1(n_1255), .B2(n_1487), .Y(n_1102) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1103), .Y(n_1487) );
XNOR2xp5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1177), .Y(n_1103) );
XOR2xp5_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1142), .Y(n_1104) );
XNOR2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1141), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1124), .Y(n_1106) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
OAI22xp5_ASAP7_75t_SL g1238 ( .A1(n_1119), .A2(n_1239), .B1(n_1240), .B2(n_1245), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1130), .C(n_1134), .Y(n_1125) );
NAND3xp33_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1155), .C(n_1158), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1149), .Y(n_1145) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
BUFx3_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
AO22x2_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1215), .B1(n_1216), .B2(n_1253), .Y(n_1178) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1179), .Y(n_1253) );
AND4x1_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1184), .C(n_1200), .D(n_1214), .Y(n_1180) );
OAI221xp5_ASAP7_75t_L g1240 ( .A1(n_1188), .A2(n_1241), .B1(n_1242), .B2(n_1243), .C(n_1244), .Y(n_1240) );
INVx3_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
OAI211xp5_ASAP7_75t_L g1209 ( .A1(n_1195), .A2(n_1210), .B(n_1212), .C(n_1213), .Y(n_1209) );
OAI221xp5_ASAP7_75t_L g1245 ( .A1(n_1196), .A2(n_1230), .B1(n_1241), .B2(n_1246), .C(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1211), .Y(n_1272) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1211), .Y(n_1407) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
AND4x1_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1237), .C(n_1249), .D(n_1252), .Y(n_1217) );
OAI21xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1228), .B(n_1236), .Y(n_1218) );
INVx2_ASAP7_75t_SL g1222 ( .A(n_1223), .Y(n_1222) );
OAI211xp5_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1231), .B(n_1234), .C(n_1235), .Y(n_1229) );
OAI211xp5_ASAP7_75t_L g1416 ( .A1(n_1231), .A2(n_1417), .B(n_1418), .C(n_1419), .Y(n_1416) );
OAI211xp5_ASAP7_75t_L g1798 ( .A1(n_1231), .A2(n_1799), .B(n_1800), .C(n_1801), .Y(n_1798) );
INVx5_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx2_ASAP7_75t_SL g1232 ( .A(n_1233), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1373 ( .A(n_1233), .B(n_1374), .Y(n_1373) );
O2A1O1Ixp5_ASAP7_75t_SL g1503 ( .A1(n_1236), .A2(n_1504), .B(n_1515), .C(n_1526), .Y(n_1503) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
AO22x2_ASAP7_75t_L g1255 ( .A1(n_1256), .A2(n_1442), .B1(n_1485), .B2(n_1486), .Y(n_1255) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1256), .Y(n_1485) );
XNOR2xp5_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1398), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1258), .A2(n_1312), .B1(n_1396), .B2(n_1397), .Y(n_1257) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1258), .Y(n_1397) );
NAND3xp33_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1305), .C(n_1309), .Y(n_1258) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1260), .Y(n_1306) );
AOI22xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B1(n_1266), .B2(n_1268), .Y(n_1263) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_1270), .A2(n_1278), .B1(n_1279), .B2(n_1280), .Y(n_1269) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AOI22xp5_ASAP7_75t_L g1404 ( .A1(n_1278), .A2(n_1279), .B1(n_1405), .B2(n_1411), .Y(n_1404) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1283), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1290), .Y(n_1283) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1292), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1299), .Y(n_1292) );
NAND2x1_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1295), .Y(n_1293) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_1296), .A2(n_1317), .B1(n_1318), .B2(n_1319), .Y(n_1316) );
AND2x4_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1300), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1422 ( .A1(n_1301), .A2(n_1303), .B1(n_1410), .B2(n_1423), .Y(n_1422) );
OAI21xp5_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B(n_1308), .Y(n_1305) );
OAI21xp33_ASAP7_75t_L g1309 ( .A1(n_1308), .A2(n_1310), .B(n_1311), .Y(n_1309) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1312), .Y(n_1396) );
XNOR2xp5_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1314), .Y(n_1312) );
NOR2x1_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1356), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1320), .Y(n_1315) );
INVx3_ASAP7_75t_L g1438 ( .A(n_1318), .Y(n_1438) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
HB1xp67_ASAP7_75t_L g1351 ( .A(n_1324), .Y(n_1351) );
OAI221xp5_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1330), .B1(n_1336), .B2(n_1339), .C(n_1345), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1332), .B1(n_1333), .B2(n_1334), .C(n_1335), .Y(n_1330) );
OR2x6_ASAP7_75t_L g1345 ( .A(n_1331), .B(n_1346), .Y(n_1345) );
OAI211xp5_ASAP7_75t_L g1378 ( .A1(n_1332), .A2(n_1379), .B(n_1381), .C(n_1382), .Y(n_1378) );
OAI21xp5_ASAP7_75t_SL g1339 ( .A1(n_1340), .A2(n_1342), .B(n_1343), .Y(n_1339) );
INVx3_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
AOI22xp5_ASAP7_75t_L g1362 ( .A1(n_1349), .A2(n_1363), .B1(n_1365), .B2(n_1366), .Y(n_1362) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx4_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
NAND3xp33_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1385), .C(n_1391), .Y(n_1356) );
NOR3xp33_ASAP7_75t_SL g1357 ( .A(n_1358), .B(n_1372), .C(n_1375), .Y(n_1357) );
OAI21xp5_ASAP7_75t_SL g1358 ( .A1(n_1359), .A2(n_1361), .B(n_1362), .Y(n_1358) );
INVx1_ASAP7_75t_SL g1363 ( .A(n_1364), .Y(n_1363) );
INVx2_ASAP7_75t_SL g1366 ( .A(n_1367), .Y(n_1366) );
NAND2x2_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1370), .Y(n_1367) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1368), .Y(n_1384) );
INVx2_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx2_ASAP7_75t_SL g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1374), .Y(n_1390) );
OAI21xp5_ASAP7_75t_L g1375 ( .A1(n_1376), .A2(n_1378), .B(n_1383), .Y(n_1375) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1387), .Y(n_1385) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1393), .Y(n_1391) );
AOI21xp5_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1420), .B(n_1421), .Y(n_1400) );
NAND4xp25_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1404), .C(n_1412), .D(n_1416), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g1516 ( .A1(n_1407), .A2(n_1517), .B1(n_1518), .B2(n_1519), .C(n_1520), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1437), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1441), .B(n_1453), .Y(n_1452) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1441), .B(n_1496), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1441), .B(n_1775), .Y(n_1774) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1442), .Y(n_1486) );
XOR2x2_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1484), .Y(n_1442) );
NAND2xp5_ASAP7_75t_SL g1443 ( .A(n_1444), .B(n_1465), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1454), .Y(n_1446) );
NOR2xp33_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1451), .Y(n_1447) );
NAND3xp33_ASAP7_75t_SL g1466 ( .A(n_1467), .B(n_1468), .C(n_1471), .Y(n_1466) );
INVx2_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx4_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1488), .Y(n_1531) );
HB1xp67_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
XOR2xp5_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1530), .Y(n_1489) );
NAND3xp33_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1503), .C(n_1528), .Y(n_1490) );
NAND4xp25_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1510), .C(n_1513), .D(n_1514), .Y(n_1504) );
OAI211xp5_ASAP7_75t_L g1505 ( .A1(n_1506), .A2(n_1507), .B(n_1508), .C(n_1509), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_1522), .A2(n_1523), .B1(n_1524), .B2(n_1525), .Y(n_1521) );
OAI221xp5_ASAP7_75t_SL g1532 ( .A1(n_1533), .A2(n_1762), .B1(n_1765), .B2(n_1805), .C(n_1808), .Y(n_1532) );
AOI21xp5_ASAP7_75t_L g1533 ( .A1(n_1534), .A2(n_1676), .B(n_1729), .Y(n_1533) );
NAND4xp25_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1646), .C(n_1662), .D(n_1668), .Y(n_1534) );
NOR5xp2_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1600), .C(n_1613), .D(n_1620), .E(n_1643), .Y(n_1535) );
OAI21xp5_ASAP7_75t_SL g1536 ( .A1(n_1537), .A2(n_1557), .B(n_1576), .Y(n_1536) );
NOR2xp33_ASAP7_75t_L g1577 ( .A(n_1537), .B(n_1558), .Y(n_1577) );
OAI31xp33_ASAP7_75t_L g1754 ( .A1(n_1537), .A2(n_1755), .A3(n_1756), .B(n_1757), .Y(n_1754) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1538), .B(n_1633), .Y(n_1675) );
AOI221xp5_ASAP7_75t_L g1692 ( .A1(n_1538), .A2(n_1616), .B1(n_1693), .B2(n_1694), .C(n_1696), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1553), .Y(n_1538) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1539), .Y(n_1603) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1539), .Y(n_1615) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1539), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1539), .B(n_1591), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1547), .Y(n_1539) );
INVx2_ASAP7_75t_L g1764 ( .A(n_1541), .Y(n_1764) );
AND2x6_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1543), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1542), .B(n_1546), .Y(n_1545) );
AND2x4_ASAP7_75t_L g1548 ( .A(n_1542), .B(n_1549), .Y(n_1548) );
AND2x6_ASAP7_75t_L g1551 ( .A(n_1542), .B(n_1552), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1542), .B(n_1546), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1542), .B(n_1546), .Y(n_1637) );
OAI21xp5_ASAP7_75t_L g1818 ( .A1(n_1543), .A2(n_1819), .B(n_1820), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1544), .B(n_1550), .Y(n_1549) );
CKINVDCx5p33_ASAP7_75t_R g1591 ( .A(n_1553), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1612 ( .A(n_1553), .B(n_1588), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1553), .B(n_1603), .Y(n_1640) );
HB1xp67_ASAP7_75t_SL g1658 ( .A(n_1553), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1553), .B(n_1633), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1553), .B(n_1560), .Y(n_1734) );
AND2x4_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1556), .Y(n_1553) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1557), .Y(n_1745) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1563), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1558), .B(n_1595), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1752 ( .A(n_1558), .B(n_1641), .Y(n_1752) );
CKINVDCx14_ASAP7_75t_R g1558 ( .A(n_1559), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1559), .B(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1559), .B(n_1588), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1626 ( .A(n_1559), .B(n_1580), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1559), .B(n_1608), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1559), .B(n_1687), .Y(n_1686) );
NOR2xp33_ASAP7_75t_L g1698 ( .A(n_1559), .B(n_1612), .Y(n_1698) );
NOR2xp33_ASAP7_75t_L g1718 ( .A(n_1559), .B(n_1654), .Y(n_1718) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_1559), .B(n_1621), .Y(n_1728) );
INVx3_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
CKINVDCx5p33_ASAP7_75t_R g1592 ( .A(n_1560), .Y(n_1592) );
NOR2xp33_ASAP7_75t_L g1629 ( .A(n_1560), .B(n_1597), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1560), .B(n_1565), .Y(n_1632) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_1560), .B(n_1581), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1560), .B(n_1674), .Y(n_1702) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1560), .B(n_1683), .Y(n_1724) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1560), .B(n_1608), .Y(n_1726) );
NAND2xp5_ASAP7_75t_L g1756 ( .A(n_1560), .B(n_1654), .Y(n_1756) );
AND2x4_ASAP7_75t_SL g1560 ( .A(n_1561), .B(n_1562), .Y(n_1560) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
OR2x2_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1568), .Y(n_1564) );
INVx2_ASAP7_75t_L g1580 ( .A(n_1565), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1565), .B(n_1573), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1565), .B(n_1582), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1657 ( .A(n_1565), .B(n_1581), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1565), .B(n_1681), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1565), .B(n_1570), .Y(n_1695) );
OAI322xp33_ASAP7_75t_L g1696 ( .A1(n_1565), .A2(n_1579), .A3(n_1674), .B1(n_1697), .B2(n_1699), .C1(n_1703), .C2(n_1705), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1732 ( .A(n_1565), .B(n_1667), .Y(n_1732) );
OR2x2_ASAP7_75t_L g1743 ( .A(n_1565), .B(n_1570), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1566), .B(n_1567), .Y(n_1565) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1568), .B(n_1580), .Y(n_1642) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1568), .Y(n_1683) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1573), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1569), .B(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
OR2x2_ASAP7_75t_L g1597 ( .A(n_1570), .B(n_1598), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1570), .B(n_1573), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1570), .B(n_1580), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1572), .Y(n_1570) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1573), .Y(n_1582) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1573), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1573), .B(n_1580), .Y(n_1715) );
NAND2x1_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1575), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_1577), .A2(n_1578), .B1(n_1584), .B2(n_1593), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1583), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1581), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1580), .B(n_1596), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1580), .B(n_1608), .Y(n_1607) );
OR2x2_ASAP7_75t_L g1652 ( .A(n_1580), .B(n_1653), .Y(n_1652) );
OR2x2_ASAP7_75t_L g1688 ( .A(n_1580), .B(n_1597), .Y(n_1688) );
NOR2xp33_ASAP7_75t_L g1700 ( .A(n_1580), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1581), .B(n_1625), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1631 ( .A(n_1581), .B(n_1632), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1581), .B(n_1592), .Y(n_1681) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1583), .Y(n_1645) );
OAI21xp5_ASAP7_75t_L g1733 ( .A1(n_1583), .A2(n_1734), .B(n_1735), .Y(n_1733) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1592), .Y(n_1585) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1586), .Y(n_1761) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1601 ( .A(n_1587), .B(n_1602), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1591), .Y(n_1587) );
INVx2_ASAP7_75t_SL g1622 ( .A(n_1588), .Y(n_1622) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1588), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1590), .Y(n_1588) );
OR2x2_ASAP7_75t_L g1621 ( .A(n_1591), .B(n_1622), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1591), .B(n_1615), .Y(n_1628) );
NOR2xp33_ASAP7_75t_L g1647 ( .A(n_1591), .B(n_1648), .Y(n_1647) );
OAI22xp5_ASAP7_75t_L g1678 ( .A1(n_1591), .A2(n_1658), .B1(n_1679), .B2(n_1682), .Y(n_1678) );
NAND3xp33_ASAP7_75t_L g1717 ( .A(n_1591), .B(n_1608), .C(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1592), .Y(n_1606) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1592), .B(n_1714), .Y(n_1713) );
INVxp33_ASAP7_75t_SL g1593 ( .A(n_1594), .Y(n_1593) );
NOR2xp33_ASAP7_75t_SL g1594 ( .A(n_1595), .B(n_1599), .Y(n_1594) );
INVx2_ASAP7_75t_L g1619 ( .A(n_1595), .Y(n_1619) );
AOI222xp33_ASAP7_75t_L g1668 ( .A1(n_1596), .A2(n_1669), .B1(n_1670), .B2(n_1671), .C1(n_1673), .C2(n_1675), .Y(n_1668) );
NOR2xp33_ASAP7_75t_L g1704 ( .A(n_1596), .B(n_1683), .Y(n_1704) );
A2O1A1Ixp33_ASAP7_75t_L g1757 ( .A1(n_1596), .A2(n_1606), .B(n_1675), .C(n_1687), .Y(n_1757) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
A2O1A1Ixp33_ASAP7_75t_L g1758 ( .A1(n_1599), .A2(n_1670), .B(n_1698), .C(n_1759), .Y(n_1758) );
OAI21xp5_ASAP7_75t_SL g1600 ( .A1(n_1601), .A2(n_1604), .B(n_1609), .Y(n_1600) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1601), .Y(n_1753) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1603), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1603), .B(n_1650), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1603), .B(n_1611), .Y(n_1693) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1603), .B(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1607), .Y(n_1605) );
AOI221xp5_ASAP7_75t_L g1744 ( .A1(n_1607), .A2(n_1710), .B1(n_1745), .B2(n_1746), .C(n_1747), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1608), .B(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1608), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1608), .B(n_1632), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1610), .B(n_1645), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1659 ( .A(n_1610), .B(n_1660), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1711 ( .A(n_1611), .B(n_1670), .Y(n_1711) );
INVx2_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
AOI21xp33_ASAP7_75t_L g1677 ( .A1(n_1612), .A2(n_1678), .B(n_1684), .Y(n_1677) );
INVxp67_ASAP7_75t_SL g1613 ( .A(n_1614), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1619), .Y(n_1616) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
OAI21xp33_ASAP7_75t_L g1639 ( .A1(n_1618), .A2(n_1640), .B(n_1641), .Y(n_1639) );
OAI211xp5_ASAP7_75t_SL g1620 ( .A1(n_1621), .A2(n_1623), .B(n_1627), .C(n_1639), .Y(n_1620) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1621), .Y(n_1746) );
INVx2_ASAP7_75t_L g1654 ( .A(n_1622), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1622), .B(n_1737), .Y(n_1736) );
O2A1O1Ixp33_ASAP7_75t_SL g1747 ( .A1(n_1622), .A2(n_1689), .B(n_1748), .C(n_1749), .Y(n_1747) );
CKINVDCx14_ASAP7_75t_R g1623 ( .A(n_1624), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1625), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
OR2x2_ASAP7_75t_L g1689 ( .A(n_1626), .B(n_1653), .Y(n_1689) );
AOI211xp5_ASAP7_75t_L g1738 ( .A1(n_1626), .A2(n_1739), .B(n_1740), .C(n_1742), .Y(n_1738) );
AOI221xp5_ASAP7_75t_L g1627 ( .A1(n_1628), .A2(n_1629), .B1(n_1630), .B2(n_1633), .C(n_1634), .Y(n_1627) );
NOR2xp33_ASAP7_75t_L g1651 ( .A(n_1628), .B(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1628), .Y(n_1705) );
O2A1O1Ixp33_ASAP7_75t_L g1750 ( .A1(n_1629), .A2(n_1751), .B(n_1753), .C(n_1754), .Y(n_1750) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1649 ( .A(n_1631), .B(n_1650), .Y(n_1649) );
INVx2_ASAP7_75t_L g1650 ( .A(n_1633), .Y(n_1650) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1634), .B(n_1717), .Y(n_1716) );
INVx3_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1636), .B(n_1638), .Y(n_1635) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1640), .Y(n_1749) );
INVx2_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVxp67_ASAP7_75t_SL g1643 ( .A(n_1644), .Y(n_1643) );
O2A1O1Ixp33_ASAP7_75t_L g1646 ( .A1(n_1647), .A2(n_1651), .B(n_1654), .C(n_1655), .Y(n_1646) );
OAI31xp33_ASAP7_75t_L g1662 ( .A1(n_1647), .A2(n_1651), .A3(n_1663), .B(n_1666), .Y(n_1662) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1650), .B(n_1674), .Y(n_1673) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1650), .B(n_1674), .Y(n_1709) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1652), .Y(n_1707) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1654), .B(n_1665), .Y(n_1664) );
O2A1O1Ixp33_ASAP7_75t_L g1655 ( .A1(n_1656), .A2(n_1658), .B(n_1659), .C(n_1661), .Y(n_1655) );
AOI21xp33_ASAP7_75t_L g1759 ( .A1(n_1656), .A2(n_1760), .B(n_1761), .Y(n_1759) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
NAND2xp5_ASAP7_75t_L g1727 ( .A(n_1660), .B(n_1728), .Y(n_1727) );
CKINVDCx14_ASAP7_75t_R g1755 ( .A(n_1660), .Y(n_1755) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1661), .Y(n_1670) );
AOI221xp5_ASAP7_75t_L g1730 ( .A1(n_1661), .A2(n_1693), .B1(n_1731), .B2(n_1733), .C(n_1738), .Y(n_1730) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1666), .Y(n_1748) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1669), .Y(n_1760) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
AOI222xp33_ASAP7_75t_L g1719 ( .A1(n_1673), .A2(n_1708), .B1(n_1720), .B2(n_1721), .C1(n_1723), .C2(n_1725), .Y(n_1719) );
NAND5xp2_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1692), .C(n_1706), .D(n_1719), .E(n_1727), .Y(n_1676) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVxp67_ASAP7_75t_SL g1739 ( .A(n_1681), .Y(n_1739) );
AOI21xp33_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1689), .B(n_1690), .Y(n_1684) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1689), .Y(n_1720) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVxp67_ASAP7_75t_SL g1697 ( .A(n_1698), .Y(n_1697) );
INVxp67_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
HB1xp67_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
AOI221xp5_ASAP7_75t_L g1706 ( .A1(n_1707), .A2(n_1708), .B1(n_1710), .B2(n_1712), .C(n_1716), .Y(n_1706) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1722), .Y(n_1741) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
INVxp67_ASAP7_75t_SL g1725 ( .A(n_1726), .Y(n_1725) );
NAND4xp25_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1744), .C(n_1750), .D(n_1758), .Y(n_1729) );
INVxp67_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
CKINVDCx20_ASAP7_75t_R g1762 ( .A(n_1763), .Y(n_1762) );
CKINVDCx20_ASAP7_75t_R g1763 ( .A(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
XNOR2x2_ASAP7_75t_L g1766 ( .A(n_1767), .B(n_1768), .Y(n_1766) );
HB1xp67_ASAP7_75t_L g1811 ( .A(n_1768), .Y(n_1811) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1785), .B(n_1789), .Y(n_1784) );
AOI21xp5_ASAP7_75t_L g1785 ( .A1(n_1786), .A2(n_1787), .B(n_1788), .Y(n_1785) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
CKINVDCx5p33_ASAP7_75t_R g1805 ( .A(n_1806), .Y(n_1805) );
INVxp33_ASAP7_75t_SL g1809 ( .A(n_1810), .Y(n_1809) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
HB1xp67_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
BUFx3_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
HB1xp67_ASAP7_75t_L g1817 ( .A(n_1818), .Y(n_1817) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
endmodule