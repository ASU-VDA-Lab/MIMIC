module fake_jpeg_5336_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

AOI21xp33_ASAP7_75t_L g10 ( 
.A1(n_4),
.A2(n_5),
.B(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_18),
.B1(n_9),
.B2(n_12),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_0),
.CON(n_15),
.SN(n_15)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_21),
.B(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_20),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_25),
.B(n_27),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_12),
.B1(n_9),
.B2(n_8),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_8),
.B1(n_11),
.B2(n_6),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_21),
.C(n_14),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_26),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_24),
.C(n_23),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_37),
.B1(n_36),
.B2(n_16),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_45)
);

OAI21x1_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_42),
.B(n_11),
.Y(n_46)
);


endmodule