module fake_jpeg_26857_n_249 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_7),
.B(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_41),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_24),
.B1(n_27),
.B2(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_52),
.B1(n_57),
.B2(n_22),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_24),
.B1(n_27),
.B2(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_62),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_22),
.B1(n_20),
.B2(n_26),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_38),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_69),
.B(n_72),
.C(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_71),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_18),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_20),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_35),
.B1(n_22),
.B2(n_42),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_90),
.B1(n_94),
.B2(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_86),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_18),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_25),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_21),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_35),
.B1(n_17),
.B2(n_29),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_23),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_74),
.B(n_30),
.Y(n_140)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_104),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_51),
.B(n_60),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_115),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_64),
.C(n_36),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_51),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_118),
.B1(n_88),
.B2(n_73),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_17),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_76),
.Y(n_127)
);

OAI22x1_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_84),
.B1(n_85),
.B2(n_53),
.Y(n_139)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_41),
.C(n_40),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_40),
.B(n_53),
.C(n_17),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_69),
.A2(n_30),
.B1(n_29),
.B2(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_130),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_139),
.B1(n_105),
.B2(n_113),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_69),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_100),
.B(n_97),
.Y(n_160)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_76),
.B1(n_72),
.B2(n_90),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_30),
.B1(n_32),
.B2(n_3),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_143),
.B(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_89),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_94),
.A3(n_72),
.B1(n_77),
.B2(n_76),
.Y(n_131)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_135),
.A3(n_141),
.B1(n_99),
.B2(n_97),
.C(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_136),
.B(n_143),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_77),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_140),
.B(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_80),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_137),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_111),
.B1(n_116),
.B2(n_105),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_70),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_96),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_96),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_146),
.C(n_109),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_108),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_106),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_150),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_126),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_160),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_103),
.B(n_119),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_153),
.B1(n_137),
.B2(n_32),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_152),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_98),
.C(n_100),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_129),
.C(n_125),
.Y(n_179)
);

BUFx4f_ASAP7_75t_SL g159 ( 
.A(n_132),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_136),
.B(n_98),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_162),
.B(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_16),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_74),
.B(n_2),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_125),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_180),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_170),
.B1(n_160),
.B2(n_153),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_146),
.C(n_130),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_13),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_182),
.C(n_152),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_132),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_159),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_129),
.C(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_124),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_133),
.B1(n_131),
.B2(n_134),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_191),
.B1(n_161),
.B2(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_152),
.B1(n_149),
.B2(n_169),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_200),
.B(n_203),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_181),
.B1(n_189),
.B2(n_183),
.Y(n_218)
);

NOR4xp25_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_156),
.C(n_157),
.D(n_171),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_197),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_148),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_199),
.Y(n_210)
);

AOI321xp33_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_156),
.A3(n_169),
.B1(n_14),
.B2(n_13),
.C(n_12),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

FAx1_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_1),
.CI(n_2),
.CON(n_204),
.SN(n_204)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_1),
.B(n_2),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_179),
.C(n_190),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_190),
.C(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_218),
.Y(n_229)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_185),
.B(n_184),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_195),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_199),
.C(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_228),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_227),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_181),
.B(n_204),
.Y(n_226)
);

AOI31xp67_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_204),
.A3(n_219),
.B(n_211),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_203),
.C(n_4),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_221),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_230),
.A2(n_220),
.B(n_226),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_5),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_229),
.A2(n_216),
.B1(n_217),
.B2(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_5),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.C(n_240),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_3),
.B(n_4),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_231),
.B(n_8),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.C(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_10),
.C(n_6),
.Y(n_245)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_231),
.B(n_7),
.Y(n_242)
);

OAI21x1_ASAP7_75t_SL g246 ( 
.A1(n_242),
.A2(n_244),
.B(n_245),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_6),
.B(n_8),
.C(n_10),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_246),
.Y(n_249)
);


endmodule