module fake_jpeg_1867_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_17),
.B1(n_36),
.B2(n_35),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_53),
.B1(n_49),
.B2(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_0),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_52),
.B(n_1),
.Y(n_72)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_48),
.B1(n_42),
.B2(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_48),
.B1(n_42),
.B2(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_48),
.B1(n_40),
.B2(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_43),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_45),
.B(n_69),
.C(n_60),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_40),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_2),
.Y(n_96)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_67),
.Y(n_86)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_67),
.B1(n_46),
.B2(n_5),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_27),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_23),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_19),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_46),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_9),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_91),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_86),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_80),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_116),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_46),
.B(n_10),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_12),
.B(n_21),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_11),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_93),
.C(n_99),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_33),
.B(n_37),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_25),
.B1(n_34),
.B2(n_13),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_11),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_127),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_121),
.C(n_130),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_133),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_147),
.B(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_124),
.B1(n_141),
.B2(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_139),
.C(n_131),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_144),
.C(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_149),
.B1(n_137),
.B2(n_136),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_150),
.B(n_129),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_129),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_128),
.C(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_134),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_128),
.Y(n_159)
);


endmodule