module fake_netlist_1_10198_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI22xp5_ASAP7_75t_SL g11 ( .A1(n_5), .A2(n_0), .B1(n_9), .B2(n_6), .Y(n_11) );
OAI21x1_ASAP7_75t_L g12 ( .A1(n_1), .A2(n_6), .B(n_5), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
OA21x2_ASAP7_75t_L g16 ( .A1(n_4), .A2(n_0), .B(n_10), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
OR2x6_ASAP7_75t_L g18 ( .A(n_11), .B(n_1), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_2), .B(n_3), .C(n_7), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_12), .B(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVxp67_ASAP7_75t_SL g22 ( .A(n_20), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_23), .B(n_13), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_18), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_18), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AOI221x1_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_11), .B1(n_15), .B2(n_14), .C(n_13), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
NOR3xp33_ASAP7_75t_L g31 ( .A(n_28), .B(n_23), .C(n_15), .Y(n_31) );
NAND4xp25_ASAP7_75t_L g32 ( .A(n_29), .B(n_2), .C(n_3), .D(n_7), .Y(n_32) );
NAND4xp25_ASAP7_75t_SL g33 ( .A(n_29), .B(n_12), .C(n_16), .D(n_20), .Y(n_33) );
OAI22xp5_ASAP7_75t_SL g34 ( .A1(n_32), .A2(n_28), .B1(n_16), .B2(n_30), .Y(n_34) );
AO21x2_ASAP7_75t_L g35 ( .A1(n_31), .A2(n_22), .B(n_30), .Y(n_35) );
AOI21xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_16), .B(n_33), .Y(n_36) );
AOI22x1_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_34), .B1(n_16), .B2(n_22), .Y(n_37) );
endmodule