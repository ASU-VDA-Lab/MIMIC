module fake_aes_204_n_1468 (n_303, n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_302, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1468);
input n_303;
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_302;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1468;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_325;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g304 ( .A(n_159), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_74), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_86), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_237), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_269), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_72), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_236), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_268), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_188), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_172), .B(n_202), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_211), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_160), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_161), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_155), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_264), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_76), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_17), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_2), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_218), .Y(n_325) );
INVxp33_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
INVxp33_ASAP7_75t_L g327 ( .A(n_164), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_69), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_227), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_151), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_176), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_289), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_12), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_139), .Y(n_334) );
INVxp67_ASAP7_75t_SL g335 ( .A(n_97), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_251), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_240), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_279), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_135), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_107), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_186), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_95), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_119), .Y(n_343) );
INVxp33_ASAP7_75t_SL g344 ( .A(n_278), .Y(n_344) );
INVx4_ASAP7_75t_R g345 ( .A(n_233), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_71), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_60), .Y(n_347) );
CKINVDCx14_ASAP7_75t_R g348 ( .A(n_19), .Y(n_348) );
BUFx10_ASAP7_75t_L g349 ( .A(n_125), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_197), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_133), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_178), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_19), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_287), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_255), .Y(n_355) );
INVxp33_ASAP7_75t_SL g356 ( .A(n_294), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_85), .B(n_219), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_96), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_243), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_216), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_169), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_106), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_162), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_259), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_101), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_254), .Y(n_366) );
BUFx10_ASAP7_75t_L g367 ( .A(n_32), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_140), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_265), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_56), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_53), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_189), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_127), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_43), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_105), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_40), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_232), .B(n_298), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_80), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_58), .Y(n_379) );
CKINVDCx14_ASAP7_75t_R g380 ( .A(n_148), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_120), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_273), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_74), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_40), .Y(n_384) );
INVxp33_ASAP7_75t_L g385 ( .A(n_54), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_249), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_26), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_200), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_204), .Y(n_389) );
INVxp33_ASAP7_75t_SL g390 ( .A(n_92), .Y(n_390) );
INVxp33_ASAP7_75t_SL g391 ( .A(n_73), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_87), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_48), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_171), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_66), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_157), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_190), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_51), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_235), .B(n_165), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_77), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_234), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_54), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_297), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_167), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_12), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_91), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_22), .Y(n_407) );
INVxp33_ASAP7_75t_SL g408 ( .A(n_131), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_203), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_112), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_276), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_224), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_115), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_215), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_207), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_103), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_9), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_256), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_93), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_113), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_199), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_166), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_24), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_214), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_290), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_2), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_175), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_116), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_122), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_141), .Y(n_430) );
INVxp33_ASAP7_75t_L g431 ( .A(n_18), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_221), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_121), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_124), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_209), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_57), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_208), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_15), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_177), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_258), .Y(n_440) );
INVxp33_ASAP7_75t_L g441 ( .A(n_49), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_48), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_25), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_7), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_68), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_138), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_28), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g448 ( .A(n_156), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_182), .Y(n_449) );
BUFx6f_ASAP7_75t_SL g450 ( .A(n_53), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_147), .Y(n_451) );
INVxp33_ASAP7_75t_L g452 ( .A(n_26), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_181), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_98), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_210), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_143), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_8), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_31), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_82), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_9), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_180), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_411), .B(n_0), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
AND2x6_ASAP7_75t_L g465 ( .A(n_392), .B(n_88), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_366), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_326), .B(n_0), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_400), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_366), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_400), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_385), .B(n_1), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_366), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_366), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_348), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_348), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_402), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_450), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_450), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_450), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_432), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_326), .B(n_1), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_349), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_432), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_354), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_310), .B(n_3), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_354), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_338), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_368), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_350), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_385), .Y(n_494) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_368), .A2(n_90), .B(n_89), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_392), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_397), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_462), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_462), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_464), .B(n_494), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_494), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_462), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_482), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_485), .B(n_419), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_464), .B(n_375), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_469), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_485), .B(n_327), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_464), .B(n_386), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_463), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_482), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
OR2x6_ASAP7_75t_L g514 ( .A(n_471), .B(n_376), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_469), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_463), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_464), .B(n_429), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_485), .B(n_327), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_485), .B(n_322), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_471), .B(n_431), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_471), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_469), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_491), .B(n_431), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_488), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_491), .B(n_441), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_468), .B(n_322), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_468), .B(n_457), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_488), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_493), .B(n_316), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_479), .B(n_362), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_472), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_480), .B(n_389), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_490), .B(n_397), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_467), .B(n_484), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_467), .B(n_394), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_472), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_470), .B(n_474), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_472), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_470), .B(n_344), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_472), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_474), .B(n_441), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_472), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_475), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_501), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_502), .B(n_476), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_504), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_504), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_512), .B(n_489), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_499), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_521), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_511), .A2(n_484), .B(n_498), .C(n_492), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_514), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_528), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_512), .B(n_359), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_521), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_511), .A2(n_498), .B(n_492), .C(n_477), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_523), .Y(n_566) );
AO22x1_ASAP7_75t_L g567 ( .A1(n_523), .A2(n_391), .B1(n_452), .B2(n_344), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_521), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_514), .A2(n_391), .B1(n_363), .B2(n_359), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_521), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_514), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_524), .B(n_324), .Y(n_572) );
NAND3xp33_ASAP7_75t_SL g573 ( .A(n_526), .B(n_363), .C(n_371), .Y(n_573) );
BUFx12f_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_529), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_509), .B(n_520), .Y(n_576) );
INVx5_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_528), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_530), .Y(n_579) );
INVx5_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
OR2x6_ASAP7_75t_L g581 ( .A(n_547), .B(n_407), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_515), .B(n_406), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_540), .A2(n_353), .B1(n_387), .B2(n_323), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_506), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_530), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_499), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_500), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_507), .B(n_410), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_507), .B(n_425), .Y(n_589) );
NOR2x2_ASAP7_75t_L g590 ( .A(n_541), .B(n_371), .Y(n_590) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_515), .B(n_448), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_530), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_510), .B(n_306), .Y(n_593) );
INVx4_ASAP7_75t_L g594 ( .A(n_506), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_517), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_528), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_510), .B(n_306), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_518), .B(n_308), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_543), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_531), .Y(n_601) );
OAI22xp5_ASAP7_75t_SL g602 ( .A1(n_505), .A2(n_460), .B1(n_383), .B2(n_305), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_518), .B(n_308), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_540), .B(n_356), .Y(n_604) );
INVx6_ASAP7_75t_L g605 ( .A(n_531), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_533), .Y(n_606) );
NAND2x1_ASAP7_75t_L g607 ( .A(n_517), .B(n_345), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_545), .B(n_311), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_500), .B(n_304), .Y(n_609) );
NOR2x2_ASAP7_75t_L g610 ( .A(n_534), .B(n_383), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_537), .B(n_311), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_531), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_531), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_503), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_503), .A2(n_492), .B1(n_498), .B2(n_465), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_522), .A2(n_465), .B1(n_486), .B2(n_477), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_528), .Y(n_617) );
INVx2_ASAP7_75t_SL g618 ( .A(n_539), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_522), .B(n_312), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_532), .B(n_452), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_532), .B(n_312), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_539), .A2(n_353), .B1(n_387), .B2(n_323), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_536), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_536), .B(n_313), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_538), .B(n_356), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_538), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_508), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_508), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_527), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_508), .B(n_307), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_513), .B(n_390), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_513), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_513), .A2(n_495), .B(n_399), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_516), .B(n_313), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_516), .B(n_315), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_516), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_519), .B(n_447), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_519), .A2(n_495), .B(n_357), .Y(n_638) );
INVx5_ASAP7_75t_L g639 ( .A(n_527), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_525), .B(n_390), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_525), .B(n_317), .Y(n_641) );
NAND2xp33_ASAP7_75t_L g642 ( .A(n_527), .B(n_465), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_525), .B(n_329), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_535), .B(n_318), .Y(n_644) );
NAND2xp33_ASAP7_75t_SL g645 ( .A(n_527), .B(n_329), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_556), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_633), .A2(n_495), .B(n_413), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_550), .A2(n_460), .B1(n_408), .B2(n_380), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_638), .A2(n_495), .B(n_454), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_552), .B(n_340), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_566), .A2(n_558), .B(n_604), .C(n_575), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_562), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_553), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_575), .B(n_447), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_604), .A2(n_408), .B1(n_380), .B2(n_465), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_618), .B(n_309), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_600), .B(n_370), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_620), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_576), .A2(n_495), .B(n_335), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_561), .A2(n_360), .B1(n_361), .B2(n_340), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_574), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_549), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_555), .B(n_328), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_551), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_564), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_557), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_614), .B(n_360), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_558), .A2(n_320), .B(n_319), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_596), .A2(n_325), .B(n_321), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_568), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_557), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_570), .Y(n_672) );
OR2x6_ASAP7_75t_L g673 ( .A(n_563), .B(n_457), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_554), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_563), .B(n_367), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_595), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
BUFx3_ASAP7_75t_L g678 ( .A(n_605), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_554), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_577), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_584), .Y(n_681) );
BUFx8_ASAP7_75t_SL g682 ( .A(n_571), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_591), .A2(n_465), .B1(n_346), .B2(n_347), .Y(n_683) );
INVx5_ASAP7_75t_L g684 ( .A(n_605), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_596), .A2(n_331), .B(n_330), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_559), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_605), .Y(n_687) );
INVx8_ASAP7_75t_L g688 ( .A(n_581), .Y(n_688) );
OAI22xp5_ASAP7_75t_SL g689 ( .A1(n_602), .A2(n_417), .B1(n_361), .B2(n_415), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_581), .B(n_486), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_591), .A2(n_465), .B1(n_374), .B2(n_378), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_642), .A2(n_334), .B(n_332), .Y(n_692) );
OR2x6_ASAP7_75t_L g693 ( .A(n_559), .B(n_333), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_562), .Y(n_694) );
BUFx8_ASAP7_75t_L g695 ( .A(n_555), .Y(n_695) );
BUFx12f_ASAP7_75t_L g696 ( .A(n_572), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_560), .B(n_379), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_567), .A2(n_395), .B1(n_398), .B2(n_393), .C(n_384), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_588), .B(n_404), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_580), .Y(n_700) );
NOR2xp33_ASAP7_75t_R g701 ( .A(n_573), .B(n_404), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_589), .B(n_415), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_572), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_579), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_581), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_560), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_582), .A2(n_337), .B(n_336), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_582), .A2(n_341), .B(n_339), .Y(n_708) );
O2A1O1Ixp5_ASAP7_75t_SL g709 ( .A1(n_609), .A2(n_496), .B(n_342), .C(n_351), .Y(n_709) );
AND2x4_ASAP7_75t_SL g710 ( .A(n_569), .B(n_367), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_637), .Y(n_711) );
BUFx12f_ASAP7_75t_L g712 ( .A(n_606), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_622), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_583), .B(n_367), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_601), .B(n_405), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_625), .A2(n_430), .B1(n_420), .B2(n_426), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_593), .B(n_420), .Y(n_717) );
INVx4_ASAP7_75t_L g718 ( .A(n_580), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_585), .Y(n_719) );
BUFx3_ASAP7_75t_L g720 ( .A(n_562), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_592), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_590), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_601), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_634), .A2(n_377), .B(n_314), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_565), .A2(n_436), .B(n_438), .C(n_423), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_598), .B(n_430), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_613), .B(n_443), .Y(n_727) );
O2A1O1Ixp33_ASAP7_75t_SL g728 ( .A1(n_565), .A2(n_352), .B(n_355), .C(n_343), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_611), .B(n_444), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_625), .A2(n_458), .B(n_459), .C(n_445), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_613), .A2(n_465), .B1(n_497), .B2(n_349), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_608), .B(n_349), .Y(n_732) );
O2A1O1Ixp33_ASAP7_75t_L g733 ( .A1(n_612), .A2(n_496), .B(n_364), .C(n_369), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_556), .A2(n_373), .B(n_381), .C(n_358), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_562), .Y(n_735) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_586), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_599), .A2(n_388), .B(n_382), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g738 ( .A(n_610), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_586), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_587), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_587), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_623), .A2(n_401), .B(n_403), .C(n_396), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_603), .Y(n_743) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_626), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_619), .A2(n_465), .B1(n_365), .B2(n_418), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_584), .Y(n_746) );
AND2x2_ASAP7_75t_SL g747 ( .A(n_594), .B(n_409), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_627), .A2(n_414), .B(n_412), .Y(n_748) );
OAI21xp5_ASAP7_75t_L g749 ( .A1(n_609), .A2(n_465), .B(n_422), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_621), .A2(n_421), .B1(n_427), .B2(n_424), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_580), .B(n_428), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_580), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_594), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_624), .B(n_3), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_578), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_627), .A2(n_435), .B(n_434), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_597), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_607), .B(n_372), .Y(n_758) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_629), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_636), .A2(n_439), .B(n_437), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_617), .Y(n_761) );
AND2x4_ASAP7_75t_L g762 ( .A(n_631), .B(n_440), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_631), .A2(n_449), .B1(n_451), .B2(n_446), .Y(n_763) );
BUFx3_ASAP7_75t_L g764 ( .A(n_640), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_640), .B(n_455), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_636), .Y(n_766) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_639), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_645), .A2(n_461), .B1(n_433), .B2(n_453), .Y(n_768) );
INVx3_ASAP7_75t_L g769 ( .A(n_639), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_616), .A2(n_433), .B1(n_453), .B2(n_416), .Y(n_770) );
INVx4_ASAP7_75t_L g771 ( .A(n_639), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_643), .A2(n_456), .B(n_416), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_630), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_616), .B(n_4), .Y(n_774) );
O2A1O1Ixp33_ASAP7_75t_L g775 ( .A1(n_630), .A2(n_456), .B(n_481), .C(n_466), .Y(n_775) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_639), .Y(n_776) );
INVx2_ASAP7_75t_SL g777 ( .A(n_635), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_644), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_635), .A2(n_542), .B(n_535), .Y(n_779) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_628), .Y(n_780) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_628), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_644), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_641), .A2(n_497), .B1(n_483), .B2(n_487), .Y(n_783) );
NAND2xp33_ASAP7_75t_L g784 ( .A(n_615), .B(n_497), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_632), .A2(n_548), .B(n_542), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_552), .Y(n_786) );
INVx3_ASAP7_75t_L g787 ( .A(n_557), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_552), .A2(n_497), .B1(n_473), .B2(n_478), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_658), .Y(n_789) );
OAI21x1_ASAP7_75t_L g790 ( .A1(n_647), .A2(n_497), .B(n_473), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_L g791 ( .A1(n_651), .A2(n_473), .B(n_478), .C(n_472), .Y(n_791) );
OR2x6_ASAP7_75t_L g792 ( .A(n_696), .B(n_4), .Y(n_792) );
OAI21x1_ASAP7_75t_L g793 ( .A1(n_649), .A2(n_478), .B(n_473), .Y(n_793) );
OAI21xp5_ASAP7_75t_L g794 ( .A1(n_659), .A2(n_478), .B(n_473), .Y(n_794) );
NOR2x1_ASAP7_75t_SL g795 ( .A(n_693), .B(n_473), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_767), .Y(n_796) );
OA21x2_ASAP7_75t_L g797 ( .A1(n_668), .A2(n_478), .B(n_546), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_715), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_747), .A2(n_478), .B1(n_7), .B2(n_5), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_646), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_693), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_801) );
NOR2x1_ASAP7_75t_SL g802 ( .A(n_703), .B(n_10), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_715), .Y(n_803) );
AO21x2_ASAP7_75t_L g804 ( .A1(n_728), .A2(n_544), .B(n_527), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_662), .B(n_10), .Y(n_805) );
AO21x2_ASAP7_75t_L g806 ( .A1(n_784), .A2(n_544), .B(n_527), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_709), .A2(n_99), .B(n_94), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_743), .B(n_11), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_713), .B(n_11), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_711), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_724), .A2(n_546), .B(n_544), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_646), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_664), .B(n_13), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_774), .A2(n_546), .B1(n_544), .B2(n_17), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_727), .Y(n_815) );
OA21x2_ASAP7_75t_L g816 ( .A1(n_772), .A2(n_546), .B(n_544), .Y(n_816) );
OAI21x1_ASAP7_75t_SL g817 ( .A1(n_739), .A2(n_14), .B(n_16), .Y(n_817) );
OAI21x1_ASAP7_75t_L g818 ( .A1(n_785), .A2(n_102), .B(n_100), .Y(n_818) );
OAI21xp33_ASAP7_75t_SL g819 ( .A1(n_740), .A2(n_16), .B(n_18), .Y(n_819) );
AO31x2_ASAP7_75t_L g820 ( .A1(n_725), .A2(n_20), .A3(n_21), .B(n_22), .Y(n_820) );
INVx5_ASAP7_75t_L g821 ( .A(n_767), .Y(n_821) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_736), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_698), .A2(n_730), .B1(n_729), .B2(n_689), .C(n_657), .Y(n_823) );
INVxp67_ASAP7_75t_L g824 ( .A(n_653), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_673), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_674), .B(n_23), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_727), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_669), .A2(n_108), .B(n_104), .Y(n_828) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_767), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_786), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_766), .Y(n_831) );
AND2x4_ASAP7_75t_L g832 ( .A(n_679), .B(n_24), .Y(n_832) );
BUFx6f_ASAP7_75t_L g833 ( .A(n_776), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_774), .A2(n_546), .B1(n_544), .B2(n_28), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_673), .A2(n_25), .B1(n_27), .B2(n_29), .Y(n_835) );
OAI21x1_ASAP7_75t_L g836 ( .A1(n_779), .A2(n_110), .B(n_109), .Y(n_836) );
INVxp67_ASAP7_75t_L g837 ( .A(n_686), .Y(n_837) );
INVxp67_ASAP7_75t_L g838 ( .A(n_706), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_766), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_741), .A2(n_27), .B1(n_29), .B2(n_30), .Y(n_840) );
OAI21x1_ASAP7_75t_L g841 ( .A1(n_692), .A2(n_114), .B(n_111), .Y(n_841) );
NOR2x1_ASAP7_75t_R g842 ( .A(n_712), .B(n_30), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_697), .B(n_31), .Y(n_843) );
OAI21x1_ASAP7_75t_L g844 ( .A1(n_749), .A2(n_118), .B(n_117), .Y(n_844) );
OR2x2_ASAP7_75t_L g845 ( .A(n_688), .B(n_32), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_690), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_655), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_847) );
INVx3_ASAP7_75t_L g848 ( .A(n_753), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_753), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g850 ( .A(n_736), .B(n_546), .Y(n_850) );
OAI21x1_ASAP7_75t_SL g851 ( .A1(n_718), .A2(n_33), .B(n_34), .Y(n_851) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_763), .A2(n_35), .B1(n_36), .B2(n_37), .C(n_38), .Y(n_852) );
OA21x2_ASAP7_75t_L g853 ( .A1(n_765), .A2(n_126), .B(n_123), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_746), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g855 ( .A1(n_742), .A2(n_36), .B1(n_37), .B2(n_38), .C(n_39), .Y(n_855) );
NAND2xp33_ASAP7_75t_R g856 ( .A(n_705), .B(n_39), .Y(n_856) );
BUFx2_ASAP7_75t_SL g857 ( .A(n_661), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_736), .Y(n_858) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_769), .A2(n_129), .B(n_128), .Y(n_859) );
CKINVDCx6p67_ASAP7_75t_R g860 ( .A(n_688), .Y(n_860) );
INVx2_ASAP7_75t_SL g861 ( .A(n_695), .Y(n_861) );
O2A1O1Ixp33_ASAP7_75t_L g862 ( .A1(n_734), .A2(n_41), .B(n_42), .C(n_43), .Y(n_862) );
AO21x2_ASAP7_75t_L g863 ( .A1(n_770), .A2(n_132), .B(n_130), .Y(n_863) );
NAND2x1p5_ASAP7_75t_L g864 ( .A(n_753), .B(n_41), .Y(n_864) );
OAI22xp33_ASAP7_75t_SL g865 ( .A1(n_738), .A2(n_42), .B1(n_44), .B2(n_45), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g866 ( .A(n_732), .B(n_44), .C(n_45), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_759), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_683), .A2(n_46), .B1(n_47), .B2(n_49), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_654), .B(n_46), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_691), .A2(n_47), .B1(n_50), .B2(n_51), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_656), .Y(n_871) );
INVxp67_ASAP7_75t_L g872 ( .A(n_697), .Y(n_872) );
BUFx2_ASAP7_75t_L g873 ( .A(n_695), .Y(n_873) );
AO31x2_ASAP7_75t_L g874 ( .A1(n_750), .A2(n_50), .A3(n_52), .B(n_55), .Y(n_874) );
OA21x2_ASAP7_75t_L g875 ( .A1(n_737), .A2(n_195), .B(n_302), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_682), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_665), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_663), .B(n_52), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_755), .A2(n_194), .B(n_301), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_764), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_880) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_685), .A2(n_198), .B(n_300), .Y(n_881) );
AO31x2_ASAP7_75t_L g882 ( .A1(n_704), .A2(n_58), .A3(n_59), .B(n_60), .Y(n_882) );
OA21x2_ASAP7_75t_L g883 ( .A1(n_788), .A2(n_201), .B(n_299), .Y(n_883) );
OA21x2_ASAP7_75t_L g884 ( .A1(n_707), .A2(n_708), .B(n_731), .Y(n_884) );
AO21x2_ASAP7_75t_L g885 ( .A1(n_768), .A2(n_196), .B(n_296), .Y(n_885) );
INVx4_ASAP7_75t_L g886 ( .A(n_776), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_744), .Y(n_887) );
AO21x2_ASAP7_75t_L g888 ( .A1(n_748), .A2(n_193), .B(n_293), .Y(n_888) );
INVx4_ASAP7_75t_L g889 ( .A(n_776), .Y(n_889) );
AO21x2_ASAP7_75t_L g890 ( .A1(n_756), .A2(n_192), .B(n_291), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_744), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_762), .A2(n_59), .B1(n_61), .B2(n_62), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_710), .B(n_61), .Y(n_893) );
OAI21x1_ASAP7_75t_SL g894 ( .A1(n_718), .A2(n_62), .B(n_63), .Y(n_894) );
AO32x2_ASAP7_75t_L g895 ( .A1(n_777), .A2(n_63), .A3(n_64), .B1(n_65), .B2(n_66), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_699), .A2(n_64), .B1(n_65), .B2(n_67), .Y(n_896) );
INVx3_ASAP7_75t_L g897 ( .A(n_771), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_744), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_719), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_670), .Y(n_900) );
BUFx3_ASAP7_75t_L g901 ( .A(n_759), .Y(n_901) );
AND2x4_ASAP7_75t_L g902 ( .A(n_684), .B(n_67), .Y(n_902) );
AO31x2_ASAP7_75t_L g903 ( .A1(n_721), .A2(n_68), .A3(n_69), .B(n_70), .Y(n_903) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_761), .A2(n_212), .B(n_288), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_652), .Y(n_905) );
OAI21x1_ASAP7_75t_L g906 ( .A1(n_775), .A2(n_206), .B(n_286), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_760), .A2(n_205), .B(n_285), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_778), .A2(n_191), .B(n_284), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_778), .A2(n_187), .B(n_283), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_672), .Y(n_910) );
O2A1O1Ixp33_ASAP7_75t_SL g911 ( .A1(n_782), .A2(n_185), .B(n_281), .C(n_280), .Y(n_911) );
AOI22xp5_ASAP7_75t_SL g912 ( .A1(n_722), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_782), .A2(n_213), .B(n_277), .Y(n_913) );
BUFx3_ASAP7_75t_L g914 ( .A(n_759), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_762), .A2(n_73), .B1(n_75), .B2(n_76), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g916 ( .A1(n_773), .A2(n_217), .B(n_275), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_714), .B(n_75), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_663), .A2(n_77), .B1(n_78), .B2(n_79), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_702), .B(n_78), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_723), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_648), .B(n_716), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_687), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_717), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_923) );
AO21x2_ASAP7_75t_L g924 ( .A1(n_754), .A2(n_220), .B(n_274), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_701), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_676), .Y(n_926) );
INVx6_ASAP7_75t_L g927 ( .A(n_684), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_675), .B(n_81), .Y(n_928) );
OAI21x1_ASAP7_75t_L g929 ( .A1(n_681), .A2(n_222), .B(n_272), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_677), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_751), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_931) );
INVx3_ASAP7_75t_L g932 ( .A(n_771), .Y(n_932) );
NOR2xp67_ASAP7_75t_L g933 ( .A(n_660), .B(n_83), .Y(n_933) );
OAI21x1_ASAP7_75t_L g934 ( .A1(n_681), .A2(n_223), .B(n_134), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_726), .A2(n_84), .B1(n_136), .B2(n_137), .Y(n_935) );
AND2x4_ASAP7_75t_L g936 ( .A(n_684), .B(n_303), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_667), .A2(n_142), .B1(n_144), .B2(n_145), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_678), .B(n_146), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_650), .B(n_787), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_733), .A2(n_149), .B1(n_150), .B2(n_152), .C(n_153), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_751), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_780), .Y(n_942) );
AOI21xp5_ASAP7_75t_L g943 ( .A1(n_758), .A2(n_154), .B(n_158), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_752), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_823), .B(n_787), .Y(n_945) );
AOI21xp5_ASAP7_75t_L g946 ( .A1(n_794), .A2(n_652), .B(n_694), .Y(n_946) );
NOR2x1_ASAP7_75t_R g947 ( .A(n_876), .B(n_720), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_814), .A2(n_757), .B1(n_745), .B2(n_652), .Y(n_948) );
O2A1O1Ixp33_ASAP7_75t_L g949 ( .A1(n_921), .A2(n_666), .B(n_671), .C(n_700), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_823), .A2(n_666), .B1(n_671), .B2(n_680), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_809), .A2(n_735), .B1(n_781), .B2(n_780), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_809), .A2(n_781), .B1(n_780), .B2(n_694), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_832), .A2(n_781), .B1(n_694), .B2(n_783), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_831), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_837), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_813), .B(n_163), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_877), .B(n_168), .Y(n_957) );
BUFx2_ASAP7_75t_L g958 ( .A(n_792), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_872), .B(n_170), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_871), .B(n_271), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_789), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_837), .B(n_173), .Y(n_962) );
A2O1A1Ixp33_ASAP7_75t_L g963 ( .A1(n_933), .A2(n_174), .B(n_179), .C(n_183), .Y(n_963) );
NOR2xp33_ASAP7_75t_R g964 ( .A(n_860), .B(n_856), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_850), .A2(n_184), .B(n_225), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_838), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_846), .Y(n_967) );
AOI21xp5_ASAP7_75t_L g968 ( .A1(n_850), .A2(n_226), .B(n_228), .Y(n_968) );
AO21x2_ASAP7_75t_L g969 ( .A1(n_791), .A2(n_229), .B(n_230), .Y(n_969) );
OAI221xp5_ASAP7_75t_SL g970 ( .A1(n_792), .A2(n_231), .B1(n_238), .B2(n_239), .C(n_241), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_838), .Y(n_971) );
INVx3_ASAP7_75t_L g972 ( .A(n_821), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_832), .A2(n_242), .B1(n_244), .B2(n_246), .Y(n_973) );
AND2x4_ASAP7_75t_L g974 ( .A(n_821), .B(n_247), .Y(n_974) );
BUFx2_ASAP7_75t_L g975 ( .A(n_792), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_839), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g977 ( .A1(n_912), .A2(n_248), .B1(n_250), .B2(n_252), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_917), .A2(n_253), .B1(n_257), .B2(n_260), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_856), .Y(n_979) );
NAND3xp33_ASAP7_75t_L g980 ( .A(n_866), .B(n_261), .C(n_262), .Y(n_980) );
OA21x2_ASAP7_75t_L g981 ( .A1(n_791), .A2(n_263), .B(n_266), .Y(n_981) );
AOI221xp5_ASAP7_75t_L g982 ( .A1(n_825), .A2(n_267), .B1(n_270), .B2(n_835), .C(n_852), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_900), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_824), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_830), .Y(n_985) );
NOR2xp33_ASAP7_75t_L g986 ( .A(n_872), .B(n_824), .Y(n_986) );
AOI221xp5_ASAP7_75t_L g987 ( .A1(n_825), .A2(n_835), .B1(n_852), .B2(n_893), .C(n_826), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_800), .Y(n_988) );
AND2x4_ASAP7_75t_L g989 ( .A(n_821), .B(n_886), .Y(n_989) );
OR2x6_ASAP7_75t_L g990 ( .A(n_857), .B(n_873), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_893), .A2(n_802), .B1(n_795), .B2(n_826), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_928), .A2(n_869), .B1(n_805), .B2(n_799), .Y(n_992) );
OA21x2_ASAP7_75t_L g993 ( .A1(n_790), .A2(n_793), .B(n_807), .Y(n_993) );
AOI21xp5_ASAP7_75t_L g994 ( .A1(n_806), .A2(n_816), .B(n_919), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_798), .A2(n_815), .B1(n_827), .B2(n_803), .C(n_810), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_899), .B(n_910), .Y(n_996) );
AO21x2_ASAP7_75t_L g997 ( .A1(n_804), .A2(n_806), .B(n_916), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_925), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_926), .Y(n_999) );
NOR2x1_ASAP7_75t_L g1000 ( .A(n_845), .B(n_901), .Y(n_1000) );
INVx3_ASAP7_75t_L g1001 ( .A(n_821), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_854), .B(n_812), .Y(n_1002) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_861), .B(n_854), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_808), .B(n_930), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_878), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_892), .B(n_915), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_902), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_843), .A2(n_847), .B1(n_834), .B2(n_814), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_834), .A2(n_915), .B1(n_892), .B2(n_931), .Y(n_1009) );
OAI322xp33_ASAP7_75t_L g1010 ( .A1(n_855), .A2(n_801), .A3(n_840), .B1(n_896), .B2(n_923), .C1(n_862), .C2(n_868), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_944), .B(n_941), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_865), .A2(n_855), .B1(n_862), .B2(n_870), .C(n_819), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_918), .A2(n_931), .B1(n_880), .B2(n_939), .C(n_940), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_864), .A2(n_918), .B1(n_880), .B2(n_940), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_867), .B(n_902), .Y(n_1015) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_901), .Y(n_1016) );
OAI22xp33_ASAP7_75t_L g1017 ( .A1(n_864), .A2(n_914), .B1(n_867), .B2(n_897), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_816), .A2(n_822), .B(n_811), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_936), .A2(n_822), .B1(n_811), .B2(n_914), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_920), .B(n_939), .Y(n_1020) );
AOI21xp5_ASAP7_75t_L g1021 ( .A1(n_816), .A2(n_811), .B(n_797), .Y(n_1021) );
AOI222xp33_ASAP7_75t_L g1022 ( .A1(n_842), .A2(n_922), .B1(n_894), .B2(n_851), .C1(n_817), .C2(n_935), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_874), .Y(n_1023) );
AOI21xp5_ASAP7_75t_L g1024 ( .A1(n_797), .A2(n_804), .B(n_884), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g1025 ( .A1(n_797), .A2(n_884), .B(n_911), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1026 ( .A1(n_943), .A2(n_907), .B1(n_881), .B2(n_828), .C(n_913), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_829), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_897), .A2(n_932), .B1(n_936), .B2(n_927), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_932), .A2(n_927), .B1(n_884), .B2(n_938), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_927), .A2(n_796), .B1(n_849), .B2(n_848), .Y(n_1030) );
BUFx4f_ASAP7_75t_SL g1031 ( .A(n_886), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_874), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_874), .B(n_889), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_829), .Y(n_1034) );
AO21x1_ASAP7_75t_L g1035 ( .A1(n_908), .A2(n_913), .B(n_943), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_848), .B(n_849), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_858), .B(n_898), .Y(n_1037) );
INVxp67_ASAP7_75t_SL g1038 ( .A(n_829), .Y(n_1038) );
AOI21xp5_ASAP7_75t_L g1039 ( .A1(n_911), .A2(n_907), .B(n_905), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_889), .Y(n_1040) );
AND2x6_ASAP7_75t_L g1041 ( .A(n_829), .B(n_833), .Y(n_1041) );
AOI21xp5_ASAP7_75t_L g1042 ( .A1(n_905), .A2(n_908), .B(n_853), .Y(n_1042) );
NAND2xp5_ASAP7_75t_SL g1043 ( .A(n_833), .B(n_796), .Y(n_1043) );
AOI21xp5_ASAP7_75t_L g1044 ( .A1(n_853), .A2(n_875), .B(n_942), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_833), .Y(n_1045) );
AO221x2_ASAP7_75t_L g1046 ( .A1(n_895), .A2(n_903), .B1(n_882), .B2(n_874), .C(n_820), .Y(n_1046) );
OAI221xp5_ASAP7_75t_L g1047 ( .A1(n_937), .A2(n_875), .B1(n_853), .B2(n_891), .C(n_887), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_924), .A2(n_833), .B1(n_890), .B2(n_888), .Y(n_1048) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_882), .Y(n_1049) );
OR2x6_ASAP7_75t_L g1050 ( .A(n_929), .B(n_934), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_924), .A2(n_888), .B1(n_890), .B2(n_863), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_863), .A2(n_885), .B1(n_875), .B2(n_883), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_883), .A2(n_895), .B1(n_820), .B2(n_882), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_820), .B(n_882), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_820), .Y(n_1055) );
INVx3_ASAP7_75t_L g1056 ( .A(n_859), .Y(n_1056) );
AOI222xp33_ASAP7_75t_L g1057 ( .A1(n_895), .A2(n_903), .B1(n_909), .B2(n_879), .C1(n_904), .C2(n_841), .Y(n_1057) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_903), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_885), .A2(n_883), .B1(n_844), .B2(n_906), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_903), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g1061 ( .A(n_818), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1062 ( .A1(n_836), .A2(n_649), .B(n_647), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_895), .A2(n_814), .B1(n_834), .B2(n_747), .Y(n_1063) );
A2O1A1Ixp33_ASAP7_75t_L g1064 ( .A1(n_933), .A2(n_651), .B(n_819), .C(n_866), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_823), .A2(n_722), .B1(n_602), .B2(n_673), .Y(n_1065) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_876), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_789), .Y(n_1067) );
AOI21xp5_ASAP7_75t_L g1068 ( .A1(n_794), .A2(n_649), .B(n_647), .Y(n_1068) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_791), .A2(n_651), .B(n_659), .Y(n_1069) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_821), .B(n_703), .Y(n_1070) );
INVx4_ASAP7_75t_SL g1071 ( .A(n_792), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_823), .A2(n_722), .B1(n_602), .B2(n_673), .Y(n_1072) );
NAND2x1_ASAP7_75t_L g1073 ( .A(n_886), .B(n_889), .Y(n_1073) );
OAI211xp5_ASAP7_75t_L g1074 ( .A1(n_823), .A2(n_698), .B(n_722), .C(n_892), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g1075 ( .A1(n_823), .A2(n_698), .B1(n_602), .B2(n_664), .C(n_662), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g1076 ( .A(n_876), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_789), .Y(n_1077) );
NOR3xp33_ASAP7_75t_SL g1078 ( .A(n_925), .B(n_738), .C(n_856), .Y(n_1078) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_837), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_837), .B(n_575), .Y(n_1080) );
INVx6_ASAP7_75t_L g1081 ( .A(n_821), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_831), .Y(n_1082) );
INVx6_ASAP7_75t_L g1083 ( .A(n_821), .Y(n_1083) );
INVx2_ASAP7_75t_SL g1084 ( .A(n_860), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g1085 ( .A1(n_823), .A2(n_698), .B1(n_602), .B2(n_664), .C(n_662), .Y(n_1085) );
OAI211xp5_ASAP7_75t_SL g1086 ( .A1(n_823), .A2(n_698), .B(n_662), .C(n_664), .Y(n_1086) );
INVx4_ASAP7_75t_L g1087 ( .A(n_792), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_988), .B(n_954), .Y(n_1088) );
INVx3_ASAP7_75t_L g1089 ( .A(n_1041), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1056), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_993), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1075), .B(n_1085), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1060), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1023), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_996), .Y(n_1095) );
AOI221xp5_ASAP7_75t_L g1096 ( .A1(n_1086), .A2(n_1072), .B1(n_1065), .B2(n_987), .C(n_1074), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_984), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1082), .B(n_976), .Y(n_1098) );
BUFx3_ASAP7_75t_L g1099 ( .A(n_989), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_996), .B(n_983), .Y(n_1100) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_989), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1006), .B(n_961), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_982), .A2(n_1009), .B1(n_1087), .B2(n_1013), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1002), .B(n_1032), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1067), .B(n_1077), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1055), .Y(n_1106) );
INVxp67_ASAP7_75t_R g1107 ( .A(n_1071), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_999), .B(n_950), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1080), .B(n_967), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1015), .B(n_945), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_985), .B(n_986), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1005), .B(n_1020), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1020), .B(n_1054), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1033), .B(n_972), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1054), .Y(n_1115) );
INVx1_ASAP7_75t_SL g1116 ( .A(n_1040), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_955), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1049), .Y(n_1118) );
INVxp67_ASAP7_75t_SL g1119 ( .A(n_1019), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_966), .B(n_971), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1058), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1079), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1003), .B(n_995), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g1124 ( .A(n_1076), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1046), .Y(n_1125) );
INVx1_ASAP7_75t_SL g1126 ( .A(n_1031), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_972), .B(n_1001), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_992), .A2(n_1087), .B1(n_1063), .B2(n_1009), .Y(n_1128) );
INVxp67_ASAP7_75t_SL g1129 ( .A(n_1019), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1046), .B(n_1063), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1027), .Y(n_1131) );
INVx3_ASAP7_75t_L g1132 ( .A(n_1041), .Y(n_1132) );
OAI33xp33_ASAP7_75t_L g1133 ( .A1(n_1053), .A2(n_979), .A3(n_1014), .B1(n_1004), .B2(n_1007), .B3(n_1011), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1001), .B(n_1070), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_997), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1070), .B(n_1016), .Y(n_1136) );
OA21x2_ASAP7_75t_L g1137 ( .A1(n_1025), .A2(n_1024), .B(n_1021), .Y(n_1137) );
BUFx3_ASAP7_75t_L g1138 ( .A(n_1081), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_1041), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1071), .B(n_974), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_991), .B(n_958), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_990), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1053), .B(n_975), .Y(n_1143) );
INVx2_ASAP7_75t_L g1144 ( .A(n_1061), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1037), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_1012), .A2(n_1014), .B1(n_1071), .B2(n_1022), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_974), .B(n_1028), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_957), .B(n_1022), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1037), .Y(n_1149) );
INVx4_ASAP7_75t_L g1150 ( .A(n_1041), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_957), .Y(n_1151) );
BUFx6f_ASAP7_75t_L g1152 ( .A(n_1050), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_1010), .A2(n_1008), .B1(n_948), .B2(n_964), .Y(n_1153) );
INVx3_ASAP7_75t_SL g1154 ( .A(n_990), .Y(n_1154) );
INVx3_ASAP7_75t_L g1155 ( .A(n_1081), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1000), .B(n_1084), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_990), .B(n_1078), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1064), .B(n_1036), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1034), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1050), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1045), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1057), .Y(n_1162) );
INVxp67_ASAP7_75t_SL g1163 ( .A(n_1017), .Y(n_1163) );
OAI21xp5_ASAP7_75t_L g1164 ( .A1(n_948), .A2(n_949), .B(n_1026), .Y(n_1164) );
AOI22xp33_ASAP7_75t_SL g1165 ( .A1(n_1083), .A2(n_962), .B1(n_981), .B2(n_969), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1083), .B(n_956), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1030), .B(n_1069), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1057), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1169 ( .A(n_1073), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1069), .B(n_1038), .Y(n_1170) );
INVx3_ASAP7_75t_SL g1171 ( .A(n_1066), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_953), .A2(n_970), .B1(n_977), .B2(n_973), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1029), .B(n_969), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_1043), .Y(n_1174) );
BUFx3_ASAP7_75t_L g1175 ( .A(n_1050), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_960), .B(n_951), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_981), .B(n_952), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1178 ( .A(n_1018), .B(n_1051), .Y(n_1178) );
AND2x4_ASAP7_75t_L g1179 ( .A(n_946), .B(n_1068), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_994), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_959), .B(n_1048), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1047), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1052), .B(n_1044), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_947), .B(n_978), .Y(n_1184) );
AND2x4_ASAP7_75t_SL g1185 ( .A(n_1059), .B(n_963), .Y(n_1185) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1035), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_980), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1062), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_1042), .B(n_1039), .Y(n_1189) );
INVx2_ASAP7_75t_L g1190 ( .A(n_965), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_968), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1113), .B(n_998), .Y(n_1192) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1150), .Y(n_1193) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1117), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1102), .B(n_1114), .Y(n_1195) );
OAI221xp5_ASAP7_75t_L g1196 ( .A1(n_1096), .A2(n_1146), .B1(n_1092), .B2(n_1153), .C(n_1103), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1105), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1113), .B(n_1130), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1122), .Y(n_1199) );
AND2x4_ASAP7_75t_L g1200 ( .A(n_1114), .B(n_1175), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_1097), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1094), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1130), .B(n_1143), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1102), .B(n_1125), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1094), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1125), .B(n_1162), .Y(n_1206) );
OR2x2_ASAP7_75t_SL g1207 ( .A(n_1143), .B(n_1142), .Y(n_1207) );
OAI31xp33_ASAP7_75t_L g1208 ( .A1(n_1128), .A2(n_1148), .A3(n_1123), .B(n_1141), .Y(n_1208) );
BUFx3_ASAP7_75t_L g1209 ( .A(n_1099), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1106), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1112), .B(n_1100), .Y(n_1211) );
AOI33xp33_ASAP7_75t_L g1212 ( .A1(n_1112), .A2(n_1162), .A3(n_1168), .B1(n_1105), .B2(n_1148), .B3(n_1100), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1168), .B(n_1115), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1106), .Y(n_1214) );
INVx4_ASAP7_75t_L g1215 ( .A(n_1154), .Y(n_1215) );
BUFx2_ASAP7_75t_L g1216 ( .A(n_1152), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1091), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1115), .B(n_1167), .Y(n_1218) );
OAI33xp33_ASAP7_75t_L g1219 ( .A1(n_1120), .A2(n_1111), .A3(n_1156), .B1(n_1157), .B2(n_1109), .B3(n_1104), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1098), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1098), .B(n_1110), .Y(n_1221) );
AND2x4_ASAP7_75t_L g1222 ( .A(n_1160), .B(n_1093), .Y(n_1222) );
AND2x2_ASAP7_75t_SL g1223 ( .A(n_1150), .B(n_1139), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1116), .B(n_1126), .Y(n_1224) );
INVx1_ASAP7_75t_SL g1225 ( .A(n_1154), .Y(n_1225) );
INVx3_ASAP7_75t_L g1226 ( .A(n_1150), .Y(n_1226) );
AND2x4_ASAP7_75t_L g1227 ( .A(n_1093), .B(n_1089), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1099), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1229 ( .A1(n_1184), .A2(n_1154), .B1(n_1164), .B2(n_1172), .C(n_1163), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1167), .B(n_1110), .Y(n_1230) );
AOI31xp33_ASAP7_75t_L g1231 ( .A1(n_1140), .A2(n_1107), .A3(n_1169), .B(n_1147), .Y(n_1231) );
AND2x4_ASAP7_75t_L g1232 ( .A(n_1089), .B(n_1132), .Y(n_1232) );
INVx4_ASAP7_75t_L g1233 ( .A(n_1150), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_1101), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1104), .B(n_1095), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1107), .A2(n_1140), .B1(n_1147), .B2(n_1101), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_1158), .A2(n_1108), .B1(n_1133), .B2(n_1181), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1088), .B(n_1170), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1145), .B(n_1149), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1088), .B(n_1108), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1118), .Y(n_1241) );
OAI31xp33_ASAP7_75t_L g1242 ( .A1(n_1158), .A2(n_1166), .A3(n_1185), .B(n_1151), .Y(n_1242) );
OR2x6_ASAP7_75t_L g1243 ( .A(n_1152), .B(n_1139), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1170), .B(n_1149), .Y(n_1244) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_1101), .Y(n_1245) );
OAI33xp33_ASAP7_75t_L g1246 ( .A1(n_1178), .A2(n_1180), .A3(n_1183), .B1(n_1121), .B2(n_1118), .B3(n_1145), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1136), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1121), .B(n_1178), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1180), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1159), .Y(n_1250) );
INVx2_ASAP7_75t_SL g1251 ( .A(n_1089), .Y(n_1251) );
AND2x4_ASAP7_75t_SL g1252 ( .A(n_1134), .B(n_1136), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1159), .B(n_1161), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1119), .B(n_1129), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1161), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_1152), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1166), .B(n_1134), .Y(n_1257) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_1151), .A2(n_1181), .B1(n_1176), .B2(n_1127), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1238), .B(n_1173), .Y(n_1259) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1217), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1238), .B(n_1173), .Y(n_1261) );
NOR2x1_ASAP7_75t_L g1262 ( .A(n_1215), .B(n_1132), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1197), .B(n_1127), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1194), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1218), .B(n_1186), .Y(n_1265) );
BUFx3_ASAP7_75t_L g1266 ( .A(n_1209), .Y(n_1266) );
NAND4xp25_ASAP7_75t_L g1267 ( .A(n_1208), .B(n_1165), .C(n_1186), .D(n_1183), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1199), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1218), .B(n_1186), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1203), .B(n_1186), .Y(n_1270) );
INVx6_ASAP7_75t_L g1271 ( .A(n_1215), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1244), .B(n_1144), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1244), .B(n_1144), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1195), .B(n_1144), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1195), .B(n_1182), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1220), .B(n_1131), .Y(n_1276) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_1201), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1202), .Y(n_1278) );
BUFx2_ASAP7_75t_L g1279 ( .A(n_1243), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1224), .B(n_1171), .Y(n_1280) );
OR2x6_ASAP7_75t_L g1281 ( .A(n_1233), .B(n_1152), .Y(n_1281) );
AND2x4_ASAP7_75t_L g1282 ( .A(n_1227), .B(n_1152), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1203), .B(n_1188), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1202), .Y(n_1284) );
NAND2x1p5_ASAP7_75t_L g1285 ( .A(n_1233), .B(n_1089), .Y(n_1285) );
NAND4xp25_ASAP7_75t_L g1286 ( .A(n_1242), .B(n_1229), .C(n_1237), .D(n_1196), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1205), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1213), .B(n_1182), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1230), .B(n_1131), .Y(n_1289) );
INVx4_ASAP7_75t_L g1290 ( .A(n_1215), .Y(n_1290) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_1192), .A2(n_1171), .B1(n_1155), .B2(n_1182), .C(n_1138), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1205), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1230), .B(n_1174), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1213), .B(n_1188), .Y(n_1294) );
INVx2_ASAP7_75t_SL g1295 ( .A(n_1252), .Y(n_1295) );
AND2x4_ASAP7_75t_L g1296 ( .A(n_1227), .B(n_1179), .Y(n_1296) );
NOR2xp33_ASAP7_75t_R g1297 ( .A(n_1223), .B(n_1124), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1298 ( .A(n_1192), .B(n_1179), .C(n_1189), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1206), .B(n_1179), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1206), .B(n_1179), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1198), .B(n_1189), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1228), .Y(n_1302) );
NAND5xp2_ASAP7_75t_SL g1303 ( .A(n_1223), .B(n_1171), .C(n_1177), .D(n_1176), .E(n_1185), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_1211), .B(n_1155), .Y(n_1304) );
NAND2xp33_ASAP7_75t_SL g1305 ( .A(n_1212), .B(n_1132), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1204), .B(n_1137), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1204), .B(n_1137), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1210), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1210), .Y(n_1309) );
NAND4xp25_ASAP7_75t_L g1310 ( .A(n_1258), .B(n_1138), .C(n_1177), .D(n_1155), .Y(n_1310) );
AOI21xp5_ASAP7_75t_SL g1311 ( .A1(n_1231), .A2(n_1138), .B(n_1090), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1214), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1222), .B(n_1137), .Y(n_1313) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1198), .B(n_1135), .Y(n_1314) );
OAI21xp33_ASAP7_75t_L g1315 ( .A1(n_1248), .A2(n_1185), .B(n_1191), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1221), .B(n_1155), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g1317 ( .A(n_1234), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1275), .B(n_1240), .Y(n_1318) );
NOR3xp33_ASAP7_75t_L g1319 ( .A(n_1286), .B(n_1219), .C(n_1225), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1277), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1264), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1301), .B(n_1248), .Y(n_1322) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_1266), .Y(n_1323) );
OAI21xp5_ASAP7_75t_SL g1324 ( .A1(n_1310), .A2(n_1252), .B(n_1236), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1299), .B(n_1222), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1268), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1301), .B(n_1254), .Y(n_1327) );
BUFx2_ASAP7_75t_L g1328 ( .A(n_1297), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1299), .B(n_1222), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1278), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1284), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1300), .B(n_1200), .Y(n_1332) );
OR3x2_ASAP7_75t_L g1333 ( .A(n_1267), .B(n_1235), .C(n_1239), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1300), .B(n_1200), .Y(n_1334) );
CKINVDCx16_ASAP7_75t_R g1335 ( .A(n_1295), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1275), .B(n_1247), .Y(n_1336) );
NAND2xp5_ASAP7_75t_SL g1337 ( .A(n_1290), .B(n_1233), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1259), .B(n_1200), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1287), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1259), .B(n_1241), .Y(n_1340) );
BUFx2_ASAP7_75t_L g1341 ( .A(n_1266), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1283), .B(n_1254), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1292), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1308), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1309), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1294), .B(n_1253), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1294), .B(n_1253), .Y(n_1347) );
INVx2_ASAP7_75t_L g1348 ( .A(n_1260), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1274), .B(n_1241), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1283), .B(n_1314), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1312), .Y(n_1351) );
INVx1_ASAP7_75t_SL g1352 ( .A(n_1295), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g1353 ( .A(n_1280), .B(n_1257), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1314), .B(n_1235), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1274), .Y(n_1355) );
INVx1_ASAP7_75t_SL g1356 ( .A(n_1271), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1270), .B(n_1207), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1261), .B(n_1249), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1293), .B(n_1214), .Y(n_1359) );
INVx1_ASAP7_75t_SL g1360 ( .A(n_1271), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1270), .B(n_1207), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1289), .B(n_1255), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1288), .B(n_1250), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1350), .B(n_1306), .Y(n_1364) );
NOR2xp33_ASAP7_75t_SL g1365 ( .A(n_1335), .B(n_1290), .Y(n_1365) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1348), .Y(n_1366) );
AOI211xp5_ASAP7_75t_SL g1367 ( .A1(n_1324), .A2(n_1311), .B(n_1291), .C(n_1315), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1330), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1331), .Y(n_1369) );
OAI322xp33_ASAP7_75t_L g1370 ( .A1(n_1327), .A2(n_1316), .A3(n_1263), .B1(n_1298), .B2(n_1304), .C1(n_1261), .C2(n_1276), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1339), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1340), .B(n_1306), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1358), .B(n_1307), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1343), .Y(n_1374) );
AOI22xp5_ASAP7_75t_L g1375 ( .A1(n_1333), .A2(n_1305), .B1(n_1269), .B2(n_1265), .Y(n_1375) );
HB1xp67_ASAP7_75t_L g1376 ( .A(n_1341), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1344), .Y(n_1377) );
AOI22xp5_ASAP7_75t_L g1378 ( .A1(n_1333), .A2(n_1305), .B1(n_1269), .B2(n_1265), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1350), .Y(n_1379) );
INVxp67_ASAP7_75t_L g1380 ( .A(n_1341), .Y(n_1380) );
INVx1_ASAP7_75t_SL g1381 ( .A(n_1352), .Y(n_1381) );
OAI21xp33_ASAP7_75t_L g1382 ( .A1(n_1319), .A2(n_1311), .B(n_1307), .Y(n_1382) );
INVxp67_ASAP7_75t_L g1383 ( .A(n_1328), .Y(n_1383) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1348), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1321), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1358), .B(n_1313), .Y(n_1386) );
INVx1_ASAP7_75t_SL g1387 ( .A(n_1323), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1340), .B(n_1288), .Y(n_1388) );
INVx1_ASAP7_75t_SL g1389 ( .A(n_1323), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1320), .B(n_1317), .Y(n_1390) );
INVx2_ASAP7_75t_L g1391 ( .A(n_1345), .Y(n_1391) );
O2A1O1Ixp33_ASAP7_75t_L g1392 ( .A1(n_1337), .A2(n_1302), .B(n_1303), .C(n_1245), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1327), .B(n_1272), .Y(n_1393) );
AOI22xp5_ASAP7_75t_L g1394 ( .A1(n_1337), .A2(n_1296), .B1(n_1271), .B2(n_1272), .Y(n_1394) );
INVx2_ASAP7_75t_L g1395 ( .A(n_1351), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1391), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1391), .Y(n_1397) );
INVx1_ASAP7_75t_SL g1398 ( .A(n_1387), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1373), .B(n_1355), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1395), .Y(n_1400) );
XOR2x2_ASAP7_75t_L g1401 ( .A(n_1367), .B(n_1353), .Y(n_1401) );
XNOR2x1_ASAP7_75t_L g1402 ( .A(n_1381), .B(n_1326), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1373), .B(n_1346), .Y(n_1403) );
NAND2xp5_ASAP7_75t_SL g1404 ( .A(n_1365), .B(n_1356), .Y(n_1404) );
AOI21xp33_ASAP7_75t_SL g1405 ( .A1(n_1382), .A2(n_1285), .B(n_1361), .Y(n_1405) );
NAND2x1_ASAP7_75t_L g1406 ( .A(n_1394), .B(n_1271), .Y(n_1406) );
INVxp67_ASAP7_75t_SL g1407 ( .A(n_1376), .Y(n_1407) );
AOI21xp5_ASAP7_75t_L g1408 ( .A1(n_1392), .A2(n_1303), .B(n_1290), .Y(n_1408) );
INVx3_ASAP7_75t_L g1409 ( .A(n_1389), .Y(n_1409) );
AOI32xp33_ASAP7_75t_L g1410 ( .A1(n_1386), .A2(n_1338), .A3(n_1360), .B1(n_1332), .B2(n_1334), .Y(n_1410) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1366), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1395), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1379), .B(n_1347), .Y(n_1413) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1364), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_1375), .A2(n_1361), .B1(n_1357), .B2(n_1322), .Y(n_1415) );
INVx1_ASAP7_75t_SL g1416 ( .A(n_1390), .Y(n_1416) );
OAI21xp33_ASAP7_75t_L g1417 ( .A1(n_1378), .A2(n_1357), .B(n_1338), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1418 ( .A1(n_1402), .A2(n_1383), .B1(n_1364), .B2(n_1380), .Y(n_1418) );
AOI22xp5_ASAP7_75t_L g1419 ( .A1(n_1401), .A2(n_1334), .B1(n_1332), .B2(n_1377), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1414), .B(n_1372), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g1421 ( .A1(n_1415), .A2(n_1370), .B1(n_1385), .B2(n_1369), .C(n_1368), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1399), .Y(n_1422) );
OAI322xp33_ASAP7_75t_L g1423 ( .A1(n_1416), .A2(n_1342), .A3(n_1322), .B1(n_1393), .B2(n_1359), .C1(n_1354), .C2(n_1388), .Y(n_1423) );
AO22x2_ASAP7_75t_L g1424 ( .A1(n_1402), .A2(n_1369), .B1(n_1371), .B2(n_1377), .Y(n_1424) );
OAI221xp5_ASAP7_75t_L g1425 ( .A1(n_1401), .A2(n_1374), .B1(n_1371), .B2(n_1368), .C(n_1342), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_1417), .A2(n_1296), .B1(n_1279), .B2(n_1282), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1427 ( .A1(n_1410), .A2(n_1386), .B1(n_1354), .B2(n_1336), .Y(n_1427) );
AOI221xp5_ASAP7_75t_L g1428 ( .A1(n_1405), .A2(n_1374), .B1(n_1362), .B2(n_1318), .C(n_1349), .Y(n_1428) );
AOI221xp5_ASAP7_75t_SL g1429 ( .A1(n_1398), .A2(n_1363), .B1(n_1329), .B2(n_1325), .C(n_1279), .Y(n_1429) );
NAND2xp5_ASAP7_75t_SL g1430 ( .A(n_1404), .B(n_1384), .Y(n_1430) );
OAI21xp5_ASAP7_75t_L g1431 ( .A1(n_1408), .A2(n_1262), .B(n_1285), .Y(n_1431) );
OAI21xp5_ASAP7_75t_L g1432 ( .A1(n_1404), .A2(n_1285), .B(n_1281), .Y(n_1432) );
OAI21xp33_ASAP7_75t_L g1433 ( .A1(n_1421), .A2(n_1407), .B(n_1406), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1422), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1420), .Y(n_1435) );
NOR3xp33_ASAP7_75t_L g1436 ( .A(n_1418), .B(n_1409), .C(n_1407), .Y(n_1436) );
OAI211xp5_ASAP7_75t_SL g1437 ( .A1(n_1425), .A2(n_1428), .B(n_1419), .C(n_1426), .Y(n_1437) );
AOI322xp5_ASAP7_75t_L g1438 ( .A1(n_1429), .A2(n_1403), .A3(n_1413), .B1(n_1409), .B2(n_1329), .C1(n_1325), .C2(n_1400), .Y(n_1438) );
NOR4xp25_ASAP7_75t_L g1439 ( .A(n_1423), .B(n_1412), .C(n_1397), .D(n_1396), .Y(n_1439) );
CKINVDCx20_ASAP7_75t_R g1440 ( .A(n_1427), .Y(n_1440) );
OAI221xp5_ASAP7_75t_L g1441 ( .A1(n_1432), .A2(n_1411), .B1(n_1281), .B2(n_1366), .C(n_1384), .Y(n_1441) );
OAI221xp5_ASAP7_75t_L g1442 ( .A1(n_1431), .A2(n_1411), .B1(n_1281), .B2(n_1251), .C(n_1226), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_1435), .B(n_1430), .Y(n_1443) );
OAI22xp33_ASAP7_75t_L g1444 ( .A1(n_1440), .A2(n_1424), .B1(n_1281), .B2(n_1226), .Y(n_1444) );
XNOR2xp5_ASAP7_75t_L g1445 ( .A(n_1436), .B(n_1424), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1434), .B(n_1296), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1438), .B(n_1273), .Y(n_1447) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1441), .Y(n_1448) );
NAND3x1_ASAP7_75t_L g1449 ( .A(n_1439), .B(n_1193), .C(n_1226), .Y(n_1449) );
HB1xp67_ASAP7_75t_L g1450 ( .A(n_1443), .Y(n_1450) );
NOR4xp25_ASAP7_75t_L g1451 ( .A(n_1449), .B(n_1433), .C(n_1437), .D(n_1442), .Y(n_1451) );
NOR3xp33_ASAP7_75t_SL g1452 ( .A(n_1445), .B(n_1246), .C(n_1191), .Y(n_1452) );
NOR3xp33_ASAP7_75t_L g1453 ( .A(n_1444), .B(n_1193), .C(n_1132), .Y(n_1453) );
NAND2xp5_ASAP7_75t_SL g1454 ( .A(n_1448), .B(n_1193), .Y(n_1454) );
AOI21x1_ASAP7_75t_L g1455 ( .A1(n_1450), .A2(n_1448), .B(n_1447), .Y(n_1455) );
NAND2xp5_ASAP7_75t_SL g1456 ( .A(n_1451), .B(n_1446), .Y(n_1456) );
INVx2_ASAP7_75t_L g1457 ( .A(n_1454), .Y(n_1457) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1453), .Y(n_1458) );
OAI21x1_ASAP7_75t_L g1459 ( .A1(n_1455), .A2(n_1452), .B(n_1187), .Y(n_1459) );
XNOR2xp5_ASAP7_75t_L g1460 ( .A(n_1456), .B(n_1232), .Y(n_1460) );
XOR2x2_ASAP7_75t_L g1461 ( .A(n_1458), .B(n_1232), .Y(n_1461) );
AOI21xp5_ASAP7_75t_L g1462 ( .A1(n_1460), .A2(n_1457), .B(n_1187), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1461), .Y(n_1463) );
OAI21x1_ASAP7_75t_L g1464 ( .A1(n_1459), .A2(n_1187), .B(n_1239), .Y(n_1464) );
AOI222xp33_ASAP7_75t_SL g1465 ( .A1(n_1463), .A2(n_1461), .B1(n_1256), .B2(n_1216), .C1(n_1249), .C2(n_1190), .Y(n_1465) );
OR2x6_ASAP7_75t_L g1466 ( .A(n_1462), .B(n_1464), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1466), .Y(n_1467) );
AOI21xp5_ASAP7_75t_L g1468 ( .A1(n_1467), .A2(n_1465), .B(n_1190), .Y(n_1468) );
endmodule