module fake_jpeg_26161_n_67 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_13),
.B1(n_23),
.B2(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_37),
.B1(n_29),
.B2(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_2),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_11),
.B1(n_21),
.B2(n_20),
.Y(n_36)
);

A2O1A1O1Ixp25_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_25),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_14),
.B(n_24),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_45),
.B(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_28),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_41),
.C(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_7),
.B(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.C(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.C(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_59),
.B1(n_31),
.B2(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_53),
.B(n_56),
.C(n_58),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_60),
.C(n_17),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_16),
.B(n_19),
.Y(n_67)
);


endmodule