module fake_aes_1203_n_43 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_43);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_10), .B(n_7), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_1), .B(n_8), .Y(n_16) );
INVx6_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_12), .Y(n_22) );
BUFx8_ASAP7_75t_L g23 ( .A(n_11), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_14), .B(n_12), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_19), .A2(n_16), .B1(n_14), .B2(n_15), .C(n_1), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_18), .B(n_0), .Y(n_27) );
NOR4xp25_ASAP7_75t_L g28 ( .A(n_26), .B(n_19), .C(n_20), .D(n_18), .Y(n_28) );
BUFx3_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
BUFx3_ASAP7_75t_L g30 ( .A(n_25), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_24), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_28), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
INVx1_ASAP7_75t_SL g37 ( .A(n_34), .Y(n_37) );
OAI221xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_28), .B1(n_16), .B2(n_23), .C(n_2), .Y(n_38) );
AOI22xp33_ASAP7_75t_R g39 ( .A1(n_36), .A2(n_34), .B1(n_2), .B2(n_0), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_37), .B1(n_36), .B2(n_23), .Y(n_40) );
BUFx2_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_40), .Y(n_42) );
AOI22xp33_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_4), .B1(n_42), .B2(n_40), .Y(n_43) );
endmodule