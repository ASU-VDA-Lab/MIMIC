module fake_jpeg_16063_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_14),
.B1(n_24),
.B2(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_52),
.B1(n_33),
.B2(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_14),
.B1(n_24),
.B2(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_46),
.B1(n_54),
.B2(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_30),
.Y(n_66)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_27),
.B1(n_15),
.B2(n_17),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_66),
.Y(n_76)
);

OR2x4_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_28),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_51),
.B(n_26),
.C(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_48),
.B1(n_38),
.B2(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_52),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_37),
.B1(n_27),
.B2(n_26),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_45),
.B1(n_38),
.B2(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_34),
.B1(n_27),
.B2(n_37),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_69),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_37),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_39),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_74),
.B(n_79),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_13),
.C(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_83),
.B1(n_72),
.B2(n_62),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_96),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_99),
.B1(n_71),
.B2(n_22),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_60),
.C(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_87),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_74),
.A2(n_72),
.B1(n_55),
.B2(n_62),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_83),
.B1(n_86),
.B2(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_126),
.B1(n_92),
.B2(n_120),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_73),
.B1(n_79),
.B2(n_76),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_119),
.B1(n_122),
.B2(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_76),
.B1(n_55),
.B2(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_77),
.B1(n_51),
.B2(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_22),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_99),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_132),
.C(n_119),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_97),
.C(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_134),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_97),
.B(n_95),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_136),
.B(n_117),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_93),
.B(n_105),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_93),
.B1(n_102),
.B2(n_67),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_143),
.Y(n_156)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_142),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_109),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_137),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_160),
.C(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_109),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_122),
.C(n_67),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_167),
.C(n_173),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_130),
.B(n_131),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_158),
.B(n_2),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_134),
.C(n_19),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_153),
.B(n_150),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_170),
.B(n_173),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_148),
.C(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_4),
.B(n_5),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_0),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_166),
.B(n_178),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_194),
.B(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_190),
.A2(n_193),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_192),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_174),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_200),
.C(n_19),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_7),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_162),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_162),
.B(n_7),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_5),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_205),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_196),
.C(n_19),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_200),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_211),
.A3(n_207),
.B1(n_208),
.B2(n_206),
.C1(n_11),
.C2(n_12),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_18),
.C(n_9),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_207),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_8),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_10),
.Y(n_216)
);


endmodule