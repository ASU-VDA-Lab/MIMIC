module fake_ariane_3351_n_6182 (n_913, n_1681, n_1486, n_1507, n_589, n_1174, n_1469, n_691, n_1353, n_1355, n_423, n_1383, n_603, n_373, n_1250, n_1169, n_789, n_850, n_610, n_245, n_1713, n_96, n_319, n_49, n_1436, n_690, n_416, n_1109, n_1430, n_525, n_187, n_1463, n_1238, n_1515, n_817, n_924, n_781, n_1566, n_189, n_717, n_72, n_952, n_864, n_1096, n_1379, n_57, n_1706, n_117, n_524, n_1214, n_634, n_1246, n_1138, n_214, n_764, n_1503, n_462, n_1196, n_1181, n_32, n_410, n_1187, n_1131, n_1225, n_737, n_137, n_1298, n_1366, n_232, n_52, n_568, n_1088, n_77, n_1424, n_766, n_1457, n_377, n_1682, n_520, n_870, n_1453, n_279, n_945, n_958, n_813, n_419, n_146, n_270, n_338, n_995, n_285, n_1184, n_202, n_1535, n_500, n_665, n_754, n_903, n_871, n_1073, n_239, n_402, n_1277, n_54, n_829, n_1062, n_339, n_738, n_1690, n_672, n_740, n_1283, n_167, n_1018, n_69, n_259, n_953, n_1364, n_143, n_1224, n_1425, n_625, n_557, n_1107, n_1688, n_989, n_242, n_645, n_331, n_559, n_267, n_495, n_350, n_381, n_795, n_721, n_1084, n_1276, n_200, n_1428, n_1284, n_1241, n_821, n_561, n_770, n_1514, n_1528, n_507, n_486, n_901, n_569, n_1145, n_971, n_787, n_1650, n_31, n_1519, n_1195, n_1522, n_518, n_1207, n_222, n_786, n_1404, n_868, n_1542, n_1314, n_1512, n_1539, n_884, n_1415, n_1034, n_1652, n_1676, n_1085, n_277, n_1636, n_432, n_293, n_823, n_620, n_93, n_1074, n_859, n_108, n_587, n_693, n_863, n_303, n_1254, n_929, n_206, n_352, n_899, n_1703, n_611, n_1295, n_238, n_365, n_1013, n_1495, n_1637, n_136, n_334, n_192, n_661, n_300, n_533, n_104, n_438, n_1560, n_1654, n_1548, n_16, n_440, n_273, n_1396, n_1230, n_612, n_333, n_376, n_512, n_1597, n_1544, n_579, n_844, n_1012, n_1267, n_1354, n_149, n_1213, n_237, n_780, n_1021, n_1443, n_491, n_1465, n_1595, n_1142, n_1140, n_705, n_570, n_260, n_942, n_1437, n_7, n_1378, n_461, n_1121, n_1416, n_209, n_490, n_1461, n_17, n_1391, n_225, n_1599, n_1006, n_575, n_546, n_503, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_1669, n_1675, n_676, n_42, n_1594, n_680, n_287, n_1716, n_302, n_380, n_1585, n_1432, n_94, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_1590, n_1351, n_1274, n_257, n_652, n_475, n_135, n_947, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_1442, n_482, n_798, n_577, n_407, n_1691, n_27, n_916, n_1386, n_912, n_460, n_1555, n_366, n_762, n_1253, n_1468, n_1661, n_555, n_804, n_1656, n_1382, n_966, n_992, n_955, n_1182, n_794, n_78, n_1692, n_1562, n_514, n_418, n_1376, n_513, n_288, n_179, n_1292, n_1178, n_1435, n_1026, n_1506, n_1610, n_306, n_92, n_203, n_436, n_150, n_324, n_669, n_931, n_1491, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_1418, n_746, n_1357, n_292, n_1079, n_1389, n_615, n_1139, n_76, n_517, n_1312, n_1717, n_0, n_824, n_428, n_159, n_892, n_959, n_30, n_1399, n_1101, n_1567, n_1343, n_563, n_144, n_990, n_1623, n_867, n_1226, n_944, n_749, n_815, n_542, n_1340, n_470, n_1240, n_1087, n_632, n_477, n_650, n_425, n_1433, n_1155, n_1071, n_712, n_976, n_909, n_1392, n_767, n_1680, n_964, n_1627, n_382, n_489, n_80, n_251, n_974, n_506, n_799, n_1147, n_397, n_471, n_351, n_965, n_155, n_934, n_1447, n_1220, n_356, n_698, n_1674, n_124, n_307, n_1209, n_1020, n_1563, n_646, n_1633, n_34, n_404, n_172, n_1058, n_347, n_1042, n_183, n_1234, n_479, n_1578, n_1455, n_299, n_836, n_1279, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_1568, n_20, n_1483, n_1363, n_367, n_1111, n_970, n_1689, n_713, n_1255, n_1646, n_598, n_345, n_1237, n_927, n_261, n_1095, n_370, n_706, n_286, n_1401, n_1419, n_1531, n_776, n_424, n_1651, n_85, n_130, n_1387, n_466, n_1263, n_346, n_348, n_552, n_670, n_379, n_138, n_162, n_264, n_441, n_1032, n_1217, n_1496, n_637, n_1592, n_73, n_327, n_1259, n_1177, n_1231, n_980, n_1618, n_905, n_207, n_720, n_926, n_41, n_194, n_1163, n_186, n_1384, n_145, n_59, n_1501, n_1173, n_1068, n_1198, n_1570, n_487, n_1518, n_1456, n_90, n_1648, n_1413, n_855, n_158, n_808, n_1365, n_553, n_1439, n_814, n_578, n_1665, n_1287, n_405, n_1611, n_120, n_320, n_1414, n_1134, n_1484, n_647, n_1423, n_481, n_600, n_1053, n_1609, n_529, n_502, n_218, n_1467, n_247, n_1304, n_1608, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1349, n_1709, n_1061, n_326, n_681, n_227, n_874, n_1278, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_545, n_1015, n_1377, n_1162, n_536, n_1614, n_325, n_1602, n_688, n_636, n_427, n_1098, n_1490, n_442, n_777, n_1553, n_1080, n_920, n_1086, n_1092, n_986, n_1104, n_729, n_887, n_1122, n_1205, n_1408, n_163, n_1693, n_1132, n_390, n_1156, n_501, n_314, n_1120, n_1202, n_627, n_1188, n_1498, n_1371, n_233, n_957, n_388, n_1402, n_1242, n_1607, n_1489, n_1218, n_221, n_321, n_86, n_1586, n_861, n_1543, n_1431, n_877, n_1119, n_1666, n_1500, n_616, n_1055, n_1395, n_1346, n_1189, n_1089, n_281, n_262, n_1502, n_1523, n_1478, n_735, n_297, n_1005, n_527, n_46, n_84, n_1294, n_1667, n_845, n_888, n_1649, n_1677, n_1297, n_178, n_551, n_417, n_1708, n_70, n_343, n_1222, n_582, n_755, n_1097, n_1219, n_1711, n_710, n_534, n_1460, n_1239, n_278, n_560, n_890, n_842, n_148, n_451, n_745, n_1572, n_61, n_742, n_1081, n_1373, n_1388, n_1266, n_1540, n_769, n_13, n_1372, n_476, n_832, n_55, n_535, n_744, n_982, n_915, n_215, n_1075, n_454, n_298, n_1331, n_1529, n_1227, n_655, n_403, n_1007, n_1580, n_1319, n_657, n_837, n_812, n_606, n_951, n_862, n_1700, n_659, n_1332, n_509, n_666, n_430, n_1206, n_722, n_1508, n_1532, n_1171, n_1030, n_785, n_1309, n_999, n_1338, n_1342, n_456, n_852, n_1394, n_704, n_1060, n_1044, n_1714, n_521, n_873, n_1301, n_1243, n_1400, n_342, n_1466, n_1513, n_1527, n_358, n_608, n_1538, n_1037, n_1329, n_317, n_1545, n_134, n_1257, n_1480, n_1668, n_1605, n_1078, n_266, n_157, n_1161, n_811, n_624, n_791, n_876, n_618, n_1191, n_736, n_1025, n_1215, n_241, n_1449, n_687, n_797, n_480, n_1327, n_1475, n_211, n_642, n_97, n_408, n_1406, n_595, n_1405, n_602, n_592, n_1499, n_854, n_1318, n_393, n_1632, n_474, n_805, n_295, n_1658, n_190, n_1072, n_695, n_1526, n_1305, n_64, n_180, n_730, n_386, n_1596, n_1281, n_516, n_1137, n_1258, n_197, n_640, n_463, n_1476, n_1524, n_943, n_1118, n_678, n_651, n_1293, n_961, n_469, n_1046, n_726, n_1123, n_1657, n_878, n_771, n_1321, n_752, n_71, n_1488, n_985, n_421, n_1330, n_906, n_1180, n_1697, n_283, n_806, n_1350, n_1556, n_649, n_1561, n_374, n_1352, n_643, n_1492, n_226, n_1441, n_682, n_36, n_1616, n_819, n_586, n_1324, n_1429, n_686, n_605, n_1154, n_584, n_1557, n_1130, n_1450, n_349, n_756, n_1016, n_1149, n_1505, n_979, n_1642, n_2, n_897, n_949, n_1493, n_515, n_807, n_891, n_885, n_1659, n_198, n_1208, n_396, n_802, n_23, n_1151, n_554, n_960, n_1256, n_87, n_714, n_790, n_354, n_140, n_725, n_1577, n_151, n_1448, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_801, n_1286, n_818, n_1685, n_779, n_594, n_1397, n_35, n_1052, n_272, n_1333, n_1306, n_833, n_1426, n_879, n_1117, n_38, n_422, n_1269, n_1303, n_1547, n_1438, n_1541, n_597, n_75, n_1047, n_95, n_1472, n_1593, n_1050, n_566, n_152, n_169, n_106, n_1201, n_1288, n_173, n_858, n_1185, n_335, n_1035, n_1143, n_344, n_426, n_433, n_398, n_62, n_210, n_1090, n_1367, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1565, n_1192, n_128, n_224, n_82, n_894, n_1380, n_1624, n_420, n_1291, n_562, n_748, n_510, n_1045, n_256, n_1160, n_1023, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_467, n_1511, n_1422, n_644, n_1197, n_276, n_497, n_1165, n_1641, n_168, n_81, n_538, n_1517, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_1307, n_1128, n_1671, n_1417, n_1048, n_775, n_667, n_1049, n_14, n_869, n_141, n_846, n_1398, n_1356, n_1341, n_1504, n_1440, n_1370, n_1603, n_305, n_312, n_56, n_60, n_728, n_413, n_715, n_889, n_1066, n_1549, n_935, n_685, n_911, n_361, n_89, n_623, n_1712, n_1403, n_1065, n_453, n_1534, n_74, n_810, n_19, n_40, n_1290, n_181, n_617, n_543, n_1362, n_1559, n_236, n_601, n_683, n_565, n_628, n_1300, n_743, n_1194, n_1647, n_1546, n_1420, n_907, n_1454, n_660, n_464, n_962, n_941, n_1210, n_847, n_747, n_1622, n_1135, n_918, n_107, n_639, n_452, n_673, n_1038, n_414, n_571, n_1521, n_1694, n_6, n_284, n_593, n_1695, n_1164, n_37, n_58, n_609, n_1193, n_1345, n_613, n_1022, n_1336, n_1033, n_409, n_171, n_519, n_384, n_1166, n_1056, n_526, n_1040, n_674, n_1158, n_316, n_125, n_1444, n_820, n_43, n_872, n_1653, n_254, n_1157, n_1584, n_234, n_848, n_1664, n_280, n_629, n_161, n_532, n_763, n_99, n_540, n_216, n_692, n_5, n_984, n_1687, n_223, n_1552, n_750, n_834, n_1612, n_800, n_1606, n_395, n_621, n_1587, n_213, n_67, n_1014, n_724, n_1427, n_1481, n_493, n_1311, n_1589, n_114, n_1100, n_585, n_875, n_1617, n_827, n_697, n_622, n_1626, n_1335, n_1715, n_296, n_880, n_793, n_1175, n_132, n_751, n_1027, n_1070, n_1621, n_739, n_1485, n_1028, n_1221, n_530, n_792, n_1262, n_580, n_1579, n_494, n_434, n_975, n_229, n_394, n_923, n_1645, n_1124, n_1381, n_1494, n_932, n_1183, n_1326, n_981, n_1110, n_243, n_1407, n_185, n_1204, n_1554, n_994, n_1360, n_973, n_268, n_972, n_164, n_184, n_856, n_1248, n_1176, n_1564, n_1054, n_508, n_118, n_121, n_1679, n_353, n_1678, n_1482, n_1361, n_1601, n_1057, n_191, n_978, n_1011, n_1520, n_1509, n_828, n_322, n_1411, n_1359, n_558, n_116, n_39, n_653, n_1445, n_1317, n_783, n_556, n_1127, n_170, n_1536, n_1471, n_160, n_119, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_987, n_936, n_1620, n_1385, n_1525, n_541, n_499, n_788, n_12, n_908, n_1036, n_341, n_1270, n_109, n_1167, n_1272, n_549, n_591, n_969, n_919, n_1663, n_50, n_1625, n_318, n_1458, n_103, n_244, n_679, n_1630, n_220, n_663, n_443, n_1412, n_1550, n_528, n_1358, n_1200, n_387, n_406, n_826, n_139, n_391, n_940, n_1537, n_1077, n_607, n_956, n_445, n_765, n_122, n_1268, n_385, n_917, n_1271, n_372, n_15, n_1530, n_631, n_399, n_1170, n_1261, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1323, n_1462, n_1064, n_633, n_900, n_1446, n_1282, n_1701, n_1093, n_1551, n_1285, n_193, n_733, n_761, n_731, n_336, n_315, n_311, n_1452, n_1573, n_8, n_668, n_758, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_1322, n_1473, n_835, n_446, n_1076, n_1348, n_753, n_701, n_1003, n_1125, n_1710, n_309, n_1344, n_115, n_1390, n_401, n_485, n_504, n_483, n_435, n_1141, n_1629, n_291, n_1640, n_822, n_1094, n_840, n_1459, n_1510, n_1099, n_839, n_79, n_3, n_759, n_567, n_91, n_240, n_369, n_44, n_1575, n_1172, n_614, n_1212, n_831, n_778, n_48, n_1619, n_188, n_323, n_550, n_1315, n_1660, n_997, n_635, n_694, n_1643, n_1320, n_1113, n_248, n_1152, n_921, n_1615, n_1236, n_228, n_1265, n_1576, n_1470, n_671, n_1533, n_1, n_1409, n_1148, n_1588, n_1684, n_1673, n_1334, n_654, n_1275, n_488, n_904, n_505, n_88, n_1696, n_498, n_1059, n_684, n_1039, n_539, n_1150, n_977, n_449, n_392, n_1628, n_1289, n_1497, n_459, n_1136, n_458, n_1190, n_1600, n_1144, n_383, n_838, n_1558, n_1316, n_175, n_950, n_1017, n_711, n_734, n_723, n_1393, n_658, n_630, n_1369, n_53, n_362, n_310, n_709, n_24, n_809, n_1686, n_235, n_881, n_1019, n_1477, n_662, n_641, n_910, n_290, n_741, n_939, n_1410, n_371, n_199, n_217, n_1114, n_1325, n_708, n_308, n_1223, n_201, n_572, n_1199, n_865, n_10, n_1273, n_1041, n_993, n_948, n_922, n_1004, n_448, n_1347, n_860, n_1043, n_255, n_450, n_896, n_1479, n_1613, n_902, n_1031, n_1638, n_853, n_716, n_1571, n_1698, n_196, n_1337, n_774, n_933, n_596, n_954, n_1168, n_219, n_1310, n_231, n_656, n_492, n_574, n_252, n_664, n_1591, n_1229, n_1683, n_68, n_415, n_63, n_1280, n_544, n_1516, n_1186, n_1705, n_599, n_768, n_1091, n_537, n_1063, n_25, n_991, n_83, n_389, n_1670, n_1707, n_1126, n_195, n_938, n_1328, n_895, n_110, n_304, n_1639, n_583, n_1302, n_1000, n_313, n_626, n_378, n_1581, n_98, n_946, n_757, n_375, n_113, n_1655, n_33, n_1146, n_1634, n_1203, n_998, n_1699, n_1598, n_472, n_937, n_1474, n_265, n_1583, n_1604, n_208, n_1631, n_1702, n_156, n_174, n_275, n_100, n_1375, n_147, n_204, n_1232, n_996, n_1211, n_1368, n_963, n_1264, n_51, n_1082, n_496, n_866, n_26, n_246, n_925, n_1313, n_1001, n_1115, n_1339, n_1002, n_1644, n_105, n_1051, n_719, n_131, n_263, n_1102, n_360, n_1129, n_1252, n_250, n_1464, n_1296, n_773, n_165, n_1010, n_882, n_1249, n_101, n_803, n_329, n_718, n_1434, n_340, n_1569, n_289, n_9, n_112, n_45, n_548, n_523, n_1662, n_457, n_1299, n_177, n_782, n_364, n_258, n_431, n_1228, n_1244, n_411, n_484, n_849, n_22, n_29, n_357, n_412, n_1251, n_447, n_1421, n_1233, n_1574, n_1672, n_1635, n_1704, n_893, n_1582, n_841, n_886, n_1069, n_359, n_1308, n_573, n_796, n_127, n_531, n_1374, n_1451, n_1487, n_675, n_6182);

input n_913;
input n_1681;
input n_1486;
input n_1507;
input n_589;
input n_1174;
input n_1469;
input n_691;
input n_1353;
input n_1355;
input n_423;
input n_1383;
input n_603;
input n_373;
input n_1250;
input n_1169;
input n_789;
input n_850;
input n_610;
input n_245;
input n_1713;
input n_96;
input n_319;
input n_49;
input n_1436;
input n_690;
input n_416;
input n_1109;
input n_1430;
input n_525;
input n_187;
input n_1463;
input n_1238;
input n_1515;
input n_817;
input n_924;
input n_781;
input n_1566;
input n_189;
input n_717;
input n_72;
input n_952;
input n_864;
input n_1096;
input n_1379;
input n_57;
input n_1706;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1246;
input n_1138;
input n_214;
input n_764;
input n_1503;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_410;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_1298;
input n_1366;
input n_232;
input n_52;
input n_568;
input n_1088;
input n_77;
input n_1424;
input n_766;
input n_1457;
input n_377;
input n_1682;
input n_520;
input n_870;
input n_1453;
input n_279;
input n_945;
input n_958;
input n_813;
input n_419;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1184;
input n_202;
input n_1535;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_1073;
input n_239;
input n_402;
input n_1277;
input n_54;
input n_829;
input n_1062;
input n_339;
input n_738;
input n_1690;
input n_672;
input n_740;
input n_1283;
input n_167;
input n_1018;
input n_69;
input n_259;
input n_953;
input n_1364;
input n_143;
input n_1224;
input n_1425;
input n_625;
input n_557;
input n_1107;
input n_1688;
input n_989;
input n_242;
input n_645;
input n_331;
input n_559;
input n_267;
input n_495;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_1276;
input n_200;
input n_1428;
input n_1284;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_1514;
input n_1528;
input n_507;
input n_486;
input n_901;
input n_569;
input n_1145;
input n_971;
input n_787;
input n_1650;
input n_31;
input n_1519;
input n_1195;
input n_1522;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_1404;
input n_868;
input n_1542;
input n_1314;
input n_1512;
input n_1539;
input n_884;
input n_1415;
input n_1034;
input n_1652;
input n_1676;
input n_1085;
input n_277;
input n_1636;
input n_432;
input n_293;
input n_823;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_108;
input n_587;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_206;
input n_352;
input n_899;
input n_1703;
input n_611;
input n_1295;
input n_238;
input n_365;
input n_1013;
input n_1495;
input n_1637;
input n_136;
input n_334;
input n_192;
input n_661;
input n_300;
input n_533;
input n_104;
input n_438;
input n_1560;
input n_1654;
input n_1548;
input n_16;
input n_440;
input n_273;
input n_1396;
input n_1230;
input n_612;
input n_333;
input n_376;
input n_512;
input n_1597;
input n_1544;
input n_579;
input n_844;
input n_1012;
input n_1267;
input n_1354;
input n_149;
input n_1213;
input n_237;
input n_780;
input n_1021;
input n_1443;
input n_491;
input n_1465;
input n_1595;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_1437;
input n_7;
input n_1378;
input n_461;
input n_1121;
input n_1416;
input n_209;
input n_490;
input n_1461;
input n_17;
input n_1391;
input n_225;
input n_1599;
input n_1006;
input n_575;
input n_546;
input n_503;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_1669;
input n_1675;
input n_676;
input n_42;
input n_1594;
input n_680;
input n_287;
input n_1716;
input n_302;
input n_380;
input n_1585;
input n_1432;
input n_94;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_1590;
input n_1351;
input n_1274;
input n_257;
input n_652;
input n_475;
input n_135;
input n_947;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_1442;
input n_482;
input n_798;
input n_577;
input n_407;
input n_1691;
input n_27;
input n_916;
input n_1386;
input n_912;
input n_460;
input n_1555;
input n_366;
input n_762;
input n_1253;
input n_1468;
input n_1661;
input n_555;
input n_804;
input n_1656;
input n_1382;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_1692;
input n_1562;
input n_514;
input n_418;
input n_1376;
input n_513;
input n_288;
input n_179;
input n_1292;
input n_1178;
input n_1435;
input n_1026;
input n_1506;
input n_1610;
input n_306;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_669;
input n_931;
input n_1491;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_1418;
input n_746;
input n_1357;
input n_292;
input n_1079;
input n_1389;
input n_615;
input n_1139;
input n_76;
input n_517;
input n_1312;
input n_1717;
input n_0;
input n_824;
input n_428;
input n_159;
input n_892;
input n_959;
input n_30;
input n_1399;
input n_1101;
input n_1567;
input n_1343;
input n_563;
input n_144;
input n_990;
input n_1623;
input n_867;
input n_1226;
input n_944;
input n_749;
input n_815;
input n_542;
input n_1340;
input n_470;
input n_1240;
input n_1087;
input n_632;
input n_477;
input n_650;
input n_425;
input n_1433;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_1392;
input n_767;
input n_1680;
input n_964;
input n_1627;
input n_382;
input n_489;
input n_80;
input n_251;
input n_974;
input n_506;
input n_799;
input n_1147;
input n_397;
input n_471;
input n_351;
input n_965;
input n_155;
input n_934;
input n_1447;
input n_1220;
input n_356;
input n_698;
input n_1674;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_1563;
input n_646;
input n_1633;
input n_34;
input n_404;
input n_172;
input n_1058;
input n_347;
input n_1042;
input n_183;
input n_1234;
input n_479;
input n_1578;
input n_1455;
input n_299;
input n_836;
input n_1279;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_1568;
input n_20;
input n_1483;
input n_1363;
input n_367;
input n_1111;
input n_970;
input n_1689;
input n_713;
input n_1255;
input n_1646;
input n_598;
input n_345;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_370;
input n_706;
input n_286;
input n_1401;
input n_1419;
input n_1531;
input n_776;
input n_424;
input n_1651;
input n_85;
input n_130;
input n_1387;
input n_466;
input n_1263;
input n_346;
input n_348;
input n_552;
input n_670;
input n_379;
input n_138;
input n_162;
input n_264;
input n_441;
input n_1032;
input n_1217;
input n_1496;
input n_637;
input n_1592;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_980;
input n_1618;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_194;
input n_1163;
input n_186;
input n_1384;
input n_145;
input n_59;
input n_1501;
input n_1173;
input n_1068;
input n_1198;
input n_1570;
input n_487;
input n_1518;
input n_1456;
input n_90;
input n_1648;
input n_1413;
input n_855;
input n_158;
input n_808;
input n_1365;
input n_553;
input n_1439;
input n_814;
input n_578;
input n_1665;
input n_1287;
input n_405;
input n_1611;
input n_120;
input n_320;
input n_1414;
input n_1134;
input n_1484;
input n_647;
input n_1423;
input n_481;
input n_600;
input n_1053;
input n_1609;
input n_529;
input n_502;
input n_218;
input n_1467;
input n_247;
input n_1304;
input n_1608;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1349;
input n_1709;
input n_1061;
input n_326;
input n_681;
input n_227;
input n_874;
input n_1278;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_545;
input n_1015;
input n_1377;
input n_1162;
input n_536;
input n_1614;
input n_325;
input n_1602;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_1490;
input n_442;
input n_777;
input n_1553;
input n_1080;
input n_920;
input n_1086;
input n_1092;
input n_986;
input n_1104;
input n_729;
input n_887;
input n_1122;
input n_1205;
input n_1408;
input n_163;
input n_1693;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_314;
input n_1120;
input n_1202;
input n_627;
input n_1188;
input n_1498;
input n_1371;
input n_233;
input n_957;
input n_388;
input n_1402;
input n_1242;
input n_1607;
input n_1489;
input n_1218;
input n_221;
input n_321;
input n_86;
input n_1586;
input n_861;
input n_1543;
input n_1431;
input n_877;
input n_1119;
input n_1666;
input n_1500;
input n_616;
input n_1055;
input n_1395;
input n_1346;
input n_1189;
input n_1089;
input n_281;
input n_262;
input n_1502;
input n_1523;
input n_1478;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_46;
input n_84;
input n_1294;
input n_1667;
input n_845;
input n_888;
input n_1649;
input n_1677;
input n_1297;
input n_178;
input n_551;
input n_417;
input n_1708;
input n_70;
input n_343;
input n_1222;
input n_582;
input n_755;
input n_1097;
input n_1219;
input n_1711;
input n_710;
input n_534;
input n_1460;
input n_1239;
input n_278;
input n_560;
input n_890;
input n_842;
input n_148;
input n_451;
input n_745;
input n_1572;
input n_61;
input n_742;
input n_1081;
input n_1373;
input n_1388;
input n_1266;
input n_1540;
input n_769;
input n_13;
input n_1372;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_982;
input n_915;
input n_215;
input n_1075;
input n_454;
input n_298;
input n_1331;
input n_1529;
input n_1227;
input n_655;
input n_403;
input n_1007;
input n_1580;
input n_1319;
input n_657;
input n_837;
input n_812;
input n_606;
input n_951;
input n_862;
input n_1700;
input n_659;
input n_1332;
input n_509;
input n_666;
input n_430;
input n_1206;
input n_722;
input n_1508;
input n_1532;
input n_1171;
input n_1030;
input n_785;
input n_1309;
input n_999;
input n_1338;
input n_1342;
input n_456;
input n_852;
input n_1394;
input n_704;
input n_1060;
input n_1044;
input n_1714;
input n_521;
input n_873;
input n_1301;
input n_1243;
input n_1400;
input n_342;
input n_1466;
input n_1513;
input n_1527;
input n_358;
input n_608;
input n_1538;
input n_1037;
input n_1329;
input n_317;
input n_1545;
input n_134;
input n_1257;
input n_1480;
input n_1668;
input n_1605;
input n_1078;
input n_266;
input n_157;
input n_1161;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_1449;
input n_687;
input n_797;
input n_480;
input n_1327;
input n_1475;
input n_211;
input n_642;
input n_97;
input n_408;
input n_1406;
input n_595;
input n_1405;
input n_602;
input n_592;
input n_1499;
input n_854;
input n_1318;
input n_393;
input n_1632;
input n_474;
input n_805;
input n_295;
input n_1658;
input n_190;
input n_1072;
input n_695;
input n_1526;
input n_1305;
input n_64;
input n_180;
input n_730;
input n_386;
input n_1596;
input n_1281;
input n_516;
input n_1137;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_1476;
input n_1524;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_1293;
input n_961;
input n_469;
input n_1046;
input n_726;
input n_1123;
input n_1657;
input n_878;
input n_771;
input n_1321;
input n_752;
input n_71;
input n_1488;
input n_985;
input n_421;
input n_1330;
input n_906;
input n_1180;
input n_1697;
input n_283;
input n_806;
input n_1350;
input n_1556;
input n_649;
input n_1561;
input n_374;
input n_1352;
input n_643;
input n_1492;
input n_226;
input n_1441;
input n_682;
input n_36;
input n_1616;
input n_819;
input n_586;
input n_1324;
input n_1429;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1557;
input n_1130;
input n_1450;
input n_349;
input n_756;
input n_1016;
input n_1149;
input n_1505;
input n_979;
input n_1642;
input n_2;
input n_897;
input n_949;
input n_1493;
input n_515;
input n_807;
input n_891;
input n_885;
input n_1659;
input n_198;
input n_1208;
input n_396;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_1256;
input n_87;
input n_714;
input n_790;
input n_354;
input n_140;
input n_725;
input n_1577;
input n_151;
input n_1448;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_801;
input n_1286;
input n_818;
input n_1685;
input n_779;
input n_594;
input n_1397;
input n_35;
input n_1052;
input n_272;
input n_1333;
input n_1306;
input n_833;
input n_1426;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_1269;
input n_1303;
input n_1547;
input n_1438;
input n_1541;
input n_597;
input n_75;
input n_1047;
input n_95;
input n_1472;
input n_1593;
input n_1050;
input n_566;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_1288;
input n_173;
input n_858;
input n_1185;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_1367;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1565;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_1380;
input n_1624;
input n_420;
input n_1291;
input n_562;
input n_748;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1023;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_467;
input n_1511;
input n_1422;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_1641;
input n_168;
input n_81;
input n_538;
input n_1517;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_1307;
input n_1128;
input n_1671;
input n_1417;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_14;
input n_869;
input n_141;
input n_846;
input n_1398;
input n_1356;
input n_1341;
input n_1504;
input n_1440;
input n_1370;
input n_1603;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_715;
input n_889;
input n_1066;
input n_1549;
input n_935;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1712;
input n_1403;
input n_1065;
input n_453;
input n_1534;
input n_74;
input n_810;
input n_19;
input n_40;
input n_1290;
input n_181;
input n_617;
input n_543;
input n_1362;
input n_1559;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_1300;
input n_743;
input n_1194;
input n_1647;
input n_1546;
input n_1420;
input n_907;
input n_1454;
input n_660;
input n_464;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1622;
input n_1135;
input n_918;
input n_107;
input n_639;
input n_452;
input n_673;
input n_1038;
input n_414;
input n_571;
input n_1521;
input n_1694;
input n_6;
input n_284;
input n_593;
input n_1695;
input n_1164;
input n_37;
input n_58;
input n_609;
input n_1193;
input n_1345;
input n_613;
input n_1022;
input n_1336;
input n_1033;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_526;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_1444;
input n_820;
input n_43;
input n_872;
input n_1653;
input n_254;
input n_1157;
input n_1584;
input n_234;
input n_848;
input n_1664;
input n_280;
input n_629;
input n_161;
input n_532;
input n_763;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_984;
input n_1687;
input n_223;
input n_1552;
input n_750;
input n_834;
input n_1612;
input n_800;
input n_1606;
input n_395;
input n_621;
input n_1587;
input n_213;
input n_67;
input n_1014;
input n_724;
input n_1427;
input n_1481;
input n_493;
input n_1311;
input n_1589;
input n_114;
input n_1100;
input n_585;
input n_875;
input n_1617;
input n_827;
input n_697;
input n_622;
input n_1626;
input n_1335;
input n_1715;
input n_296;
input n_880;
input n_793;
input n_1175;
input n_132;
input n_751;
input n_1027;
input n_1070;
input n_1621;
input n_739;
input n_1485;
input n_1028;
input n_1221;
input n_530;
input n_792;
input n_1262;
input n_580;
input n_1579;
input n_494;
input n_434;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1645;
input n_1124;
input n_1381;
input n_1494;
input n_932;
input n_1183;
input n_1326;
input n_981;
input n_1110;
input n_243;
input n_1407;
input n_185;
input n_1204;
input n_1554;
input n_994;
input n_1360;
input n_973;
input n_268;
input n_972;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1564;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_1679;
input n_353;
input n_1678;
input n_1482;
input n_1361;
input n_1601;
input n_1057;
input n_191;
input n_978;
input n_1011;
input n_1520;
input n_1509;
input n_828;
input n_322;
input n_1411;
input n_1359;
input n_558;
input n_116;
input n_39;
input n_653;
input n_1445;
input n_1317;
input n_783;
input n_556;
input n_1127;
input n_170;
input n_1536;
input n_1471;
input n_160;
input n_119;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_987;
input n_936;
input n_1620;
input n_1385;
input n_1525;
input n_541;
input n_499;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_341;
input n_1270;
input n_109;
input n_1167;
input n_1272;
input n_549;
input n_591;
input n_969;
input n_919;
input n_1663;
input n_50;
input n_1625;
input n_318;
input n_1458;
input n_103;
input n_244;
input n_679;
input n_1630;
input n_220;
input n_663;
input n_443;
input n_1412;
input n_1550;
input n_528;
input n_1358;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_391;
input n_940;
input n_1537;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_765;
input n_122;
input n_1268;
input n_385;
input n_917;
input n_1271;
input n_372;
input n_15;
input n_1530;
input n_631;
input n_399;
input n_1170;
input n_1261;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1323;
input n_1462;
input n_1064;
input n_633;
input n_900;
input n_1446;
input n_1282;
input n_1701;
input n_1093;
input n_1551;
input n_1285;
input n_193;
input n_733;
input n_761;
input n_731;
input n_336;
input n_315;
input n_311;
input n_1452;
input n_1573;
input n_8;
input n_668;
input n_758;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_1322;
input n_1473;
input n_835;
input n_446;
input n_1076;
input n_1348;
input n_753;
input n_701;
input n_1003;
input n_1125;
input n_1710;
input n_309;
input n_1344;
input n_115;
input n_1390;
input n_401;
input n_485;
input n_504;
input n_483;
input n_435;
input n_1141;
input n_1629;
input n_291;
input n_1640;
input n_822;
input n_1094;
input n_840;
input n_1459;
input n_1510;
input n_1099;
input n_839;
input n_79;
input n_3;
input n_759;
input n_567;
input n_91;
input n_240;
input n_369;
input n_44;
input n_1575;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_1619;
input n_188;
input n_323;
input n_550;
input n_1315;
input n_1660;
input n_997;
input n_635;
input n_694;
input n_1643;
input n_1320;
input n_1113;
input n_248;
input n_1152;
input n_921;
input n_1615;
input n_1236;
input n_228;
input n_1265;
input n_1576;
input n_1470;
input n_671;
input n_1533;
input n_1;
input n_1409;
input n_1148;
input n_1588;
input n_1684;
input n_1673;
input n_1334;
input n_654;
input n_1275;
input n_488;
input n_904;
input n_505;
input n_88;
input n_1696;
input n_498;
input n_1059;
input n_684;
input n_1039;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_392;
input n_1628;
input n_1289;
input n_1497;
input n_459;
input n_1136;
input n_458;
input n_1190;
input n_1600;
input n_1144;
input n_383;
input n_838;
input n_1558;
input n_1316;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_723;
input n_1393;
input n_658;
input n_630;
input n_1369;
input n_53;
input n_362;
input n_310;
input n_709;
input n_24;
input n_809;
input n_1686;
input n_235;
input n_881;
input n_1019;
input n_1477;
input n_662;
input n_641;
input n_910;
input n_290;
input n_741;
input n_939;
input n_1410;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_1325;
input n_708;
input n_308;
input n_1223;
input n_201;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1273;
input n_1041;
input n_993;
input n_948;
input n_922;
input n_1004;
input n_448;
input n_1347;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_896;
input n_1479;
input n_1613;
input n_902;
input n_1031;
input n_1638;
input n_853;
input n_716;
input n_1571;
input n_1698;
input n_196;
input n_1337;
input n_774;
input n_933;
input n_596;
input n_954;
input n_1168;
input n_219;
input n_1310;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1591;
input n_1229;
input n_1683;
input n_68;
input n_415;
input n_63;
input n_1280;
input n_544;
input n_1516;
input n_1186;
input n_1705;
input n_599;
input n_768;
input n_1091;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_83;
input n_389;
input n_1670;
input n_1707;
input n_1126;
input n_195;
input n_938;
input n_1328;
input n_895;
input n_110;
input n_304;
input n_1639;
input n_583;
input n_1302;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_1581;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_1655;
input n_33;
input n_1146;
input n_1634;
input n_1203;
input n_998;
input n_1699;
input n_1598;
input n_472;
input n_937;
input n_1474;
input n_265;
input n_1583;
input n_1604;
input n_208;
input n_1631;
input n_1702;
input n_156;
input n_174;
input n_275;
input n_100;
input n_1375;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_1368;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_496;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1313;
input n_1001;
input n_1115;
input n_1339;
input n_1002;
input n_1644;
input n_105;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_1129;
input n_1252;
input n_250;
input n_1464;
input n_1296;
input n_773;
input n_165;
input n_1010;
input n_882;
input n_1249;
input n_101;
input n_803;
input n_329;
input n_718;
input n_1434;
input n_340;
input n_1569;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_523;
input n_1662;
input n_457;
input n_1299;
input n_177;
input n_782;
input n_364;
input n_258;
input n_431;
input n_1228;
input n_1244;
input n_411;
input n_484;
input n_849;
input n_22;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_447;
input n_1421;
input n_1233;
input n_1574;
input n_1672;
input n_1635;
input n_1704;
input n_893;
input n_1582;
input n_841;
input n_886;
input n_1069;
input n_359;
input n_1308;
input n_573;
input n_796;
input n_127;
input n_531;
input n_1374;
input n_1451;
input n_1487;
input n_675;

output n_6182;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_2680;
wire n_3264;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_2002;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_5302;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_5712;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_5479;
wire n_2646;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_2482;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_2807;
wire n_4512;
wire n_4132;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_4741;
wire n_4143;
wire n_4273;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_5896;
wire n_4567;
wire n_5833;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_3749;
wire n_5691;
wire n_3482;
wire n_5403;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_2956;
wire n_5210;
wire n_2382;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_3458;
wire n_5843;
wire n_3511;
wire n_2077;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_6156;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_5913;
wire n_4530;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_5968;
wire n_3549;
wire n_3914;
wire n_5586;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_5056;
wire n_2015;
wire n_5984;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_1787;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_2257;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_3559;
wire n_5778;
wire n_5179;
wire n_2435;
wire n_5680;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_5549;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_2954;
wire n_4438;
wire n_3814;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_2019;
wire n_5708;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2649;
wire n_6033;
wire n_2919;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_2632;
wire n_5557;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_3087;
wire n_6009;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_5773;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_5149;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_5858;
wire n_5985;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_4292;
wire n_2118;
wire n_5552;
wire n_6074;
wire n_3764;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_2125;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_2707;
wire n_5596;
wire n_2849;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_3713;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_5889;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_2821;
wire n_3696;
wire n_4781;
wire n_6031;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_2448;
wire n_2211;
wire n_5904;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_2958;
wire n_4429;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_5511;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_6036;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_3753;
wire n_4846;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_3421;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_5921;
wire n_1849;
wire n_4966;
wire n_2250;
wire n_6104;
wire n_3321;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_4202;
wire n_2044;
wire n_5679;
wire n_3886;
wire n_2619;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_2613;
wire n_5667;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_5027;
wire n_2343;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_1921;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_5999;
wire n_2110;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_4355;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_4060;
wire n_2459;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_6075;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_3630;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2672;
wire n_2018;
wire n_2602;
wire n_5780;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_5743;
wire n_1956;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_6022;
wire n_2828;
wire n_5950;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_5705;
wire n_4996;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_5848;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_3963;
wire n_3091;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_4628;
wire n_5982;
wire n_1775;
wire n_4083;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_3940;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_5763;
wire n_3633;
wire n_6061;
wire n_4001;
wire n_2584;
wire n_5701;
wire n_3111;
wire n_1813;
wire n_2997;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_1996;
wire n_2009;
wire n_5907;
wire n_4339;
wire n_6013;
wire n_4690;
wire n_2987;
wire n_5895;
wire n_2651;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_3632;
wire n_2522;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_3457;
wire n_5384;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_3768;
wire n_4295;
wire n_4100;
wire n_2372;
wire n_3445;
wire n_2105;
wire n_1806;
wire n_4087;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_4266;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_5844;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_4976;
wire n_3555;
wire n_5938;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_2148;
wire n_5548;
wire n_4663;
wire n_5840;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_4686;
wire n_2384;
wire n_3707;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_3058;
wire n_5355;
wire n_2047;
wire n_3398;
wire n_3709;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_3399;
wire n_4772;
wire n_5915;
wire n_4120;
wire n_2880;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_5116;
wire n_3771;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_6046;
wire n_4493;
wire n_6055;
wire n_1808;
wire n_6091;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_6144;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_4901;
wire n_3480;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_4602;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_5901;
wire n_2837;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_3154;
wire n_3938;
wire n_2278;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_2579;
wire n_1961;
wire n_2960;
wire n_3270;
wire n_2844;
wire n_1979;
wire n_4814;
wire n_6178;
wire n_2221;
wire n_5502;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_6000;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_4831;
wire n_4782;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_5703;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_4147;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_2685;
wire n_2061;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_5264;
wire n_2595;
wire n_3084;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_2981;
wire n_4995;
wire n_5873;
wire n_4498;
wire n_5741;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_2466;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_3460;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_2693;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_5130;
wire n_4175;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_5992;
wire n_2601;
wire n_2172;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_5981;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_3046;
wire n_2293;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_4003;
wire n_1832;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_2495;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_2535;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_3138;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_2296;
wire n_5735;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_6037;
wire n_4186;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_3377;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_5935;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_5488;
wire n_5727;
wire n_3599;
wire n_5988;
wire n_5646;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_5832;
wire n_3401;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_5470;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_2218;
wire n_2593;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_3995;
wire n_3908;
wire n_3892;
wire n_3501;
wire n_3216;
wire n_2555;
wire n_3568;
wire n_2708;
wire n_4844;
wire n_4049;
wire n_2661;
wire n_2470;
wire n_3551;
wire n_5037;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_4324;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_3459;
wire n_2576;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_3735;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_2900;
wire n_2912;
wire n_5936;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_2928;
wire n_5505;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_5504;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_2730;
wire n_5129;
wire n_4704;
wire n_2720;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_2700;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_3317;
wire n_5653;
wire n_4835;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_4727;
wire n_3654;
wire n_5627;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_6026;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_5697;
wire n_2020;
wire n_5606;
wire n_2310;
wire n_5911;
wire n_3600;
wire n_6139;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_3967;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_5841;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_3344;
wire n_4754;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_3117;
wire n_4684;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_5043;
wire n_4241;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6107;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_5035;
wire n_3037;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_2007;
wire n_3363;
wire n_1803;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_5631;
wire n_3481;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_5608;
wire n_2204;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_4217;
wire n_5277;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_2428;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_4592;
wire n_4999;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_2589;
wire n_4086;
wire n_4656;
wire n_4862;
wire n_5687;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_4177;
wire n_2501;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_6105;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_3278;
wire n_2375;
wire n_5579;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_6163;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_2358;
wire n_3546;
wire n_2355;
wire n_5887;
wire n_3068;
wire n_5683;
wire n_3002;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_2351;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_1941;
wire n_3637;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_6015;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_2297;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_4698;
wire n_3674;
wire n_5349;
wire n_3763;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_2421;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_6120;
wire n_3557;
wire n_2269;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_2361;
wire n_1752;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_2239;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_2304;
wire n_2514;
wire n_5932;
wire n_6121;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_5823;
wire n_2423;
wire n_2208;
wire n_5422;
wire n_5944;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_4834;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_2346;
wire n_4692;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_4299;
wire n_5625;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_5570;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_5978;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_4625;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_5575;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_2735;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_2109;
wire n_2709;
wire n_3419;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_5607;
wire n_2782;
wire n_3929;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6005;
wire n_2060;
wire n_3883;
wire n_4032;
wire n_2571;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_5140;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_5847;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_4884;
wire n_3580;
wire n_4276;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_5718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_5658;
wire n_4174;
wire n_5131;
wire n_5546;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_4394;
wire n_5544;
wire n_5660;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_5610;
wire n_2810;
wire n_1884;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_5808;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_2925;
wire n_1750;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_5710;
wire n_2628;
wire n_3219;
wire n_5333;
wire n_5799;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_3688;
wire n_5008;
wire n_3871;
wire n_3757;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_3479;
wire n_5499;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_2755;
wire n_5109;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_2220;
wire n_6108;
wire n_6100;
wire n_4433;
wire n_2829;
wire n_5862;
wire n_1914;
wire n_2253;
wire n_5886;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_5883;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_5630;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_2113;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_5132;
wire n_3498;
wire n_2350;
wire n_5535;
wire n_4506;
wire n_6097;
wire n_6057;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_2187;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_4359;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_5793;
wire n_1798;
wire n_3057;
wire n_5761;
wire n_3983;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_4348;
wire n_3139;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_4084;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_3984;
wire n_4389;
wire n_1763;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_2660;
wire n_1859;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_5657;
wire n_2379;
wire n_3579;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_4387;
wire n_3186;
wire n_2508;
wire n_2594;
wire n_5298;
wire n_3417;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1729;
wire n_6067;
wire n_2893;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_2280;
wire n_5867;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_5798;
wire n_4137;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_4535;
wire n_4385;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1733;
wire n_4651;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_3050;
wire n_3919;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_3718;
wire n_3390;
wire n_2298;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_5903;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_5446;
wire n_4561;
wire n_3291;
wire n_2578;
wire n_2475;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_3358;
wire n_2533;
wire n_2003;
wire n_4682;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_3289;
wire n_1955;
wire n_6127;
wire n_5005;
wire n_6126;
wire n_6151;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_3131;
wire n_1973;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_6007;
wire n_1772;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_5996;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_5652;
wire n_5805;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_4973;
wire n_4792;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_6093;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_5902;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_5952;
wire n_2086;
wire n_1926;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2597;
wire n_2321;
wire n_5980;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_2186;
wire n_5790;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_5485;
wire n_5525;
wire n_3004;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_5850;
wire n_4564;
wire n_1848;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_4080;
wire n_2206;
wire n_4185;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_5860;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_6143;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_5859;
wire n_4390;
wire n_1782;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_6175;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_5172;
wire n_1982;
wire n_5311;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2982;
wire n_5495;
wire n_4483;
wire n_3061;
wire n_3504;
wire n_2587;
wire n_5547;
wire n_4693;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_3779;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_1891;
wire n_5348;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_3045;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_1905;
wire n_5448;
wire n_2573;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_3033;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_5900;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_5851;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_2461;
wire n_3719;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_5295;
wire n_6088;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_3965;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_2323;
wire n_4549;
wire n_1746;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_5656;
wire n_1988;
wire n_5678;
wire n_5865;
wire n_6050;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_4809;
wire n_4012;
wire n_2049;
wire n_5212;
wire n_4760;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_5965;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_5042;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_5368;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_4360;
wire n_4540;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_3089;
wire n_4854;
wire n_5477;
wire n_2727;
wire n_5234;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_2499;
wire n_2549;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_5659;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_5598;
wire n_2753;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_5783;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_2378;
wire n_5530;
wire n_5809;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_5993;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_3170;
wire n_2311;
wire n_2287;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_3467;
wire n_5821;
wire n_3179;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_3699;
wire n_6118;
wire n_2120;
wire n_6028;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2757;
wire n_2168;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_5943;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_2801;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_1869;
wire n_3623;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_3471;
wire n_4075;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_5209;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_3009;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_3957;
wire n_3418;
wire n_5673;
wire n_5814;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_6040;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_5769;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_5181;
wire n_3208;
wire n_5768;
wire n_2737;
wire n_3282;
wire n_2916;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_5972;
wire n_3400;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1993;
wire n_4035;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5577;
wire n_5872;
wire n_5017;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_5838;
wire n_3694;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_4065;
wire n_4705;
wire n_1971;
wire n_2945;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_6039;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_5401;
wire n_4595;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_6021;
wire n_4617;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_3769;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_5986;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_3509;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_5863;
wire n_3790;
wire n_6152;
wire n_5734;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_5600;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_5767;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_2600;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_3686;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_2141;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_3677;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_2488;
wire n_6134;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_5714;
wire n_2169;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_2724;
wire n_2258;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_2268;
wire n_3469;
wire n_2835;
wire n_5835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_6092;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_3898;
wire n_4749;
wire n_5924;
wire n_1845;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_4238;
wire n_2005;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_4668;
wire n_5782;
wire n_4168;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_5034;
wire n_3312;
wire n_2451;
wire n_2913;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_5927;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_4890;
wire n_2485;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_5226;
wire n_2081;
wire n_1794;
wire n_5696;
wire n_5014;
wire n_3053;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_4516;
wire n_5235;
wire n_2798;
wire n_3217;
wire n_6081;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

INVx2_ASAP7_75t_L g1718 ( 
.A(n_983),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_459),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1169),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_813),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_530),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1574),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_74),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_582),
.Y(n_1725)
);

CKINVDCx16_ASAP7_75t_R g1726 ( 
.A(n_1374),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_898),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1687),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_884),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1120),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1567),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_465),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1291),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1586),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1637),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_132),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_999),
.Y(n_1737)
);

CKINVDCx14_ASAP7_75t_R g1738 ( 
.A(n_1619),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_84),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_947),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_902),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1215),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1035),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1209),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_649),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1059),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1074),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1568),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1493),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1584),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1468),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1653),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1392),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1058),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1114),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_289),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1616),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_80),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_27),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_426),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_919),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_200),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_739),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1547),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1274),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_938),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1425),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_63),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_800),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1550),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_354),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_650),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_150),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_941),
.Y(n_1774)
);

BUFx10_ASAP7_75t_L g1775 ( 
.A(n_1436),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_220),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1256),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1331),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_499),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1530),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_480),
.Y(n_1781)
);

BUFx10_ASAP7_75t_L g1782 ( 
.A(n_1539),
.Y(n_1782)
);

BUFx10_ASAP7_75t_L g1783 ( 
.A(n_350),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1400),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1558),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_585),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_556),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_851),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_304),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_521),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_859),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_649),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_816),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_37),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_365),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1477),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_139),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_977),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_1434),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1516),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1569),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1112),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_178),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_852),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1406),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_34),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_644),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_595),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1315),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_596),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1511),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1068),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1491),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_449),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1110),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1548),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1252),
.Y(n_1817)
);

BUFx10_ASAP7_75t_L g1818 ( 
.A(n_164),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_865),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1015),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_749),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1617),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_874),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_91),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1216),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1008),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1129),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1591),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_230),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_889),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1519),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_879),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_328),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1104),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1604),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1112),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_773),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1505),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_523),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1461),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_625),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1543),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1560),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1606),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1244),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_470),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1010),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_29),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1678),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_506),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_622),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_548),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1302),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1254),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1509),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_600),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1646),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1188),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_665),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1479),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_638),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_126),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_361),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_269),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1231),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1709),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1667),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1324),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_1258),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1075),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_290),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_650),
.Y(n_1872)
);

CKINVDCx16_ASAP7_75t_R g1873 ( 
.A(n_1399),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1370),
.Y(n_1874)
);

BUFx2_ASAP7_75t_R g1875 ( 
.A(n_1451),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1077),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_698),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1593),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1684),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_464),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1334),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1579),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_634),
.Y(n_1883)
);

BUFx10_ASAP7_75t_L g1884 ( 
.A(n_1343),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_588),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1711),
.Y(n_1886)
);

BUFx2_ASAP7_75t_R g1887 ( 
.A(n_1073),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1253),
.Y(n_1888)
);

BUFx10_ASAP7_75t_L g1889 ( 
.A(n_1478),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_758),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1241),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_914),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_374),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1575),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_710),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_780),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1009),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1541),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_917),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1384),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1639),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_22),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1677),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_69),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1588),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1360),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_851),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1647),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_698),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1399),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1345),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_425),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1659),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1301),
.Y(n_1914)
);

INVx2_ASAP7_75t_SL g1915 ( 
.A(n_805),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1638),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1589),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1510),
.Y(n_1918)
);

BUFx10_ASAP7_75t_L g1919 ( 
.A(n_520),
.Y(n_1919)
);

CKINVDCx20_ASAP7_75t_R g1920 ( 
.A(n_169),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1101),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1630),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_288),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_449),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1457),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1163),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1556),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1609),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_550),
.Y(n_1929)
);

CKINVDCx20_ASAP7_75t_R g1930 ( 
.A(n_919),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1007),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_811),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_526),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1666),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_731),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_50),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_799),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1018),
.Y(n_1938)
);

CKINVDCx16_ASAP7_75t_R g1939 ( 
.A(n_1498),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1042),
.Y(n_1940)
);

BUFx8_ASAP7_75t_SL g1941 ( 
.A(n_66),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1533),
.Y(n_1942)
);

CKINVDCx20_ASAP7_75t_R g1943 ( 
.A(n_551),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_747),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_961),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1063),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_776),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1610),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1323),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1380),
.Y(n_1950)
);

CKINVDCx16_ASAP7_75t_R g1951 ( 
.A(n_68),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_525),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1589),
.Y(n_1953)
);

CKINVDCx14_ASAP7_75t_R g1954 ( 
.A(n_1168),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_861),
.Y(n_1955)
);

INVx2_ASAP7_75t_SL g1956 ( 
.A(n_1537),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1165),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1586),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_573),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1623),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_926),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1307),
.Y(n_1962)
);

BUFx8_ASAP7_75t_SL g1963 ( 
.A(n_770),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1420),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1118),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_914),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_752),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1518),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1611),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1095),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1038),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1526),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_358),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_159),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1191),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_323),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_71),
.Y(n_1977)
);

CKINVDCx14_ASAP7_75t_R g1978 ( 
.A(n_541),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_936),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1433),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_349),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_543),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1655),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1324),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1287),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1180),
.Y(n_1986)
);

CKINVDCx14_ASAP7_75t_R g1987 ( 
.A(n_1514),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_673),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1385),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_928),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_647),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1494),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_498),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_965),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1522),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_849),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_495),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1686),
.Y(n_1998)
);

CKINVDCx16_ASAP7_75t_R g1999 ( 
.A(n_247),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1267),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_244),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_223),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1680),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1419),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1305),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1665),
.Y(n_2006)
);

CKINVDCx20_ASAP7_75t_R g2007 ( 
.A(n_1691),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1513),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1296),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1510),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_440),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1454),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_784),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_948),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1117),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1030),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_60),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1391),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1668),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_441),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1654),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_706),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_31),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1585),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_765),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_406),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_925),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_906),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1362),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_866),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1500),
.Y(n_2031)
);

CKINVDCx20_ASAP7_75t_R g2032 ( 
.A(n_1551),
.Y(n_2032)
);

BUFx3_ASAP7_75t_L g2033 ( 
.A(n_1405),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_777),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_456),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_151),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1600),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1566),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_91),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_385),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1133),
.Y(n_2041)
);

CKINVDCx16_ASAP7_75t_R g2042 ( 
.A(n_579),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1366),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_1651),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_15),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1283),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1693),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1578),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1580),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1067),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_976),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1656),
.Y(n_2052)
);

INVx2_ASAP7_75t_SL g2053 ( 
.A(n_445),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_801),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_911),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_365),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1272),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_113),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_290),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1052),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_262),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1063),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_996),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_881),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_37),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_621),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1216),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1308),
.Y(n_2068)
);

CKINVDCx20_ASAP7_75t_R g2069 ( 
.A(n_1146),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1662),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_829),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1511),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1458),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1053),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_70),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_431),
.Y(n_2076)
);

BUFx5_ASAP7_75t_L g2077 ( 
.A(n_1494),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_185),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1512),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_428),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1310),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_437),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1555),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1068),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1109),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_466),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1587),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1396),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1621),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1209),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1645),
.Y(n_2091)
);

CKINVDCx16_ASAP7_75t_R g2092 ( 
.A(n_807),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1658),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1620),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_344),
.Y(n_2095)
);

CKINVDCx20_ASAP7_75t_R g2096 ( 
.A(n_203),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1649),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1139),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_559),
.Y(n_2099)
);

CKINVDCx20_ASAP7_75t_R g2100 ( 
.A(n_1042),
.Y(n_2100)
);

CKINVDCx14_ASAP7_75t_R g2101 ( 
.A(n_1598),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1504),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1313),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1487),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1403),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_555),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1102),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_396),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_610),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_508),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_1410),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_297),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_668),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1264),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_964),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1398),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1174),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_154),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_1599),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1583),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1608),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1428),
.Y(n_2122)
);

INVxp67_ASAP7_75t_L g2123 ( 
.A(n_1607),
.Y(n_2123)
);

BUFx10_ASAP7_75t_L g2124 ( 
.A(n_699),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1627),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_720),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1453),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1122),
.Y(n_2128)
);

BUFx10_ASAP7_75t_L g2129 ( 
.A(n_849),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_982),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_294),
.Y(n_2131)
);

CKINVDCx20_ASAP7_75t_R g2132 ( 
.A(n_1338),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1591),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1526),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_200),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_799),
.Y(n_2136)
);

BUFx10_ASAP7_75t_L g2137 ( 
.A(n_35),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_558),
.Y(n_2138)
);

BUFx10_ASAP7_75t_L g2139 ( 
.A(n_1091),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1495),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_1382),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_645),
.Y(n_2142)
);

CKINVDCx20_ASAP7_75t_R g2143 ( 
.A(n_1282),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1211),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1546),
.Y(n_2145)
);

INVx1_ASAP7_75t_SL g2146 ( 
.A(n_448),
.Y(n_2146)
);

BUFx10_ASAP7_75t_L g2147 ( 
.A(n_284),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_617),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_317),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_1528),
.Y(n_2150)
);

BUFx10_ASAP7_75t_L g2151 ( 
.A(n_1206),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1178),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1703),
.Y(n_2153)
);

BUFx10_ASAP7_75t_L g2154 ( 
.A(n_146),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1565),
.Y(n_2155)
);

INVx1_ASAP7_75t_SL g2156 ( 
.A(n_607),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_415),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_529),
.Y(n_2158)
);

BUFx10_ASAP7_75t_L g2159 ( 
.A(n_1017),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_609),
.Y(n_2160)
);

INVx2_ASAP7_75t_SL g2161 ( 
.A(n_1030),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1698),
.Y(n_2162)
);

CKINVDCx20_ASAP7_75t_R g2163 ( 
.A(n_1309),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_1260),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1677),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_791),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1155),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1386),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1576),
.Y(n_2169)
);

CKINVDCx20_ASAP7_75t_R g2170 ( 
.A(n_1707),
.Y(n_2170)
);

CKINVDCx20_ASAP7_75t_R g2171 ( 
.A(n_268),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1181),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_465),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1015),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1197),
.Y(n_2175)
);

INVx1_ASAP7_75t_SL g2176 ( 
.A(n_1652),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_923),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1598),
.Y(n_2178)
);

CKINVDCx20_ASAP7_75t_R g2179 ( 
.A(n_1611),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_622),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_859),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_16),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_413),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1198),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1709),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1602),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_1132),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_662),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1445),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_1692),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1573),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_65),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_333),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_347),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_367),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_106),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_235),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1508),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1532),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_254),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_839),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1492),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1219),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_1527),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_312),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1428),
.Y(n_2206)
);

CKINVDCx5p33_ASAP7_75t_R g2207 ( 
.A(n_1582),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1116),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1660),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1618),
.Y(n_2210)
);

INVxp67_ASAP7_75t_L g2211 ( 
.A(n_1207),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_917),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1549),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1471),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_942),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1202),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_308),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1320),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_639),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_774),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1626),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1529),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_534),
.Y(n_2223)
);

CKINVDCx5p33_ASAP7_75t_R g2224 ( 
.A(n_771),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_1602),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_161),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_293),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_548),
.Y(n_2228)
);

BUFx10_ASAP7_75t_L g2229 ( 
.A(n_1424),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_148),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_792),
.Y(n_2231)
);

BUFx2_ASAP7_75t_L g2232 ( 
.A(n_795),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_270),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_881),
.Y(n_2234)
);

BUFx8_ASAP7_75t_SL g2235 ( 
.A(n_1536),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1184),
.Y(n_2236)
);

CKINVDCx20_ASAP7_75t_R g2237 ( 
.A(n_1633),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_504),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1592),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1644),
.Y(n_2240)
);

BUFx10_ASAP7_75t_L g2241 ( 
.A(n_847),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_666),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_28),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_259),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_1515),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_971),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_719),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1499),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_507),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_287),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_295),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1692),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_86),
.Y(n_2253)
);

INVxp33_ASAP7_75t_R g2254 ( 
.A(n_1597),
.Y(n_2254)
);

BUFx5_ASAP7_75t_L g2255 ( 
.A(n_1503),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_1052),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1298),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1083),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_1322),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1321),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1529),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_1026),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1236),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_707),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_876),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_995),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1541),
.Y(n_2267)
);

BUFx10_ASAP7_75t_L g2268 ( 
.A(n_556),
.Y(n_2268)
);

BUFx10_ASAP7_75t_L g2269 ( 
.A(n_1433),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_511),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_271),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1405),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1628),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_655),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_1272),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_53),
.Y(n_2276)
);

CKINVDCx5p33_ASAP7_75t_R g2277 ( 
.A(n_1497),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1668),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_942),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_980),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1046),
.Y(n_2281)
);

CKINVDCx16_ASAP7_75t_R g2282 ( 
.A(n_1205),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1563),
.Y(n_2283)
);

CKINVDCx16_ASAP7_75t_R g2284 ( 
.A(n_1506),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_38),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_1060),
.Y(n_2286)
);

BUFx10_ASAP7_75t_L g2287 ( 
.A(n_319),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_753),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_1502),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_585),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_251),
.Y(n_2291)
);

BUFx10_ASAP7_75t_L g2292 ( 
.A(n_1158),
.Y(n_2292)
);

BUFx2_ASAP7_75t_SL g2293 ( 
.A(n_1623),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_507),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_141),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1394),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_162),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1263),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_1348),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_872),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_1142),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_1595),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_982),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_193),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_545),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_74),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_1590),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_1033),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1629),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1648),
.Y(n_2310)
);

BUFx10_ASAP7_75t_L g2311 ( 
.A(n_84),
.Y(n_2311)
);

CKINVDCx20_ASAP7_75t_R g2312 ( 
.A(n_57),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1637),
.Y(n_2313)
);

CKINVDCx20_ASAP7_75t_R g2314 ( 
.A(n_101),
.Y(n_2314)
);

BUFx10_ASAP7_75t_L g2315 ( 
.A(n_1596),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_605),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_1201),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1188),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_1214),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_87),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_941),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_175),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_938),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_545),
.Y(n_2324)
);

CKINVDCx16_ASAP7_75t_R g2325 ( 
.A(n_1501),
.Y(n_2325)
);

CKINVDCx14_ASAP7_75t_R g2326 ( 
.A(n_1235),
.Y(n_2326)
);

CKINVDCx5p33_ASAP7_75t_R g2327 ( 
.A(n_1372),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1576),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_1128),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_181),
.Y(n_2330)
);

CKINVDCx20_ASAP7_75t_R g2331 ( 
.A(n_35),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_339),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_77),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1650),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_299),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1119),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_1636),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_1538),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1631),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_328),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_522),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_1357),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_1115),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1133),
.Y(n_2344)
);

CKINVDCx16_ASAP7_75t_R g2345 ( 
.A(n_145),
.Y(n_2345)
);

BUFx10_ASAP7_75t_L g2346 ( 
.A(n_1545),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_1344),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_857),
.Y(n_2348)
);

BUFx2_ASAP7_75t_SL g2349 ( 
.A(n_1041),
.Y(n_2349)
);

INVxp67_ASAP7_75t_SL g2350 ( 
.A(n_1560),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_863),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_772),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1056),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_923),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_329),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1159),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_519),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_1170),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1002),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_798),
.Y(n_2360)
);

CKINVDCx20_ASAP7_75t_R g2361 ( 
.A(n_1407),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_242),
.Y(n_2362)
);

INVx1_ASAP7_75t_SL g2363 ( 
.A(n_1299),
.Y(n_2363)
);

CKINVDCx20_ASAP7_75t_R g2364 ( 
.A(n_1121),
.Y(n_2364)
);

INVx1_ASAP7_75t_SL g2365 ( 
.A(n_58),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_1212),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_1699),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1520),
.Y(n_2368)
);

INVxp67_ASAP7_75t_L g2369 ( 
.A(n_676),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_699),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_824),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_996),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_1669),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_467),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_1232),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1379),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_130),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_1224),
.Y(n_2378)
);

BUFx5_ASAP7_75t_L g2379 ( 
.A(n_915),
.Y(n_2379)
);

CKINVDCx20_ASAP7_75t_R g2380 ( 
.A(n_1081),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1438),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_1554),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_445),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_1603),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_1408),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_554),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_1204),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_1282),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_739),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_1520),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_1594),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_276),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_751),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1613),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_554),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1679),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1534),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_525),
.Y(n_2398)
);

BUFx10_ASAP7_75t_L g2399 ( 
.A(n_1682),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_1705),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_1250),
.Y(n_2401)
);

HB1xp67_ASAP7_75t_L g2402 ( 
.A(n_1606),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_662),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1326),
.Y(n_2404)
);

CKINVDCx20_ASAP7_75t_R g2405 ( 
.A(n_1441),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_1199),
.Y(n_2406)
);

BUFx3_ASAP7_75t_L g2407 ( 
.A(n_620),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_1570),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_358),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_4),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_1625),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_222),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_276),
.Y(n_2413)
);

CKINVDCx20_ASAP7_75t_R g2414 ( 
.A(n_482),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1085),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_1158),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_1504),
.Y(n_2417)
);

CKINVDCx16_ASAP7_75t_R g2418 ( 
.A(n_1465),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_1571),
.Y(n_2419)
);

BUFx3_ASAP7_75t_L g2420 ( 
.A(n_320),
.Y(n_2420)
);

CKINVDCx20_ASAP7_75t_R g2421 ( 
.A(n_486),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_845),
.Y(n_2422)
);

CKINVDCx5p33_ASAP7_75t_R g2423 ( 
.A(n_575),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_1027),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_595),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1542),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1501),
.Y(n_2427)
);

CKINVDCx14_ASAP7_75t_R g2428 ( 
.A(n_1523),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_1124),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_199),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_829),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_66),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_224),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_1018),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_1031),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_530),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_788),
.Y(n_2437)
);

CKINVDCx20_ASAP7_75t_R g2438 ( 
.A(n_1552),
.Y(n_2438)
);

CKINVDCx20_ASAP7_75t_R g2439 ( 
.A(n_1553),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_443),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_634),
.Y(n_2441)
);

INVx2_ASAP7_75t_SL g2442 ( 
.A(n_1664),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_1026),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_1634),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_1674),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_1260),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_1011),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_1134),
.Y(n_2448)
);

INVxp33_ASAP7_75t_R g2449 ( 
.A(n_1521),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_862),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_1479),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_182),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_883),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_1115),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_241),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_42),
.Y(n_2456)
);

INVx1_ASAP7_75t_SL g2457 ( 
.A(n_674),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_1496),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_1657),
.Y(n_2459)
);

INVx2_ASAP7_75t_SL g2460 ( 
.A(n_597),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_5),
.Y(n_2461)
);

BUFx8_ASAP7_75t_SL g2462 ( 
.A(n_1034),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_1582),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_248),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_909),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_1540),
.Y(n_2466)
);

CKINVDCx20_ASAP7_75t_R g2467 ( 
.A(n_939),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_1614),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1469),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_1568),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_70),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_1632),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_800),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_1154),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_825),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_1643),
.Y(n_2476)
);

HB1xp67_ASAP7_75t_L g2477 ( 
.A(n_541),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_1103),
.Y(n_2478)
);

CKINVDCx20_ASAP7_75t_R g2479 ( 
.A(n_1019),
.Y(n_2479)
);

BUFx5_ASAP7_75t_L g2480 ( 
.A(n_175),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1196),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_779),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_274),
.Y(n_2483)
);

CKINVDCx20_ASAP7_75t_R g2484 ( 
.A(n_185),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_499),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_1470),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_51),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_474),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_308),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_1700),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_1665),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_695),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_765),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_302),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_1635),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_1035),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_1588),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_1449),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_1174),
.Y(n_2499)
);

BUFx5_ASAP7_75t_L g2500 ( 
.A(n_978),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_484),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_1204),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_1321),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_283),
.Y(n_2504)
);

INVx1_ASAP7_75t_SL g2505 ( 
.A(n_125),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_1601),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_1664),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_412),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_931),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_14),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_1564),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_385),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_990),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_1281),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_1373),
.Y(n_2515)
);

CKINVDCx14_ASAP7_75t_R g2516 ( 
.A(n_1185),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_1020),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_1346),
.Y(n_2518)
);

BUFx3_ASAP7_75t_L g2519 ( 
.A(n_1072),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_270),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_157),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_1561),
.Y(n_2522)
);

CKINVDCx20_ASAP7_75t_R g2523 ( 
.A(n_375),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_977),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_46),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_771),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_495),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_134),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_1507),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_1601),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1327),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_1393),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_1605),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_1183),
.Y(n_2534)
);

INVxp67_ASAP7_75t_L g2535 ( 
.A(n_1506),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_559),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_527),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_968),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_1407),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_1391),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_1297),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_1319),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_1378),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_631),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_1022),
.Y(n_2545)
);

BUFx2_ASAP7_75t_L g2546 ( 
.A(n_776),
.Y(n_2546)
);

CKINVDCx20_ASAP7_75t_R g2547 ( 
.A(n_184),
.Y(n_2547)
);

CKINVDCx16_ASAP7_75t_R g2548 ( 
.A(n_1289),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_1531),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_112),
.Y(n_2550)
);

BUFx2_ASAP7_75t_L g2551 ( 
.A(n_27),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_1306),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_388),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_1612),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_802),
.Y(n_2555)
);

INVx1_ASAP7_75t_SL g2556 ( 
.A(n_265),
.Y(n_2556)
);

INVx2_ASAP7_75t_SL g2557 ( 
.A(n_285),
.Y(n_2557)
);

CKINVDCx20_ASAP7_75t_R g2558 ( 
.A(n_1103),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_1615),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_1685),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1559),
.Y(n_2561)
);

CKINVDCx16_ASAP7_75t_R g2562 ( 
.A(n_961),
.Y(n_2562)
);

BUFx2_ASAP7_75t_L g2563 ( 
.A(n_910),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_1661),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_1517),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_562),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_1410),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_880),
.Y(n_2568)
);

BUFx5_ASAP7_75t_L g2569 ( 
.A(n_70),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_626),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_576),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_246),
.Y(n_2572)
);

CKINVDCx14_ASAP7_75t_R g2573 ( 
.A(n_470),
.Y(n_2573)
);

CKINVDCx20_ASAP7_75t_R g2574 ( 
.A(n_995),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_259),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_623),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_1581),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_1525),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_314),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_173),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_258),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_1076),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_130),
.Y(n_2583)
);

CKINVDCx5p33_ASAP7_75t_R g2584 ( 
.A(n_1624),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_1078),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_1259),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_1311),
.Y(n_2587)
);

CKINVDCx20_ASAP7_75t_R g2588 ( 
.A(n_1150),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_558),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_543),
.Y(n_2590)
);

CKINVDCx20_ASAP7_75t_R g2591 ( 
.A(n_866),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_464),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_232),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_870),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_404),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_1615),
.Y(n_2596)
);

BUFx10_ASAP7_75t_L g2597 ( 
.A(n_157),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_1376),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_1498),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_1524),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_1447),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_857),
.Y(n_2602)
);

BUFx3_ASAP7_75t_L g2603 ( 
.A(n_608),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_1594),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_701),
.Y(n_2605)
);

CKINVDCx20_ASAP7_75t_R g2606 ( 
.A(n_762),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_970),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_547),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_1081),
.Y(n_2609)
);

CKINVDCx20_ASAP7_75t_R g2610 ( 
.A(n_1557),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_1400),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_1361),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_1680),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_798),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_404),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_1572),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_1622),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_1034),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_1610),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1640),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_964),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_1641),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_1241),
.Y(n_2623)
);

BUFx6f_ASAP7_75t_L g2624 ( 
.A(n_679),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_22),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_604),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_940),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_557),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_1377),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_1390),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_1562),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_1392),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_32),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_15),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_1577),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_1131),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_901),
.Y(n_2637)
);

INVx1_ASAP7_75t_SL g2638 ( 
.A(n_288),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_557),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_1538),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_1032),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_149),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_5),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_588),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_1593),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_1530),
.Y(n_2646)
);

INVx2_ASAP7_75t_SL g2647 ( 
.A(n_1366),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_1454),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_1458),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_540),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_33),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_1425),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_837),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_198),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_1663),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_1389),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_1448),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_1535),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_1544),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_433),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_1642),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_311),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_1192),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_1883),
.Y(n_2664)
);

INVxp33_ASAP7_75t_SL g2665 ( 
.A(n_1785),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_1951),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1892),
.Y(n_2667)
);

INVxp33_ASAP7_75t_L g2668 ( 
.A(n_1941),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2187),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_1963),
.Y(n_2670)
);

INVxp67_ASAP7_75t_L g2671 ( 
.A(n_1757),
.Y(n_2671)
);

CKINVDCx16_ASAP7_75t_R g2672 ( 
.A(n_1738),
.Y(n_2672)
);

INVxp33_ASAP7_75t_SL g2673 ( 
.A(n_2177),
.Y(n_2673)
);

INVxp67_ASAP7_75t_SL g2674 ( 
.A(n_2461),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2235),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2480),
.Y(n_2676)
);

INVxp67_ASAP7_75t_SL g2677 ( 
.A(n_2461),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2480),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2462),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2480),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2345),
.Y(n_2681)
);

INVxp67_ASAP7_75t_L g2682 ( 
.A(n_1912),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_1726),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2480),
.Y(n_2684)
);

INVxp33_ASAP7_75t_L g2685 ( 
.A(n_2337),
.Y(n_2685)
);

CKINVDCx20_ASAP7_75t_R g2686 ( 
.A(n_1954),
.Y(n_2686)
);

INVxp67_ASAP7_75t_SL g2687 ( 
.A(n_2461),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_1873),
.Y(n_2688)
);

BUFx2_ASAP7_75t_L g2689 ( 
.A(n_2551),
.Y(n_2689)
);

INVxp67_ASAP7_75t_SL g2690 ( 
.A(n_1724),
.Y(n_2690)
);

INVxp67_ASAP7_75t_L g2691 ( 
.A(n_1940),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2569),
.Y(n_2692)
);

INVxp33_ASAP7_75t_L g2693 ( 
.A(n_2402),
.Y(n_2693)
);

INVxp67_ASAP7_75t_SL g2694 ( 
.A(n_1758),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2569),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2569),
.Y(n_2696)
);

INVxp33_ASAP7_75t_L g2697 ( 
.A(n_2464),
.Y(n_2697)
);

INVxp67_ASAP7_75t_SL g2698 ( 
.A(n_1794),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2077),
.Y(n_2699)
);

INVxp33_ASAP7_75t_SL g2700 ( 
.A(n_2477),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2077),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2077),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2077),
.Y(n_2703)
);

CKINVDCx16_ASAP7_75t_R g2704 ( 
.A(n_1978),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2255),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_1939),
.Y(n_2706)
);

INVxp67_ASAP7_75t_SL g2707 ( 
.A(n_1797),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2255),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_1999),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2255),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_1987),
.Y(n_2711)
);

INVxp67_ASAP7_75t_SL g2712 ( 
.A(n_1848),
.Y(n_2712)
);

CKINVDCx16_ASAP7_75t_R g2713 ( 
.A(n_2101),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2255),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2379),
.Y(n_2715)
);

CKINVDCx20_ASAP7_75t_R g2716 ( 
.A(n_2326),
.Y(n_2716)
);

INVxp33_ASAP7_75t_SL g2717 ( 
.A(n_1739),
.Y(n_2717)
);

CKINVDCx16_ASAP7_75t_R g2718 ( 
.A(n_2428),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2379),
.Y(n_2719)
);

INVxp67_ASAP7_75t_SL g2720 ( 
.A(n_1862),
.Y(n_2720)
);

INVxp67_ASAP7_75t_SL g2721 ( 
.A(n_1902),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2042),
.Y(n_2722)
);

INVxp67_ASAP7_75t_SL g2723 ( 
.A(n_1977),
.Y(n_2723)
);

INVxp33_ASAP7_75t_SL g2724 ( 
.A(n_1759),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_1779),
.Y(n_2725)
);

CKINVDCx20_ASAP7_75t_R g2726 ( 
.A(n_2516),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2379),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2379),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_1779),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2500),
.Y(n_2730)
);

CKINVDCx20_ASAP7_75t_R g2731 ( 
.A(n_2573),
.Y(n_2731)
);

CKINVDCx20_ASAP7_75t_R g2732 ( 
.A(n_1721),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2500),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2092),
.Y(n_2734)
);

BUFx2_ASAP7_75t_L g2735 ( 
.A(n_1976),
.Y(n_2735)
);

BUFx2_ASAP7_75t_L g2736 ( 
.A(n_1989),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2500),
.Y(n_2737)
);

INVxp67_ASAP7_75t_SL g2738 ( 
.A(n_2023),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2500),
.Y(n_2739)
);

INVxp67_ASAP7_75t_SL g2740 ( 
.A(n_2036),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2039),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2045),
.Y(n_2742)
);

CKINVDCx16_ASAP7_75t_R g2743 ( 
.A(n_2282),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2058),
.Y(n_2744)
);

CKINVDCx20_ASAP7_75t_R g2745 ( 
.A(n_1799),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2065),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2075),
.Y(n_2747)
);

INVxp33_ASAP7_75t_L g2748 ( 
.A(n_2232),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2118),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2196),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2297),
.Y(n_2751)
);

CKINVDCx16_ASAP7_75t_R g2752 ( 
.A(n_2284),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2410),
.Y(n_2753)
);

CKINVDCx20_ASAP7_75t_R g2754 ( 
.A(n_1802),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2452),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2456),
.Y(n_2756)
);

INVxp67_ASAP7_75t_L g2757 ( 
.A(n_2416),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_2659),
.Y(n_2758)
);

CKINVDCx14_ASAP7_75t_R g2759 ( 
.A(n_1818),
.Y(n_2759)
);

CKINVDCx20_ASAP7_75t_R g2760 ( 
.A(n_1869),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_1736),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2521),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2525),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2243),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2471),
.Y(n_2765)
);

CKINVDCx20_ASAP7_75t_R g2766 ( 
.A(n_1893),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2510),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2651),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_1779),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_1722),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_1725),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_1868),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_2325),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_1727),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2546),
.B(n_0),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_1729),
.Y(n_2776)
);

CKINVDCx20_ASAP7_75t_R g2777 ( 
.A(n_1921),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2418),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_1731),
.Y(n_2779)
);

CKINVDCx20_ASAP7_75t_R g2780 ( 
.A(n_1930),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_1868),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_1733),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_1934),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_1868),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_1745),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_2548),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_1751),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_1753),
.Y(n_2788)
);

INVxp67_ASAP7_75t_SL g2789 ( 
.A(n_2078),
.Y(n_2789)
);

INVxp67_ASAP7_75t_SL g2790 ( 
.A(n_1946),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_1754),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_1763),
.Y(n_2792)
);

INVxp33_ASAP7_75t_L g2793 ( 
.A(n_2563),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_1766),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_1769),
.Y(n_2795)
);

INVxp67_ASAP7_75t_L g2796 ( 
.A(n_1818),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_2562),
.Y(n_2797)
);

INVxp33_ASAP7_75t_SL g2798 ( 
.A(n_1773),
.Y(n_2798)
);

CKINVDCx20_ASAP7_75t_R g2799 ( 
.A(n_1935),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1770),
.Y(n_2800)
);

CKINVDCx16_ASAP7_75t_R g2801 ( 
.A(n_2137),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_1719),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_1774),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_1778),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_1787),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_1790),
.Y(n_2806)
);

INVxp67_ASAP7_75t_SL g2807 ( 
.A(n_1946),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_1946),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2000),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_1792),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2655),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_1795),
.Y(n_2812)
);

INVxp33_ASAP7_75t_SL g2813 ( 
.A(n_1803),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_1814),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_2660),
.Y(n_2815)
);

HB1xp67_ASAP7_75t_L g2816 ( 
.A(n_1824),
.Y(n_2816)
);

INVxp67_ASAP7_75t_SL g2817 ( 
.A(n_2000),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_1819),
.Y(n_2818)
);

BUFx6f_ASAP7_75t_L g2819 ( 
.A(n_2000),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_1827),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_1832),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_2648),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_1833),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_1839),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_1840),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1841),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_1875),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2060),
.Y(n_2828)
);

NOR2xp33_ASAP7_75t_L g2829 ( 
.A(n_1899),
.B(n_0),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_1842),
.Y(n_2830)
);

CKINVDCx16_ASAP7_75t_R g2831 ( 
.A(n_2137),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_1844),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2060),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_1849),
.Y(n_2834)
);

BUFx6f_ASAP7_75t_L g2835 ( 
.A(n_2060),
.Y(n_2835)
);

INVxp67_ASAP7_75t_SL g2836 ( 
.A(n_2121),
.Y(n_2836)
);

INVxp67_ASAP7_75t_L g2837 ( 
.A(n_2154),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_1855),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_1720),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_1723),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_1859),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_1861),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_1864),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_1866),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_1867),
.Y(n_2845)
);

INVxp67_ASAP7_75t_SL g2846 ( 
.A(n_2121),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_1871),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_1872),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2121),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2656),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_1874),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_2657),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_1880),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_1943),
.Y(n_2854)
);

INVxp67_ASAP7_75t_SL g2855 ( 
.A(n_2126),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_1882),
.Y(n_2856)
);

INVxp67_ASAP7_75t_SL g2857 ( 
.A(n_2126),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_1885),
.Y(n_2858)
);

INVxp67_ASAP7_75t_L g2859 ( 
.A(n_2154),
.Y(n_2859)
);

INVxp67_ASAP7_75t_SL g2860 ( 
.A(n_2390),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2645),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_1894),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_1898),
.Y(n_2863)
);

HB1xp67_ASAP7_75t_L g2864 ( 
.A(n_1904),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_1909),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_1914),
.Y(n_2866)
);

INVxp33_ASAP7_75t_L g2867 ( 
.A(n_1718),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_2654),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_1916),
.Y(n_2869)
);

CKINVDCx16_ASAP7_75t_R g2870 ( 
.A(n_2311),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_1917),
.Y(n_2871)
);

CKINVDCx16_ASAP7_75t_R g2872 ( 
.A(n_2311),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_1924),
.Y(n_2873)
);

INVxp33_ASAP7_75t_SL g2874 ( 
.A(n_1936),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_1926),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_1728),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_1927),
.Y(n_2877)
);

CKINVDCx20_ASAP7_75t_R g2878 ( 
.A(n_1965),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2390),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_1887),
.Y(n_2880)
);

INVxp67_ASAP7_75t_SL g2881 ( 
.A(n_2390),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_1932),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_1933),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_1945),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_1952),
.Y(n_2885)
);

CKINVDCx20_ASAP7_75t_R g2886 ( 
.A(n_1971),
.Y(n_2886)
);

CKINVDCx20_ASAP7_75t_R g2887 ( 
.A(n_1979),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_1953),
.Y(n_2888)
);

HB1xp67_ASAP7_75t_L g2889 ( 
.A(n_1974),
.Y(n_2889)
);

INVxp33_ASAP7_75t_SL g2890 ( 
.A(n_2017),
.Y(n_2890)
);

CKINVDCx5p33_ASAP7_75t_R g2891 ( 
.A(n_1730),
.Y(n_2891)
);

INVxp67_ASAP7_75t_L g2892 ( 
.A(n_2597),
.Y(n_2892)
);

CKINVDCx20_ASAP7_75t_R g2893 ( 
.A(n_1983),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_1967),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_1975),
.Y(n_2895)
);

INVxp33_ASAP7_75t_SL g2896 ( 
.A(n_2182),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_1986),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_1995),
.Y(n_2898)
);

CKINVDCx5p33_ASAP7_75t_R g2899 ( 
.A(n_2649),
.Y(n_2899)
);

CKINVDCx5p33_ASAP7_75t_R g2900 ( 
.A(n_2650),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2002),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2597),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_2670),
.Y(n_2903)
);

INVx5_ASAP7_75t_L g2904 ( 
.A(n_2801),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2725),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2674),
.B(n_1776),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2677),
.B(n_1821),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2687),
.B(n_1831),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2725),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2790),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2807),
.B(n_1905),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2725),
.Y(n_2912)
);

BUFx2_ASAP7_75t_L g2913 ( 
.A(n_2683),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2729),
.Y(n_2914)
);

AND2x4_ASAP7_75t_L g2915 ( 
.A(n_2796),
.B(n_2837),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2729),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2817),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2675),
.Y(n_2918)
);

CKINVDCx20_ASAP7_75t_R g2919 ( 
.A(n_2732),
.Y(n_2919)
);

INVx3_ASAP7_75t_L g2920 ( 
.A(n_2758),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_2859),
.B(n_1737),
.Y(n_2921)
);

HB1xp67_ASAP7_75t_L g2922 ( 
.A(n_2666),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2729),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_2717),
.B(n_2123),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2781),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2781),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2836),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2781),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2846),
.B(n_2855),
.Y(n_2929)
);

OA21x2_ASAP7_75t_L g2930 ( 
.A1(n_2678),
.A2(n_2008),
.B(n_2006),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2819),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2857),
.Y(n_2932)
);

OAI22x1_ASAP7_75t_L g2933 ( 
.A1(n_2827),
.A2(n_2254),
.B1(n_2449),
.B2(n_2365),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2665),
.A2(n_1920),
.B1(n_2312),
.B2(n_1768),
.Y(n_2934)
);

OAI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2671),
.A2(n_2192),
.B1(n_2230),
.B2(n_2226),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2860),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2867),
.B(n_1775),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_L g2938 ( 
.A(n_2819),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2682),
.A2(n_2253),
.B1(n_2285),
.B2(n_2276),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2881),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2819),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2835),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2835),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_L g2944 ( 
.A(n_2769),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_2679),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2690),
.B(n_1915),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2772),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2724),
.B(n_2211),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2692),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2672),
.B(n_1775),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2784),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2694),
.B(n_1956),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2695),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2698),
.B(n_2013),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2691),
.A2(n_2295),
.B1(n_2320),
.B2(n_2306),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2676),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2696),
.Y(n_2957)
);

BUFx3_ASAP7_75t_L g2958 ( 
.A(n_2699),
.Y(n_2958)
);

OAI22xp5_ASAP7_75t_SL g2959 ( 
.A1(n_2745),
.A2(n_2331),
.B1(n_2484),
.B2(n_2314),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2808),
.Y(n_2960)
);

INVxp67_ASAP7_75t_L g2961 ( 
.A(n_2761),
.Y(n_2961)
);

AND2x6_ASAP7_75t_L g2962 ( 
.A(n_2764),
.B(n_2770),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2664),
.Y(n_2963)
);

HB1xp67_ASAP7_75t_L g2964 ( 
.A(n_2681),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2798),
.B(n_2369),
.Y(n_2965)
);

BUFx2_ASAP7_75t_L g2966 ( 
.A(n_2688),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2704),
.B(n_1782),
.Y(n_2967)
);

HB1xp67_ASAP7_75t_L g2968 ( 
.A(n_2706),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2680),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2667),
.Y(n_2970)
);

HB1xp67_ASAP7_75t_L g2971 ( 
.A(n_2709),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2809),
.Y(n_2972)
);

BUFx6f_ASAP7_75t_L g2973 ( 
.A(n_2828),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2684),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2833),
.Y(n_2975)
);

BUFx2_ASAP7_75t_L g2976 ( 
.A(n_2722),
.Y(n_2976)
);

BUFx6f_ASAP7_75t_L g2977 ( 
.A(n_2849),
.Y(n_2977)
);

OAI21xp33_ASAP7_75t_L g2978 ( 
.A1(n_2775),
.A2(n_2330),
.B(n_2322),
.Y(n_2978)
);

INVxp67_ASAP7_75t_L g2979 ( 
.A(n_2816),
.Y(n_2979)
);

CKINVDCx5p33_ASAP7_75t_R g2980 ( 
.A(n_2802),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2879),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2719),
.Y(n_2982)
);

HB1xp67_ASAP7_75t_L g2983 ( 
.A(n_2734),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2701),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_2811),
.Y(n_2985)
);

INVx4_ASAP7_75t_L g2986 ( 
.A(n_2815),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2702),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2713),
.B(n_1782),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2669),
.Y(n_2989)
);

OA22x2_ASAP7_75t_SL g2990 ( 
.A1(n_2789),
.A2(n_2350),
.B1(n_2547),
.B2(n_2022),
.Y(n_2990)
);

AND2x4_ASAP7_75t_L g2991 ( 
.A(n_2892),
.B(n_1749),
.Y(n_2991)
);

OAI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2757),
.A2(n_2333),
.B1(n_2432),
.B2(n_2377),
.Y(n_2992)
);

AND2x4_ASAP7_75t_L g2993 ( 
.A(n_2902),
.B(n_1903),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2735),
.B(n_2001),
.Y(n_2994)
);

BUFx2_ASAP7_75t_L g2995 ( 
.A(n_2773),
.Y(n_2995)
);

HB1xp67_ASAP7_75t_L g2996 ( 
.A(n_2778),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2703),
.Y(n_2997)
);

XNOR2xp5_ASAP7_75t_L g2998 ( 
.A(n_2754),
.B(n_1990),
.Y(n_2998)
);

INVx3_ASAP7_75t_L g2999 ( 
.A(n_2742),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2707),
.B(n_2049),
.Y(n_3000)
);

OAI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2705),
.A2(n_1793),
.B(n_1742),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2712),
.B(n_2053),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2718),
.B(n_2429),
.Y(n_3003)
);

INVx3_ASAP7_75t_L g3004 ( 
.A(n_2771),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2765),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2673),
.A2(n_2007),
.B1(n_2032),
.B2(n_2031),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2708),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2748),
.B(n_1783),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2720),
.B(n_2161),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2774),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2710),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_2767),
.Y(n_3012)
);

INVx3_ASAP7_75t_L g3013 ( 
.A(n_2776),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2714),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2715),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2793),
.B(n_1783),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_SL g3017 ( 
.A1(n_2760),
.A2(n_2044),
.B1(n_2096),
.B2(n_2069),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2721),
.B(n_2225),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2723),
.B(n_2301),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_SL g3020 ( 
.A1(n_2766),
.A2(n_2100),
.B1(n_2143),
.B2(n_2132),
.Y(n_3020)
);

INVx4_ASAP7_75t_L g3021 ( 
.A(n_2822),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2727),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2759),
.B(n_1884),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2728),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2685),
.B(n_1884),
.Y(n_3025)
);

BUFx3_ASAP7_75t_L g3026 ( 
.A(n_2730),
.Y(n_3026)
);

AOI22x1_ASAP7_75t_SL g3027 ( 
.A1(n_2777),
.A2(n_2170),
.B1(n_2171),
.B2(n_2163),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2779),
.Y(n_3028)
);

OAI21x1_ASAP7_75t_L g3029 ( 
.A1(n_2733),
.A2(n_1820),
.B(n_1816),
.Y(n_3029)
);

CKINVDCx6p67_ASAP7_75t_R g3030 ( 
.A(n_2686),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2693),
.B(n_1889),
.Y(n_3031)
);

OA21x2_ASAP7_75t_L g3032 ( 
.A1(n_2737),
.A2(n_2027),
.B(n_2021),
.Y(n_3032)
);

BUFx6f_ASAP7_75t_L g3033 ( 
.A(n_2768),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2739),
.Y(n_3034)
);

INVx6_ASAP7_75t_L g3035 ( 
.A(n_2831),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2741),
.Y(n_3036)
);

AOI22xp5_ASAP7_75t_SL g3037 ( 
.A1(n_2780),
.A2(n_2179),
.B1(n_2237),
.B2(n_2204),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2744),
.Y(n_3038)
);

INVx3_ASAP7_75t_L g3039 ( 
.A(n_2782),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2700),
.A2(n_2487),
.B1(n_2550),
.B2(n_2528),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2746),
.Y(n_3041)
);

BUFx6f_ASAP7_75t_L g3042 ( 
.A(n_2747),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2749),
.Y(n_3043)
);

AND2x4_ASAP7_75t_L g3044 ( 
.A(n_2736),
.B(n_2689),
.Y(n_3044)
);

INVxp33_ASAP7_75t_SL g3045 ( 
.A(n_2786),
.Y(n_3045)
);

INVx6_ASAP7_75t_L g3046 ( 
.A(n_2870),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2750),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2785),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2738),
.B(n_2308),
.Y(n_3049)
);

OA21x2_ASAP7_75t_L g3050 ( 
.A1(n_2751),
.A2(n_2755),
.B(n_2753),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2787),
.Y(n_3051)
);

BUFx6f_ASAP7_75t_L g3052 ( 
.A(n_2756),
.Y(n_3052)
);

INVx5_ASAP7_75t_L g3053 ( 
.A(n_2872),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2762),
.Y(n_3054)
);

INVx3_ASAP7_75t_L g3055 ( 
.A(n_2788),
.Y(n_3055)
);

INVx3_ASAP7_75t_L g3056 ( 
.A(n_2791),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2763),
.Y(n_3057)
);

OA21x2_ASAP7_75t_L g3058 ( 
.A1(n_2740),
.A2(n_2048),
.B(n_2046),
.Y(n_3058)
);

AND2x4_ASAP7_75t_L g3059 ( 
.A(n_2864),
.B(n_2889),
.Y(n_3059)
);

INVxp33_ASAP7_75t_SL g3060 ( 
.A(n_2797),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2792),
.Y(n_3061)
);

OA21x2_ASAP7_75t_L g3062 ( 
.A1(n_2794),
.A2(n_2800),
.B(n_2795),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2803),
.Y(n_3063)
);

AND2x4_ASAP7_75t_L g3064 ( 
.A(n_2839),
.B(n_2016),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2804),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2697),
.B(n_2743),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2805),
.Y(n_3067)
);

AND2x6_ASAP7_75t_L g3068 ( 
.A(n_2806),
.B(n_2033),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2810),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2812),
.Y(n_3070)
);

AOI22x1_ASAP7_75t_SL g3071 ( 
.A1(n_2783),
.A2(n_2364),
.B1(n_2380),
.B2(n_2361),
.Y(n_3071)
);

INVx4_ASAP7_75t_L g3072 ( 
.A(n_2840),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_SL g3073 ( 
.A(n_2711),
.B(n_1806),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2752),
.Y(n_3074)
);

INVx3_ASAP7_75t_L g3075 ( 
.A(n_2814),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2818),
.Y(n_3076)
);

OAI21x1_ASAP7_75t_L g3077 ( 
.A1(n_2820),
.A2(n_1852),
.B(n_1822),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2821),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2823),
.B(n_2442),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2824),
.Y(n_3080)
);

BUFx2_ASAP7_75t_L g3081 ( 
.A(n_2850),
.Y(n_3081)
);

OA21x2_ASAP7_75t_L g3082 ( 
.A1(n_2825),
.A2(n_2068),
.B(n_2054),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2826),
.Y(n_3083)
);

HB1xp67_ASAP7_75t_L g3084 ( 
.A(n_2852),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2830),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2832),
.Y(n_3086)
);

INVx5_ASAP7_75t_L g3087 ( 
.A(n_2668),
.Y(n_3087)
);

OAI21x1_ASAP7_75t_L g3088 ( 
.A1(n_2901),
.A2(n_1856),
.B(n_1854),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2861),
.B(n_1889),
.Y(n_3089)
);

BUFx2_ASAP7_75t_L g3090 ( 
.A(n_2868),
.Y(n_3090)
);

AND2x4_ASAP7_75t_L g3091 ( 
.A(n_2876),
.B(n_2891),
.Y(n_3091)
);

AND2x4_ASAP7_75t_L g3092 ( 
.A(n_2899),
.B(n_2063),
.Y(n_3092)
);

AND2x4_ASAP7_75t_L g3093 ( 
.A(n_2900),
.B(n_2079),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_2834),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2963),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2958),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2970),
.Y(n_3097)
);

INVx2_ASAP7_75t_SL g3098 ( 
.A(n_3066),
.Y(n_3098)
);

HB1xp67_ASAP7_75t_L g3099 ( 
.A(n_2964),
.Y(n_3099)
);

CKINVDCx16_ASAP7_75t_R g3100 ( 
.A(n_2919),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_R g3101 ( 
.A(n_2903),
.B(n_2918),
.Y(n_3101)
);

CKINVDCx20_ASAP7_75t_R g3102 ( 
.A(n_2980),
.Y(n_3102)
);

CKINVDCx5p33_ASAP7_75t_R g3103 ( 
.A(n_2985),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2956),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_2945),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2969),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_3045),
.Y(n_3107)
);

CKINVDCx5p33_ASAP7_75t_R g3108 ( 
.A(n_3060),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_3081),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2974),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_R g3111 ( 
.A(n_3090),
.B(n_2716),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_3030),
.Y(n_3112)
);

CKINVDCx5p33_ASAP7_75t_R g3113 ( 
.A(n_2998),
.Y(n_3113)
);

NAND2xp33_ASAP7_75t_R g3114 ( 
.A(n_2913),
.B(n_2813),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_2966),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2976),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2982),
.Y(n_3117)
);

CKINVDCx5p33_ASAP7_75t_R g3118 ( 
.A(n_2995),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_3035),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2949),
.B(n_2874),
.Y(n_3120)
);

NOR2x1p5_ASAP7_75t_L g3121 ( 
.A(n_2915),
.B(n_2580),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2989),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_3046),
.Y(n_3123)
);

CKINVDCx5p33_ASAP7_75t_R g3124 ( 
.A(n_2986),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_3021),
.Y(n_3125)
);

CKINVDCx5p33_ASAP7_75t_R g3126 ( 
.A(n_3072),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_2937),
.B(n_2726),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_3084),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_2904),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_3053),
.Y(n_3130)
);

CKINVDCx5p33_ASAP7_75t_R g3131 ( 
.A(n_3091),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_2968),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_2920),
.B(n_2838),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_2971),
.Y(n_3134)
);

BUFx2_ASAP7_75t_L g3135 ( 
.A(n_3074),
.Y(n_3135)
);

BUFx3_ASAP7_75t_L g3136 ( 
.A(n_3067),
.Y(n_3136)
);

CKINVDCx5p33_ASAP7_75t_R g3137 ( 
.A(n_2983),
.Y(n_3137)
);

CKINVDCx5p33_ASAP7_75t_R g3138 ( 
.A(n_2996),
.Y(n_3138)
);

CKINVDCx20_ASAP7_75t_R g3139 ( 
.A(n_2922),
.Y(n_3139)
);

CKINVDCx16_ASAP7_75t_R g3140 ( 
.A(n_3073),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2924),
.B(n_2890),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3078),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3083),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3042),
.Y(n_3144)
);

AND2x4_ASAP7_75t_L g3145 ( 
.A(n_3064),
.B(n_3092),
.Y(n_3145)
);

CKINVDCx5p33_ASAP7_75t_R g3146 ( 
.A(n_3017),
.Y(n_3146)
);

CKINVDCx5p33_ASAP7_75t_R g3147 ( 
.A(n_3020),
.Y(n_3147)
);

CKINVDCx5p33_ASAP7_75t_R g3148 ( 
.A(n_3087),
.Y(n_3148)
);

CKINVDCx5p33_ASAP7_75t_R g3149 ( 
.A(n_2959),
.Y(n_3149)
);

CKINVDCx5p33_ASAP7_75t_R g3150 ( 
.A(n_3037),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_3052),
.Y(n_3151)
);

CKINVDCx5p33_ASAP7_75t_R g3152 ( 
.A(n_3027),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_3071),
.Y(n_3153)
);

CKINVDCx5p33_ASAP7_75t_R g3154 ( 
.A(n_2948),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_R g3155 ( 
.A(n_3004),
.B(n_2731),
.Y(n_3155)
);

CKINVDCx5p33_ASAP7_75t_R g3156 ( 
.A(n_2965),
.Y(n_3156)
);

NOR2xp67_ASAP7_75t_L g3157 ( 
.A(n_2961),
.B(n_2841),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2953),
.B(n_2896),
.Y(n_3158)
);

CKINVDCx5p33_ASAP7_75t_R g3159 ( 
.A(n_3023),
.Y(n_3159)
);

CKINVDCx5p33_ASAP7_75t_R g3160 ( 
.A(n_3006),
.Y(n_3160)
);

CKINVDCx5p33_ASAP7_75t_R g3161 ( 
.A(n_3040),
.Y(n_3161)
);

CKINVDCx16_ASAP7_75t_R g3162 ( 
.A(n_2950),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2944),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3036),
.Y(n_3164)
);

CKINVDCx5p33_ASAP7_75t_R g3165 ( 
.A(n_2979),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_R g3166 ( 
.A(n_3010),
.B(n_2799),
.Y(n_3166)
);

CKINVDCx5p33_ASAP7_75t_R g3167 ( 
.A(n_3093),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_R g3168 ( 
.A(n_3013),
.B(n_2854),
.Y(n_3168)
);

AOI21x1_ASAP7_75t_L g3169 ( 
.A1(n_2957),
.A2(n_2843),
.B(n_2842),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_2935),
.Y(n_3170)
);

CKINVDCx20_ASAP7_75t_R g3171 ( 
.A(n_2934),
.Y(n_3171)
);

CKINVDCx5p33_ASAP7_75t_R g3172 ( 
.A(n_2939),
.Y(n_3172)
);

NAND2xp33_ASAP7_75t_R g3173 ( 
.A(n_3059),
.B(n_2829),
.Y(n_3173)
);

CKINVDCx5p33_ASAP7_75t_R g3174 ( 
.A(n_2955),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2947),
.Y(n_3175)
);

CKINVDCx5p33_ASAP7_75t_R g3176 ( 
.A(n_2992),
.Y(n_3176)
);

CKINVDCx5p33_ASAP7_75t_R g3177 ( 
.A(n_3089),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3038),
.Y(n_3178)
);

CKINVDCx5p33_ASAP7_75t_R g3179 ( 
.A(n_3076),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2973),
.Y(n_3180)
);

CKINVDCx5p33_ASAP7_75t_R g3181 ( 
.A(n_3094),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3041),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2929),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3043),
.Y(n_3184)
);

HB1xp67_ASAP7_75t_L g3185 ( 
.A(n_3008),
.Y(n_3185)
);

CKINVDCx5p33_ASAP7_75t_R g3186 ( 
.A(n_2967),
.Y(n_3186)
);

BUFx2_ASAP7_75t_L g3187 ( 
.A(n_3016),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_2988),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3047),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3054),
.Y(n_3190)
);

CKINVDCx5p33_ASAP7_75t_R g3191 ( 
.A(n_3026),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3007),
.B(n_3011),
.Y(n_3192)
);

CKINVDCx5p33_ASAP7_75t_R g3193 ( 
.A(n_3025),
.Y(n_3193)
);

CKINVDCx5p33_ASAP7_75t_R g3194 ( 
.A(n_3031),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3057),
.Y(n_3195)
);

CKINVDCx5p33_ASAP7_75t_R g3196 ( 
.A(n_3068),
.Y(n_3196)
);

NOR2x1_ASAP7_75t_L g3197 ( 
.A(n_3028),
.B(n_2844),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3048),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_3068),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_R g3200 ( 
.A(n_3039),
.B(n_2878),
.Y(n_3200)
);

CKINVDCx5p33_ASAP7_75t_R g3201 ( 
.A(n_2962),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_2962),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3051),
.Y(n_3203)
);

CKINVDCx5p33_ASAP7_75t_R g3204 ( 
.A(n_3055),
.Y(n_3204)
);

CKINVDCx20_ASAP7_75t_R g3205 ( 
.A(n_3003),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_3056),
.Y(n_3206)
);

CKINVDCx20_ASAP7_75t_R g3207 ( 
.A(n_3058),
.Y(n_3207)
);

CKINVDCx5p33_ASAP7_75t_R g3208 ( 
.A(n_3075),
.Y(n_3208)
);

CKINVDCx5p33_ASAP7_75t_R g3209 ( 
.A(n_3086),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_R g3210 ( 
.A(n_2910),
.B(n_2886),
.Y(n_3210)
);

CKINVDCx20_ASAP7_75t_R g3211 ( 
.A(n_2946),
.Y(n_3211)
);

AND2x6_ASAP7_75t_L g3212 ( 
.A(n_3061),
.B(n_2845),
.Y(n_3212)
);

HB1xp67_ASAP7_75t_L g3213 ( 
.A(n_2994),
.Y(n_3213)
);

HB1xp67_ASAP7_75t_SL g3214 ( 
.A(n_2933),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3063),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3065),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_2917),
.Y(n_3217)
);

CKINVDCx5p33_ASAP7_75t_R g3218 ( 
.A(n_2927),
.Y(n_3218)
);

CKINVDCx5p33_ASAP7_75t_R g3219 ( 
.A(n_2932),
.Y(n_3219)
);

CKINVDCx5p33_ASAP7_75t_R g3220 ( 
.A(n_2936),
.Y(n_3220)
);

AOI21x1_ASAP7_75t_L g3221 ( 
.A1(n_3014),
.A2(n_2848),
.B(n_2847),
.Y(n_3221)
);

INVx3_ASAP7_75t_L g3222 ( 
.A(n_2930),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_2940),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3069),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_R g3225 ( 
.A(n_3070),
.B(n_2887),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2975),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3015),
.B(n_2851),
.Y(n_3227)
);

CKINVDCx5p33_ASAP7_75t_R g3228 ( 
.A(n_2921),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_2991),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_2993),
.Y(n_3230)
);

CKINVDCx5p33_ASAP7_75t_R g3231 ( 
.A(n_3005),
.Y(n_3231)
);

OAI22xp33_ASAP7_75t_SL g3232 ( 
.A1(n_2952),
.A2(n_2583),
.B1(n_2633),
.B2(n_2625),
.Y(n_3232)
);

CKINVDCx5p33_ASAP7_75t_R g3233 ( 
.A(n_3012),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2977),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_3033),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2951),
.Y(n_3236)
);

AO22x2_ASAP7_75t_L g3237 ( 
.A1(n_2990),
.A2(n_2880),
.B1(n_2505),
.B2(n_1746),
.Y(n_3237)
);

CKINVDCx5p33_ASAP7_75t_R g3238 ( 
.A(n_3080),
.Y(n_3238)
);

CKINVDCx5p33_ASAP7_75t_R g3239 ( 
.A(n_3085),
.Y(n_3239)
);

CKINVDCx20_ASAP7_75t_R g3240 ( 
.A(n_2954),
.Y(n_3240)
);

CKINVDCx20_ASAP7_75t_R g3241 ( 
.A(n_3000),
.Y(n_3241)
);

CKINVDCx5p33_ASAP7_75t_R g3242 ( 
.A(n_3002),
.Y(n_3242)
);

CKINVDCx5p33_ASAP7_75t_R g3243 ( 
.A(n_3009),
.Y(n_3243)
);

INVxp67_ASAP7_75t_SL g3244 ( 
.A(n_2911),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3022),
.Y(n_3245)
);

CKINVDCx5p33_ASAP7_75t_R g3246 ( 
.A(n_3018),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3034),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_R g3248 ( 
.A(n_2999),
.B(n_2893),
.Y(n_3248)
);

CKINVDCx5p33_ASAP7_75t_R g3249 ( 
.A(n_3019),
.Y(n_3249)
);

CKINVDCx5p33_ASAP7_75t_R g3250 ( 
.A(n_3049),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_R g3251 ( 
.A(n_2906),
.B(n_2853),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2984),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2960),
.Y(n_3253)
);

CKINVDCx5p33_ASAP7_75t_R g3254 ( 
.A(n_2978),
.Y(n_3254)
);

CKINVDCx5p33_ASAP7_75t_R g3255 ( 
.A(n_2987),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_3062),
.Y(n_3256)
);

CKINVDCx5p33_ASAP7_75t_R g3257 ( 
.A(n_2997),
.Y(n_3257)
);

INVxp67_ASAP7_75t_L g3258 ( 
.A(n_2907),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2972),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3024),
.B(n_2856),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2981),
.Y(n_3261)
);

HB1xp67_ASAP7_75t_L g3262 ( 
.A(n_3050),
.Y(n_3262)
);

BUFx2_ASAP7_75t_L g3263 ( 
.A(n_3082),
.Y(n_3263)
);

BUFx3_ASAP7_75t_L g3264 ( 
.A(n_3032),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3077),
.Y(n_3265)
);

CKINVDCx20_ASAP7_75t_R g3266 ( 
.A(n_2908),
.Y(n_3266)
);

CKINVDCx20_ASAP7_75t_R g3267 ( 
.A(n_3079),
.Y(n_3267)
);

CKINVDCx5p33_ASAP7_75t_R g3268 ( 
.A(n_2925),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3088),
.Y(n_3269)
);

NAND2xp33_ASAP7_75t_R g3270 ( 
.A(n_3001),
.B(n_2634),
.Y(n_3270)
);

CKINVDCx5p33_ASAP7_75t_R g3271 ( 
.A(n_2938),
.Y(n_3271)
);

HB1xp67_ASAP7_75t_L g3272 ( 
.A(n_3029),
.Y(n_3272)
);

CKINVDCx20_ASAP7_75t_R g3273 ( 
.A(n_2905),
.Y(n_3273)
);

CKINVDCx5p33_ASAP7_75t_R g3274 ( 
.A(n_2909),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2912),
.Y(n_3275)
);

CKINVDCx5p33_ASAP7_75t_R g3276 ( 
.A(n_2914),
.Y(n_3276)
);

CKINVDCx5p33_ASAP7_75t_R g3277 ( 
.A(n_2916),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_2923),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_2926),
.Y(n_3279)
);

CKINVDCx5p33_ASAP7_75t_R g3280 ( 
.A(n_2928),
.Y(n_3280)
);

CKINVDCx20_ASAP7_75t_R g3281 ( 
.A(n_2931),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_2941),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2942),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_R g3284 ( 
.A(n_2943),
.B(n_2858),
.Y(n_3284)
);

OR2x2_ASAP7_75t_L g3285 ( 
.A(n_3044),
.B(n_2862),
.Y(n_3285)
);

OAI21x1_ASAP7_75t_L g3286 ( 
.A1(n_3001),
.A2(n_2865),
.B(n_2863),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2956),
.Y(n_3287)
);

HB1xp67_ASAP7_75t_L g3288 ( 
.A(n_2964),
.Y(n_3288)
);

INVx3_ASAP7_75t_L g3289 ( 
.A(n_2958),
.Y(n_3289)
);

BUFx2_ASAP7_75t_L g3290 ( 
.A(n_3066),
.Y(n_3290)
);

BUFx3_ASAP7_75t_L g3291 ( 
.A(n_2920),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_2980),
.Y(n_3292)
);

CKINVDCx5p33_ASAP7_75t_R g3293 ( 
.A(n_2980),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_2956),
.Y(n_3294)
);

CKINVDCx20_ASAP7_75t_R g3295 ( 
.A(n_2919),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_2980),
.Y(n_3296)
);

CKINVDCx20_ASAP7_75t_R g3297 ( 
.A(n_2919),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3286),
.Y(n_3298)
);

CKINVDCx20_ASAP7_75t_R g3299 ( 
.A(n_3102),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3290),
.B(n_2405),
.Y(n_3300)
);

AND2x6_ASAP7_75t_L g3301 ( 
.A(n_3145),
.B(n_3127),
.Y(n_3301)
);

INVx5_ASAP7_75t_L g3302 ( 
.A(n_3145),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3169),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3124),
.B(n_1732),
.Y(n_3304)
);

INVx2_ASAP7_75t_SL g3305 ( 
.A(n_3119),
.Y(n_3305)
);

AND2x4_ASAP7_75t_L g3306 ( 
.A(n_3123),
.B(n_2866),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3221),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_3154),
.B(n_1734),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3244),
.B(n_2459),
.Y(n_3309)
);

INVx2_ASAP7_75t_SL g3310 ( 
.A(n_3135),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3104),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3183),
.B(n_2460),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_3099),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3106),
.Y(n_3314)
);

INVx5_ASAP7_75t_L g3315 ( 
.A(n_3100),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3245),
.Y(n_3316)
);

BUFx2_ASAP7_75t_L g3317 ( 
.A(n_3295),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3247),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_3263),
.A2(n_3256),
.B1(n_3254),
.B2(n_3212),
.Y(n_3319)
);

BUFx10_ASAP7_75t_L g3320 ( 
.A(n_3103),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3242),
.B(n_2502),
.Y(n_3321)
);

INVx1_ASAP7_75t_SL g3322 ( 
.A(n_3297),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3110),
.Y(n_3323)
);

OR2x6_ASAP7_75t_L g3324 ( 
.A(n_3098),
.B(n_2293),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_L g3325 ( 
.A(n_3136),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3243),
.B(n_2557),
.Y(n_3326)
);

BUFx6f_ASAP7_75t_L g3327 ( 
.A(n_3291),
.Y(n_3327)
);

BUFx6f_ASAP7_75t_L g3328 ( 
.A(n_3268),
.Y(n_3328)
);

BUFx6f_ASAP7_75t_L g3329 ( 
.A(n_3271),
.Y(n_3329)
);

AND2x4_ASAP7_75t_L g3330 ( 
.A(n_3105),
.B(n_3292),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_3125),
.B(n_1735),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3198),
.Y(n_3332)
);

CKINVDCx5p33_ASAP7_75t_R g3333 ( 
.A(n_3101),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3117),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3246),
.B(n_2567),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3287),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3294),
.Y(n_3337)
);

AND2x6_ASAP7_75t_L g3338 ( 
.A(n_3120),
.B(n_2869),
.Y(n_3338)
);

CKINVDCx20_ASAP7_75t_R g3339 ( 
.A(n_3293),
.Y(n_3339)
);

NOR2x1p5_ASAP7_75t_L g3340 ( 
.A(n_3107),
.B(n_2871),
.Y(n_3340)
);

BUFx2_ASAP7_75t_L g3341 ( 
.A(n_3139),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_3133),
.Y(n_3342)
);

INVx3_ASAP7_75t_R g3343 ( 
.A(n_3285),
.Y(n_3343)
);

NAND3xp33_ASAP7_75t_L g3344 ( 
.A(n_3156),
.B(n_2643),
.C(n_2642),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3203),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3187),
.B(n_2408),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3165),
.B(n_2414),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3249),
.B(n_2589),
.Y(n_3348)
);

INVx2_ASAP7_75t_SL g3349 ( 
.A(n_3248),
.Y(n_3349)
);

AND2x6_ASAP7_75t_L g3350 ( 
.A(n_3158),
.B(n_2873),
.Y(n_3350)
);

OR2x2_ASAP7_75t_L g3351 ( 
.A(n_3288),
.B(n_1835),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_3126),
.B(n_3191),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3215),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3142),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_L g3355 ( 
.A1(n_3212),
.A2(n_2438),
.B1(n_2439),
.B2(n_2421),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3250),
.B(n_2593),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3143),
.Y(n_3357)
);

AND2x4_ASAP7_75t_L g3358 ( 
.A(n_3296),
.B(n_2875),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3216),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3224),
.Y(n_3360)
);

AND2x6_ASAP7_75t_L g3361 ( 
.A(n_3144),
.B(n_2877),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3193),
.B(n_2467),
.Y(n_3362)
);

INVx3_ASAP7_75t_L g3363 ( 
.A(n_3181),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3164),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_3141),
.B(n_1836),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3194),
.B(n_2479),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3258),
.B(n_3096),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3096),
.B(n_2647),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3185),
.B(n_2499),
.Y(n_3369)
);

INVx3_ASAP7_75t_L g3370 ( 
.A(n_3231),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3178),
.Y(n_3371)
);

HB1xp67_ASAP7_75t_L g3372 ( 
.A(n_3166),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_3204),
.B(n_1740),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3182),
.Y(n_3374)
);

CKINVDCx5p33_ASAP7_75t_R g3375 ( 
.A(n_3108),
.Y(n_3375)
);

AND2x4_ASAP7_75t_L g3376 ( 
.A(n_3115),
.B(n_2882),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_3116),
.B(n_2883),
.Y(n_3377)
);

OAI22x1_ASAP7_75t_L g3378 ( 
.A1(n_3161),
.A2(n_1881),
.B1(n_1907),
.B2(n_1863),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3184),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3095),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3097),
.Y(n_3381)
);

AND2x2_ASAP7_75t_SL g3382 ( 
.A(n_3140),
.B(n_1876),
.Y(n_3382)
);

AO21x2_ASAP7_75t_L g3383 ( 
.A1(n_3262),
.A2(n_2885),
.B(n_2884),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3189),
.Y(n_3384)
);

INVx3_ASAP7_75t_L g3385 ( 
.A(n_3233),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3122),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_3170),
.B(n_3172),
.Y(n_3387)
);

AND2x2_ASAP7_75t_SL g3388 ( 
.A(n_3162),
.B(n_1928),
.Y(n_3388)
);

BUFx4f_ASAP7_75t_L g3389 ( 
.A(n_3151),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_3174),
.B(n_2019),
.Y(n_3390)
);

CKINVDCx20_ASAP7_75t_R g3391 ( 
.A(n_3109),
.Y(n_3391)
);

AND2x2_ASAP7_75t_SL g3392 ( 
.A(n_3213),
.B(n_1947),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3190),
.Y(n_3393)
);

AND2x4_ASAP7_75t_L g3394 ( 
.A(n_3118),
.B(n_3112),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3176),
.B(n_2020),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_3211),
.B(n_2056),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3195),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3206),
.B(n_1741),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_SL g3399 ( 
.A(n_3208),
.B(n_1743),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_3235),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3209),
.B(n_3238),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3252),
.Y(n_3402)
);

BUFx10_ASAP7_75t_L g3403 ( 
.A(n_3129),
.Y(n_3403)
);

BUFx3_ASAP7_75t_L g3404 ( 
.A(n_3273),
.Y(n_3404)
);

INVx4_ASAP7_75t_L g3405 ( 
.A(n_3131),
.Y(n_3405)
);

CKINVDCx16_ASAP7_75t_R g3406 ( 
.A(n_3111),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3236),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3128),
.B(n_2523),
.Y(n_3408)
);

BUFx6f_ASAP7_75t_L g3409 ( 
.A(n_3163),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_3240),
.B(n_2138),
.Y(n_3410)
);

INVx6_ASAP7_75t_L g3411 ( 
.A(n_3121),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_SL g3412 ( 
.A(n_3239),
.B(n_1744),
.Y(n_3412)
);

AOI21x1_ASAP7_75t_L g3413 ( 
.A1(n_3272),
.A2(n_2894),
.B(n_2888),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3241),
.B(n_2146),
.Y(n_3414)
);

INVx4_ASAP7_75t_L g3415 ( 
.A(n_3130),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3289),
.B(n_2498),
.Y(n_3416)
);

INVx3_ASAP7_75t_L g3417 ( 
.A(n_3167),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3260),
.Y(n_3418)
);

AO22x2_ASAP7_75t_L g3419 ( 
.A1(n_3171),
.A2(n_2164),
.B1(n_2176),
.B2(n_2156),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_3157),
.B(n_1747),
.Y(n_3420)
);

BUFx2_ASAP7_75t_L g3421 ( 
.A(n_3168),
.Y(n_3421)
);

AND2x6_ASAP7_75t_L g3422 ( 
.A(n_3197),
.B(n_2895),
.Y(n_3422)
);

OR2x2_ASAP7_75t_SL g3423 ( 
.A(n_3114),
.B(n_2558),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3192),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3132),
.B(n_2574),
.Y(n_3425)
);

INVx6_ASAP7_75t_L g3426 ( 
.A(n_3148),
.Y(n_3426)
);

INVx3_ASAP7_75t_L g3427 ( 
.A(n_3175),
.Y(n_3427)
);

BUFx3_ASAP7_75t_L g3428 ( 
.A(n_3281),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3253),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3134),
.B(n_2588),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3259),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3261),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3255),
.B(n_2498),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3266),
.B(n_2190),
.Y(n_3434)
);

AND2x6_ASAP7_75t_L g3435 ( 
.A(n_3180),
.B(n_3226),
.Y(n_3435)
);

BUFx6f_ASAP7_75t_L g3436 ( 
.A(n_3234),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3228),
.B(n_3229),
.Y(n_3437)
);

INVx4_ASAP7_75t_L g3438 ( 
.A(n_3137),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3282),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3227),
.Y(n_3440)
);

BUFx4f_ASAP7_75t_L g3441 ( 
.A(n_3212),
.Y(n_3441)
);

BUFx2_ASAP7_75t_L g3442 ( 
.A(n_3200),
.Y(n_3442)
);

INVxp67_ASAP7_75t_L g3443 ( 
.A(n_3173),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3264),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3138),
.B(n_2591),
.Y(n_3445)
);

AND2x4_ASAP7_75t_L g3446 ( 
.A(n_3230),
.B(n_2897),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_3212),
.A2(n_2610),
.B1(n_2606),
.B2(n_2304),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3217),
.B(n_2299),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3218),
.B(n_2362),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3257),
.B(n_2517),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3275),
.Y(n_3451)
);

CKINVDCx5p33_ASAP7_75t_R g3452 ( 
.A(n_3113),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3186),
.B(n_2898),
.Y(n_3453)
);

BUFx3_ASAP7_75t_L g3454 ( 
.A(n_3274),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_3225),
.Y(n_3455)
);

INVx3_ASAP7_75t_L g3456 ( 
.A(n_3201),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3283),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3219),
.B(n_2363),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_3220),
.B(n_2366),
.Y(n_3459)
);

AND3x4_ASAP7_75t_L g3460 ( 
.A(n_3177),
.B(n_2099),
.C(n_2090),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3205),
.B(n_2117),
.Y(n_3461)
);

AND2x2_ASAP7_75t_L g3462 ( 
.A(n_3188),
.B(n_1919),
.Y(n_3462)
);

INVx3_ASAP7_75t_L g3463 ( 
.A(n_3202),
.Y(n_3463)
);

BUFx3_ASAP7_75t_L g3464 ( 
.A(n_3276),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3265),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3269),
.Y(n_3466)
);

AND3x2_ASAP7_75t_L g3467 ( 
.A(n_3155),
.B(n_2535),
.C(n_2004),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3196),
.B(n_1748),
.Y(n_3468)
);

NAND2xp33_ASAP7_75t_L g3469 ( 
.A(n_3199),
.B(n_1750),
.Y(n_3469)
);

INVxp67_ASAP7_75t_L g3470 ( 
.A(n_3159),
.Y(n_3470)
);

BUFx6f_ASAP7_75t_L g3471 ( 
.A(n_3277),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_3278),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_3210),
.Y(n_3473)
);

INVx2_ASAP7_75t_SL g3474 ( 
.A(n_3284),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3222),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3223),
.A2(n_1755),
.B1(n_1756),
.B2(n_1752),
.Y(n_3476)
);

OR2x2_ASAP7_75t_L g3477 ( 
.A(n_3160),
.B(n_2371),
.Y(n_3477)
);

AOI22xp5_ASAP7_75t_L g3478 ( 
.A1(n_3267),
.A2(n_2457),
.B1(n_2518),
.B2(n_2391),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3222),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_SL g3480 ( 
.A(n_3146),
.B(n_2556),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3279),
.Y(n_3481)
);

BUFx6f_ASAP7_75t_L g3482 ( 
.A(n_3280),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3207),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3251),
.B(n_1919),
.Y(n_3484)
);

INVx4_ASAP7_75t_SL g3485 ( 
.A(n_3214),
.Y(n_3485)
);

OR2x2_ASAP7_75t_SL g3486 ( 
.A(n_3147),
.B(n_1962),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3232),
.Y(n_3487)
);

INVxp67_ASAP7_75t_L g3488 ( 
.A(n_3270),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3237),
.Y(n_3489)
);

BUFx6f_ASAP7_75t_L g3490 ( 
.A(n_3150),
.Y(n_3490)
);

AND2x4_ASAP7_75t_L g3491 ( 
.A(n_3149),
.B(n_2217),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_3152),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3153),
.Y(n_3493)
);

CKINVDCx5p33_ASAP7_75t_R g3494 ( 
.A(n_3101),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3104),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3104),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3286),
.Y(n_3497)
);

HB1xp67_ASAP7_75t_L g3498 ( 
.A(n_3135),
.Y(n_3498)
);

INVx4_ASAP7_75t_SL g3499 ( 
.A(n_3145),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3244),
.B(n_2600),
.Y(n_3500)
);

INVx1_ASAP7_75t_SL g3501 ( 
.A(n_3297),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3104),
.Y(n_3502)
);

NAND2xp33_ASAP7_75t_L g3503 ( 
.A(n_3124),
.B(n_1760),
.Y(n_3503)
);

BUFx3_ASAP7_75t_L g3504 ( 
.A(n_3119),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3286),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3286),
.Y(n_3506)
);

BUFx3_ASAP7_75t_L g3507 ( 
.A(n_3119),
.Y(n_3507)
);

INVx4_ASAP7_75t_L g3508 ( 
.A(n_3119),
.Y(n_3508)
);

BUFx6f_ASAP7_75t_L g3509 ( 
.A(n_3119),
.Y(n_3509)
);

BUFx6f_ASAP7_75t_L g3510 ( 
.A(n_3119),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3104),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3290),
.B(n_2124),
.Y(n_3512)
);

INVx3_ASAP7_75t_L g3513 ( 
.A(n_3179),
.Y(n_3513)
);

AOI22xp5_ASAP7_75t_L g3514 ( 
.A1(n_3242),
.A2(n_2641),
.B1(n_2638),
.B2(n_1761),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3244),
.B(n_2600),
.Y(n_3515)
);

AND2x4_ASAP7_75t_L g3516 ( 
.A(n_3119),
.B(n_2319),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3286),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3244),
.B(n_2624),
.Y(n_3518)
);

AND2x4_ASAP7_75t_L g3519 ( 
.A(n_3119),
.B(n_2401),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3286),
.Y(n_3520)
);

CKINVDCx20_ASAP7_75t_R g3521 ( 
.A(n_3102),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3154),
.B(n_1762),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_3154),
.B(n_1764),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_SL g3524 ( 
.A(n_3124),
.B(n_1765),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3104),
.Y(n_3525)
);

BUFx2_ASAP7_75t_L g3526 ( 
.A(n_3295),
.Y(n_3526)
);

AND2x4_ASAP7_75t_L g3527 ( 
.A(n_3119),
.B(n_2407),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3290),
.B(n_2124),
.Y(n_3528)
);

INVx4_ASAP7_75t_L g3529 ( 
.A(n_3119),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_3154),
.B(n_1767),
.Y(n_3530)
);

AND2x2_ASAP7_75t_SL g3531 ( 
.A(n_3140),
.B(n_2010),
.Y(n_3531)
);

AND2x4_ASAP7_75t_SL g3532 ( 
.A(n_3102),
.B(n_2129),
.Y(n_3532)
);

AND2x4_ASAP7_75t_L g3533 ( 
.A(n_3119),
.B(n_2420),
.Y(n_3533)
);

CKINVDCx5p33_ASAP7_75t_R g3534 ( 
.A(n_3101),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3135),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_L g3536 ( 
.A(n_3154),
.B(n_1771),
.Y(n_3536)
);

INVx1_ASAP7_75t_SL g3537 ( 
.A(n_3297),
.Y(n_3537)
);

INVx4_ASAP7_75t_L g3538 ( 
.A(n_3119),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3104),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_L g3540 ( 
.A(n_3154),
.B(n_1772),
.Y(n_3540)
);

HB1xp67_ASAP7_75t_L g3541 ( 
.A(n_3135),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3104),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3104),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3244),
.B(n_2624),
.Y(n_3544)
);

INVx3_ASAP7_75t_L g3545 ( 
.A(n_3179),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3367),
.B(n_1777),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3358),
.B(n_1780),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3311),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3424),
.B(n_2071),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3440),
.B(n_2076),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3314),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3316),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3323),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3318),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3298),
.A2(n_2088),
.B(n_2087),
.Y(n_3555)
);

INVx3_ASAP7_75t_L g3556 ( 
.A(n_3504),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_L g3557 ( 
.A1(n_3390),
.A2(n_2349),
.B1(n_2139),
.B2(n_2147),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3448),
.B(n_2098),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_L g3559 ( 
.A(n_3395),
.B(n_1781),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3449),
.B(n_2104),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3334),
.Y(n_3561)
);

INVx2_ASAP7_75t_SL g3562 ( 
.A(n_3302),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3458),
.B(n_2110),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_3443),
.B(n_1784),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3459),
.B(n_2113),
.Y(n_3565)
);

NOR2xp67_ASAP7_75t_L g3566 ( 
.A(n_3508),
.B(n_1786),
.Y(n_3566)
);

AOI22xp5_ASAP7_75t_L g3567 ( 
.A1(n_3522),
.A2(n_1789),
.B1(n_1791),
.B2(n_1788),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3418),
.B(n_2115),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3523),
.B(n_2127),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3453),
.B(n_3387),
.Y(n_3570)
);

NOR2xp33_ASAP7_75t_L g3571 ( 
.A(n_3530),
.B(n_1796),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3536),
.B(n_2128),
.Y(n_3572)
);

OR2x6_ASAP7_75t_L g3573 ( 
.A(n_3509),
.B(n_3510),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3355),
.A2(n_2139),
.B1(n_2147),
.B2(n_2129),
.Y(n_3574)
);

AND2x2_ASAP7_75t_SL g3575 ( 
.A(n_3406),
.B(n_2043),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3310),
.B(n_1798),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3540),
.B(n_3338),
.Y(n_3577)
);

NAND2x1_ASAP7_75t_L g3578 ( 
.A(n_3465),
.B(n_2135),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3336),
.Y(n_3579)
);

NAND2xp33_ASAP7_75t_L g3580 ( 
.A(n_3333),
.B(n_1800),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3332),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3302),
.B(n_1801),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3350),
.B(n_2136),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3345),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3353),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3359),
.B(n_2149),
.Y(n_3586)
);

BUFx3_ASAP7_75t_L g3587 ( 
.A(n_3507),
.Y(n_3587)
);

INVx8_ASAP7_75t_L g3588 ( 
.A(n_3509),
.Y(n_3588)
);

NOR2xp67_ASAP7_75t_L g3589 ( 
.A(n_3529),
.B(n_1804),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3360),
.B(n_2153),
.Y(n_3590)
);

NAND2xp33_ASAP7_75t_L g3591 ( 
.A(n_3494),
.B(n_1805),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3337),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_3342),
.B(n_1807),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_SL g3594 ( 
.A(n_3534),
.B(n_2151),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3380),
.B(n_3381),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3510),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_3342),
.B(n_1808),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3495),
.Y(n_3598)
);

AOI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3365),
.A2(n_1810),
.B1(n_1811),
.B2(n_1809),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3496),
.Y(n_3600)
);

NAND2xp33_ASAP7_75t_SL g3601 ( 
.A(n_3538),
.B(n_1812),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3347),
.B(n_2151),
.Y(n_3602)
);

AND2x4_ASAP7_75t_L g3603 ( 
.A(n_3499),
.B(n_2178),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_3535),
.B(n_1813),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3502),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3511),
.Y(n_3606)
);

OAI22xp33_ASAP7_75t_L g3607 ( 
.A1(n_3447),
.A2(n_1817),
.B1(n_1823),
.B2(n_1815),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3386),
.Y(n_3608)
);

NAND3xp33_ASAP7_75t_L g3609 ( 
.A(n_3375),
.B(n_1826),
.C(n_1825),
.Y(n_3609)
);

INVxp67_ASAP7_75t_L g3610 ( 
.A(n_3541),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_3441),
.B(n_1828),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3525),
.Y(n_3612)
);

INVx2_ASAP7_75t_SL g3613 ( 
.A(n_3404),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3539),
.Y(n_3614)
);

OAI221xp5_ASAP7_75t_L g3615 ( 
.A1(n_3514),
.A2(n_2205),
.B1(n_2206),
.B2(n_2198),
.C(n_2195),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3542),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_3438),
.B(n_1829),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3354),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3488),
.B(n_2208),
.Y(n_3619)
);

INVxp67_ASAP7_75t_SL g3620 ( 
.A(n_3444),
.Y(n_3620)
);

HB1xp67_ASAP7_75t_L g3621 ( 
.A(n_3313),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3484),
.B(n_2209),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_3470),
.B(n_1830),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3312),
.B(n_2214),
.Y(n_3624)
);

O2A1O1Ixp5_ASAP7_75t_L g3625 ( 
.A1(n_3420),
.A2(n_2064),
.B(n_2066),
.C(n_2051),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_L g3626 ( 
.A(n_3477),
.B(n_1834),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3543),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3357),
.Y(n_3628)
);

BUFx6f_ASAP7_75t_L g3629 ( 
.A(n_3328),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3376),
.B(n_1837),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3364),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3309),
.B(n_2215),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3321),
.B(n_3326),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3335),
.B(n_2220),
.Y(n_3634)
);

OR2x2_ASAP7_75t_L g3635 ( 
.A(n_3322),
.B(n_2519),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3348),
.B(n_2221),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3356),
.B(n_2240),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_3339),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3422),
.B(n_2252),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3422),
.B(n_2260),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_SL g3641 ( 
.A(n_3377),
.B(n_1838),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3371),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3374),
.Y(n_3643)
);

INVx2_ASAP7_75t_SL g3644 ( 
.A(n_3428),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3379),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3384),
.Y(n_3646)
);

NAND2xp33_ASAP7_75t_L g3647 ( 
.A(n_3466),
.B(n_1843),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_SL g3648 ( 
.A(n_3330),
.B(n_1845),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3393),
.Y(n_3649)
);

INVx2_ASAP7_75t_SL g3650 ( 
.A(n_3317),
.Y(n_3650)
);

AOI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3301),
.A2(n_1847),
.B1(n_1850),
.B2(n_1846),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3397),
.Y(n_3652)
);

INVx4_ASAP7_75t_L g3653 ( 
.A(n_3328),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_3306),
.B(n_1851),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3362),
.B(n_1853),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3402),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3408),
.B(n_2159),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3451),
.Y(n_3658)
);

BUFx6f_ASAP7_75t_L g3659 ( 
.A(n_3329),
.Y(n_3659)
);

INVxp33_ASAP7_75t_L g3660 ( 
.A(n_3396),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3497),
.A2(n_2266),
.B(n_2263),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3433),
.B(n_3450),
.Y(n_3662)
);

AOI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_3301),
.A2(n_1858),
.B1(n_1860),
.B2(n_1857),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3366),
.B(n_1865),
.Y(n_3664)
);

NOR2xp33_ASAP7_75t_R g3665 ( 
.A(n_3299),
.B(n_1870),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3457),
.Y(n_3666)
);

BUFx3_ASAP7_75t_L g3667 ( 
.A(n_3521),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_3425),
.B(n_1877),
.Y(n_3668)
);

BUFx6f_ASAP7_75t_L g3669 ( 
.A(n_3329),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_L g3670 ( 
.A1(n_3487),
.A2(n_2229),
.B1(n_2241),
.B2(n_2159),
.Y(n_3670)
);

BUFx8_ASAP7_75t_L g3671 ( 
.A(n_3341),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3429),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3325),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3431),
.Y(n_3674)
);

OAI221xp5_ASAP7_75t_L g3675 ( 
.A1(n_3480),
.A2(n_2272),
.B1(n_2278),
.B2(n_2270),
.C(n_2267),
.Y(n_3675)
);

AOI22xp33_ASAP7_75t_L g3676 ( 
.A1(n_3392),
.A2(n_2241),
.B1(n_2268),
.B2(n_2229),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3474),
.B(n_2281),
.Y(n_3677)
);

INVx2_ASAP7_75t_SL g3678 ( 
.A(n_3526),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3407),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_SL g3680 ( 
.A(n_3320),
.B(n_1878),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3512),
.B(n_2283),
.Y(n_3681)
);

NOR2xp33_ASAP7_75t_L g3682 ( 
.A(n_3430),
.B(n_1879),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3432),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3475),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3528),
.B(n_3503),
.Y(n_3685)
);

O2A1O1Ixp5_ASAP7_75t_L g3686 ( 
.A1(n_3413),
.A2(n_2122),
.B(n_2133),
.C(n_2114),
.Y(n_3686)
);

AOI22xp33_ASAP7_75t_L g3687 ( 
.A1(n_3388),
.A2(n_2269),
.B1(n_2287),
.B2(n_2268),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3479),
.Y(n_3688)
);

CKINVDCx5p33_ASAP7_75t_R g3689 ( 
.A(n_3391),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3439),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3319),
.B(n_2305),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3481),
.B(n_2318),
.Y(n_3692)
);

HB1xp67_ASAP7_75t_L g3693 ( 
.A(n_3501),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3303),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3500),
.B(n_2323),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3445),
.B(n_1886),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3401),
.B(n_1888),
.Y(n_3697)
);

OAI22xp5_ASAP7_75t_SL g3698 ( 
.A1(n_3460),
.A2(n_1891),
.B1(n_1895),
.B2(n_1890),
.Y(n_3698)
);

NAND2x1_ASAP7_75t_L g3699 ( 
.A(n_3307),
.B(n_2324),
.Y(n_3699)
);

OR2x2_ASAP7_75t_L g3700 ( 
.A(n_3537),
.B(n_2533),
.Y(n_3700)
);

CKINVDCx20_ASAP7_75t_R g3701 ( 
.A(n_3452),
.Y(n_3701)
);

AOI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3352),
.A2(n_3340),
.B1(n_3412),
.B2(n_3469),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3515),
.B(n_2332),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3518),
.B(n_2334),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3300),
.B(n_2292),
.Y(n_3705)
);

NAND2xp33_ASAP7_75t_L g3706 ( 
.A(n_3305),
.B(n_1896),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3544),
.B(n_2336),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3368),
.B(n_2341),
.Y(n_3708)
);

CKINVDCx5p33_ASAP7_75t_R g3709 ( 
.A(n_3473),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_L g3710 ( 
.A(n_3410),
.B(n_1897),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3446),
.B(n_3456),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3463),
.B(n_2344),
.Y(n_3712)
);

BUFx6f_ASAP7_75t_L g3713 ( 
.A(n_3325),
.Y(n_3713)
);

NOR2xp33_ASAP7_75t_SL g3714 ( 
.A(n_3405),
.B(n_2315),
.Y(n_3714)
);

NOR2xp33_ASAP7_75t_L g3715 ( 
.A(n_3414),
.B(n_1900),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3462),
.B(n_2353),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3434),
.B(n_3361),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3416),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_SL g3719 ( 
.A(n_3363),
.B(n_3370),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3383),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3505),
.A2(n_2359),
.B(n_2356),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3385),
.B(n_1901),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3361),
.B(n_2360),
.Y(n_3723)
);

INVxp67_ASAP7_75t_L g3724 ( 
.A(n_3421),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3491),
.B(n_2368),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3351),
.B(n_2370),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3427),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3454),
.B(n_2374),
.Y(n_3728)
);

NOR2xp67_ASAP7_75t_L g3729 ( 
.A(n_3315),
.B(n_1906),
.Y(n_3729)
);

INVx2_ASAP7_75t_SL g3730 ( 
.A(n_3315),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3464),
.B(n_2376),
.Y(n_3731)
);

HB1xp67_ASAP7_75t_L g3732 ( 
.A(n_3343),
.Y(n_3732)
);

AOI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3344),
.A2(n_1910),
.B1(n_1911),
.B2(n_1908),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3409),
.Y(n_3734)
);

NOR2xp67_ASAP7_75t_L g3735 ( 
.A(n_3455),
.B(n_1913),
.Y(n_3735)
);

O2A1O1Ixp33_ASAP7_75t_L g3736 ( 
.A1(n_3476),
.A2(n_2387),
.B(n_2394),
.C(n_2381),
.Y(n_3736)
);

NAND2xp33_ASAP7_75t_L g3737 ( 
.A(n_3304),
.B(n_1918),
.Y(n_3737)
);

NOR2xp67_ASAP7_75t_L g3738 ( 
.A(n_3415),
.B(n_3400),
.Y(n_3738)
);

NAND3xp33_ASAP7_75t_L g3739 ( 
.A(n_3346),
.B(n_1923),
.C(n_1922),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3382),
.B(n_2396),
.Y(n_3740)
);

AND2x6_ASAP7_75t_SL g3741 ( 
.A(n_3394),
.B(n_3437),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3531),
.B(n_3471),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3436),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3471),
.B(n_2397),
.Y(n_3744)
);

NOR2xp67_ASAP7_75t_L g3745 ( 
.A(n_3513),
.B(n_1925),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3436),
.Y(n_3746)
);

AOI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3331),
.A2(n_1931),
.B1(n_1937),
.B2(n_1929),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3327),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_SL g3749 ( 
.A(n_3545),
.B(n_1938),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3426),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3472),
.B(n_2403),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_3403),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3472),
.B(n_2404),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3417),
.B(n_3482),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3369),
.B(n_2315),
.Y(n_3755)
);

BUFx8_ASAP7_75t_L g3756 ( 
.A(n_3442),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3327),
.Y(n_3757)
);

NOR2xp33_ASAP7_75t_L g3758 ( 
.A(n_3372),
.B(n_1942),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3483),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3482),
.B(n_2413),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3524),
.B(n_2415),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3349),
.B(n_1944),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_L g3763 ( 
.A(n_3373),
.B(n_1948),
.Y(n_3763)
);

A2O1A1Ixp33_ASAP7_75t_L g3764 ( 
.A1(n_3398),
.A2(n_2419),
.B(n_2426),
.C(n_2417),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_SL g3765 ( 
.A(n_3389),
.B(n_1949),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3399),
.B(n_1950),
.Y(n_3766)
);

AOI21x1_ASAP7_75t_L g3767 ( 
.A1(n_3506),
.A2(n_2431),
.B(n_2427),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3324),
.B(n_1955),
.Y(n_3768)
);

OR2x2_ASAP7_75t_L g3769 ( 
.A(n_3486),
.B(n_2592),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3435),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3435),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3489),
.B(n_2441),
.Y(n_3772)
);

AOI22xp33_ASAP7_75t_L g3773 ( 
.A1(n_3378),
.A2(n_2399),
.B1(n_2346),
.B2(n_2603),
.Y(n_3773)
);

OR2x2_ASAP7_75t_L g3774 ( 
.A(n_3461),
.B(n_2614),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3516),
.B(n_2450),
.Y(n_3775)
);

BUFx6f_ASAP7_75t_SL g3776 ( 
.A(n_3519),
.Y(n_3776)
);

BUFx3_ASAP7_75t_L g3777 ( 
.A(n_3532),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_SL g3778 ( 
.A(n_3527),
.B(n_3533),
.Y(n_3778)
);

AOI22xp33_ASAP7_75t_L g3779 ( 
.A1(n_3478),
.A2(n_2399),
.B1(n_2631),
.B2(n_2629),
.Y(n_3779)
);

AOI22xp5_ASAP7_75t_L g3780 ( 
.A1(n_3468),
.A2(n_1958),
.B1(n_1959),
.B2(n_1957),
.Y(n_3780)
);

OR2x2_ASAP7_75t_L g3781 ( 
.A(n_3423),
.B(n_2458),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3517),
.Y(n_3782)
);

AND2x6_ASAP7_75t_L g3783 ( 
.A(n_3490),
.B(n_2469),
.Y(n_3783)
);

NOR2xp33_ASAP7_75t_L g3784 ( 
.A(n_3411),
.B(n_1960),
.Y(n_3784)
);

BUFx3_ASAP7_75t_L g3785 ( 
.A(n_3490),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3467),
.B(n_2475),
.Y(n_3786)
);

NAND3xp33_ASAP7_75t_L g3787 ( 
.A(n_3520),
.B(n_1964),
.C(n_1961),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3493),
.B(n_1966),
.Y(n_3788)
);

HB1xp67_ASAP7_75t_L g3789 ( 
.A(n_3485),
.Y(n_3789)
);

AOI22xp33_ASAP7_75t_SL g3790 ( 
.A1(n_3419),
.A2(n_1969),
.B1(n_1970),
.B2(n_1968),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3492),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3492),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3424),
.A2(n_1973),
.B1(n_1980),
.B2(n_1972),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3424),
.A2(n_1982),
.B1(n_1984),
.B2(n_1981),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3424),
.B(n_2481),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3367),
.B(n_1985),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3424),
.B(n_2482),
.Y(n_3797)
);

NOR2xp33_ASAP7_75t_L g3798 ( 
.A(n_3308),
.B(n_1988),
.Y(n_3798)
);

BUFx3_ASAP7_75t_L g3799 ( 
.A(n_3504),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3308),
.B(n_1991),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3316),
.Y(n_3801)
);

AOI22xp5_ASAP7_75t_L g3802 ( 
.A1(n_3308),
.A2(n_1993),
.B1(n_1994),
.B2(n_1992),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3424),
.B(n_2485),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3424),
.B(n_2489),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3316),
.Y(n_3805)
);

BUFx2_ASAP7_75t_L g3806 ( 
.A(n_3498),
.Y(n_3806)
);

AOI22xp33_ASAP7_75t_L g3807 ( 
.A1(n_3390),
.A2(n_2183),
.B1(n_2219),
.B2(n_2152),
.Y(n_3807)
);

O2A1O1Ixp5_ASAP7_75t_L g3808 ( 
.A1(n_3420),
.A2(n_2279),
.B(n_2291),
.C(n_2223),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3367),
.B(n_1996),
.Y(n_3809)
);

NOR2x1p5_ASAP7_75t_L g3810 ( 
.A(n_3504),
.B(n_1997),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3424),
.B(n_2490),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_3367),
.B(n_1998),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3424),
.B(n_2496),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3316),
.Y(n_3814)
);

O2A1O1Ixp5_ASAP7_75t_L g3815 ( 
.A1(n_3420),
.A2(n_2358),
.B(n_2372),
.C(n_2321),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3424),
.B(n_2508),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3424),
.B(n_2509),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_SL g3818 ( 
.A(n_3333),
.B(n_2003),
.Y(n_3818)
);

NAND3xp33_ASAP7_75t_L g3819 ( 
.A(n_3308),
.B(n_2009),
.C(n_2005),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3316),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3311),
.Y(n_3821)
);

INVx2_ASAP7_75t_SL g3822 ( 
.A(n_3302),
.Y(n_3822)
);

HB1xp67_ASAP7_75t_L g3823 ( 
.A(n_3498),
.Y(n_3823)
);

CKINVDCx5p33_ASAP7_75t_R g3824 ( 
.A(n_3375),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3316),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3424),
.B(n_2524),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3311),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3311),
.Y(n_3828)
);

AOI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3308),
.A2(n_2012),
.B1(n_2014),
.B2(n_2011),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3424),
.B(n_2530),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3424),
.B(n_2531),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3424),
.B(n_2537),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3424),
.B(n_2543),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3367),
.B(n_2015),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3424),
.B(n_2555),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3316),
.Y(n_3836)
);

OR2x2_ASAP7_75t_L g3837 ( 
.A(n_3310),
.B(n_2572),
.Y(n_3837)
);

NOR2xp33_ASAP7_75t_L g3838 ( 
.A(n_3308),
.B(n_2018),
.Y(n_3838)
);

BUFx6f_ASAP7_75t_L g3839 ( 
.A(n_3750),
.Y(n_3839)
);

INVxp67_ASAP7_75t_L g3840 ( 
.A(n_3806),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3570),
.B(n_2024),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3782),
.A2(n_2581),
.B(n_2578),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3559),
.B(n_2025),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3798),
.B(n_2026),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3552),
.Y(n_3845)
);

AOI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3800),
.A2(n_3838),
.B1(n_3571),
.B2(n_3715),
.Y(n_3846)
);

HB1xp67_ASAP7_75t_L g3847 ( 
.A(n_3823),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3633),
.B(n_2028),
.Y(n_3848)
);

A2O1A1Ixp33_ASAP7_75t_L g3849 ( 
.A1(n_3710),
.A2(n_2602),
.B(n_2604),
.C(n_2601),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3554),
.Y(n_3850)
);

BUFx2_ASAP7_75t_L g3851 ( 
.A(n_3667),
.Y(n_3851)
);

OAI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3686),
.A2(n_3661),
.B(n_3555),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3628),
.Y(n_3853)
);

HB1xp67_ASAP7_75t_L g3854 ( 
.A(n_3621),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_SL g3855 ( 
.A(n_3689),
.B(n_2029),
.Y(n_3855)
);

AND2x4_ASAP7_75t_L g3856 ( 
.A(n_3587),
.B(n_2618),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3631),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3662),
.A2(n_2622),
.B(n_2620),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3569),
.B(n_2030),
.Y(n_3859)
);

NAND2xp33_ASAP7_75t_L g3860 ( 
.A(n_3824),
.B(n_2034),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3652),
.Y(n_3861)
);

O2A1O1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3572),
.A2(n_2639),
.B(n_2640),
.C(n_2637),
.Y(n_3862)
);

BUFx6f_ASAP7_75t_L g3863 ( 
.A(n_3588),
.Y(n_3863)
);

NAND2xp33_ASAP7_75t_L g3864 ( 
.A(n_3709),
.B(n_2035),
.Y(n_3864)
);

OAI321xp33_ASAP7_75t_L g3865 ( 
.A1(n_3615),
.A2(n_2663),
.A3(n_2658),
.B1(n_2662),
.B2(n_2644),
.C(n_2474),
.Y(n_3865)
);

AOI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3626),
.A2(n_3682),
.B1(n_3696),
.B2(n_3668),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_L g3867 ( 
.A1(n_3607),
.A2(n_2038),
.B1(n_2040),
.B2(n_2037),
.Y(n_3867)
);

BUFx6f_ASAP7_75t_L g3868 ( 
.A(n_3588),
.Y(n_3868)
);

O2A1O1Ixp33_ASAP7_75t_L g3869 ( 
.A1(n_3577),
.A2(n_2513),
.B(n_2514),
.C(n_2488),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3558),
.B(n_2041),
.Y(n_3870)
);

OAI22xp5_ASAP7_75t_L g3871 ( 
.A1(n_3595),
.A2(n_2050),
.B1(n_2052),
.B2(n_2047),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3560),
.B(n_2055),
.Y(n_3872)
);

INVx3_ASAP7_75t_L g3873 ( 
.A(n_3799),
.Y(n_3873)
);

INVx2_ASAP7_75t_SL g3874 ( 
.A(n_3756),
.Y(n_3874)
);

NOR2xp33_ASAP7_75t_L g3875 ( 
.A(n_3660),
.B(n_2057),
.Y(n_3875)
);

AOI22xp5_ASAP7_75t_L g3876 ( 
.A1(n_3655),
.A2(n_2061),
.B1(n_2062),
.B2(n_2059),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3563),
.B(n_2067),
.Y(n_3877)
);

INVx1_ASAP7_75t_SL g3878 ( 
.A(n_3693),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3565),
.B(n_2070),
.Y(n_3879)
);

BUFx6f_ASAP7_75t_L g3880 ( 
.A(n_3629),
.Y(n_3880)
);

A2O1A1Ixp33_ASAP7_75t_L g3881 ( 
.A1(n_3736),
.A2(n_2073),
.B(n_2074),
.C(n_2072),
.Y(n_3881)
);

OR2x6_ASAP7_75t_L g3882 ( 
.A(n_3573),
.B(n_0),
.Y(n_3882)
);

OAI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3721),
.A2(n_2081),
.B(n_2080),
.Y(n_3883)
);

NOR2xp33_ASAP7_75t_L g3884 ( 
.A(n_3610),
.B(n_2082),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3581),
.B(n_2083),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3718),
.A2(n_2085),
.B(n_2084),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3705),
.B(n_2086),
.Y(n_3887)
);

BUFx6f_ASAP7_75t_L g3888 ( 
.A(n_3629),
.Y(n_3888)
);

AO21x1_ASAP7_75t_L g3889 ( 
.A1(n_3767),
.A2(n_1),
.B(n_2),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3584),
.B(n_2089),
.Y(n_3890)
);

OAI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3585),
.A2(n_2093),
.B1(n_2094),
.B2(n_2091),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3714),
.B(n_3818),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3685),
.B(n_2095),
.Y(n_3893)
);

NOR2xp33_ASAP7_75t_L g3894 ( 
.A(n_3717),
.B(n_2097),
.Y(n_3894)
);

OR2x2_ASAP7_75t_L g3895 ( 
.A(n_3650),
.B(n_3678),
.Y(n_3895)
);

AOI21x1_ASAP7_75t_L g3896 ( 
.A1(n_3699),
.A2(n_191),
.B(n_190),
.Y(n_3896)
);

AOI21xp33_ASAP7_75t_L g3897 ( 
.A1(n_3664),
.A2(n_2103),
.B(n_2102),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3755),
.B(n_2105),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_3647),
.A2(n_2107),
.B(n_2106),
.Y(n_3899)
);

NAND3xp33_ASAP7_75t_L g3900 ( 
.A(n_3567),
.B(n_3829),
.C(n_3802),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3546),
.A2(n_2109),
.B(n_2108),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3796),
.A2(n_2112),
.B(n_2111),
.Y(n_3902)
);

NOR2xp67_ASAP7_75t_L g3903 ( 
.A(n_3556),
.B(n_2116),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3608),
.B(n_2119),
.Y(n_3904)
);

AO21x2_ASAP7_75t_L g3905 ( 
.A1(n_3720),
.A2(n_2125),
.B(n_2120),
.Y(n_3905)
);

OAI22xp5_ASAP7_75t_L g3906 ( 
.A1(n_3801),
.A2(n_3805),
.B1(n_3820),
.B2(n_3814),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3825),
.B(n_2130),
.Y(n_3907)
);

OAI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3684),
.A2(n_2134),
.B(n_2131),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3618),
.Y(n_3909)
);

BUFx6f_ASAP7_75t_L g3910 ( 
.A(n_3659),
.Y(n_3910)
);

AOI21xp5_ASAP7_75t_L g3911 ( 
.A1(n_3809),
.A2(n_3834),
.B(n_3812),
.Y(n_3911)
);

INVxp67_ASAP7_75t_L g3912 ( 
.A(n_3635),
.Y(n_3912)
);

CKINVDCx5p33_ASAP7_75t_R g3913 ( 
.A(n_3701),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3836),
.A2(n_2141),
.B1(n_2142),
.B2(n_2140),
.Y(n_3914)
);

AOI21xp33_ASAP7_75t_L g3915 ( 
.A1(n_3564),
.A2(n_2145),
.B(n_2144),
.Y(n_3915)
);

OAI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_3658),
.A2(n_2150),
.B1(n_2155),
.B2(n_2148),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3694),
.A2(n_2158),
.B(n_2157),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3622),
.B(n_2160),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3673),
.B(n_2162),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3642),
.Y(n_3920)
);

AND2x4_ASAP7_75t_L g3921 ( 
.A(n_3777),
.B(n_2165),
.Y(n_3921)
);

INVx3_ASAP7_75t_L g3922 ( 
.A(n_3573),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3666),
.B(n_2166),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3549),
.A2(n_2168),
.B(n_2167),
.Y(n_3924)
);

OAI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3688),
.A2(n_2172),
.B(n_2169),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3643),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3795),
.A2(n_2174),
.B(n_2173),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3797),
.B(n_2175),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3645),
.Y(n_3929)
);

INVx5_ASAP7_75t_L g3930 ( 
.A(n_3741),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3803),
.A2(n_2181),
.B(n_2180),
.Y(n_3931)
);

NOR2xp33_ASAP7_75t_L g3932 ( 
.A(n_3724),
.B(n_3623),
.Y(n_3932)
);

AOI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_3804),
.A2(n_2185),
.B(n_2184),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3811),
.B(n_3813),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3816),
.B(n_2186),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3817),
.A2(n_2189),
.B(n_2188),
.Y(n_3936)
);

BUFx4f_ASAP7_75t_L g3937 ( 
.A(n_3659),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_SL g3938 ( 
.A(n_3673),
.B(n_2191),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3646),
.Y(n_3939)
);

OAI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3787),
.A2(n_2194),
.B(n_2193),
.Y(n_3940)
);

NAND3xp33_ASAP7_75t_L g3941 ( 
.A(n_3758),
.B(n_2199),
.C(n_2197),
.Y(n_3941)
);

OAI22xp5_ASAP7_75t_L g3942 ( 
.A1(n_3702),
.A2(n_2201),
.B1(n_2202),
.B2(n_2200),
.Y(n_3942)
);

BUFx6f_ASAP7_75t_L g3943 ( 
.A(n_3669),
.Y(n_3943)
);

INVx3_ASAP7_75t_L g3944 ( 
.A(n_3669),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3826),
.B(n_2203),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3830),
.A2(n_3832),
.B(n_3831),
.Y(n_3946)
);

AOI22xp5_ASAP7_75t_L g3947 ( 
.A1(n_3604),
.A2(n_3617),
.B1(n_3657),
.B2(n_3602),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3833),
.B(n_2207),
.Y(n_3948)
);

BUFx6f_ASAP7_75t_L g3949 ( 
.A(n_3596),
.Y(n_3949)
);

AOI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3835),
.A2(n_2212),
.B(n_2210),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3550),
.B(n_2213),
.Y(n_3951)
);

INVx3_ASAP7_75t_L g3952 ( 
.A(n_3653),
.Y(n_3952)
);

OAI21xp33_ASAP7_75t_L g3953 ( 
.A1(n_3599),
.A2(n_2218),
.B(n_2216),
.Y(n_3953)
);

INVx3_ASAP7_75t_L g3954 ( 
.A(n_3713),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3568),
.A2(n_2224),
.B(n_2222),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3649),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3575),
.B(n_2227),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3656),
.Y(n_3958)
);

OAI21xp33_ASAP7_75t_L g3959 ( 
.A1(n_3697),
.A2(n_2231),
.B(n_2228),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3672),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3726),
.B(n_3624),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3634),
.B(n_2233),
.Y(n_3962)
);

OAI321xp33_ASAP7_75t_L g3963 ( 
.A1(n_3675),
.A2(n_2239),
.A3(n_2236),
.B1(n_2242),
.B2(n_2238),
.C(n_2234),
.Y(n_3963)
);

NOR2xp33_ASAP7_75t_L g3964 ( 
.A(n_3742),
.B(n_2244),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3632),
.A2(n_2246),
.B(n_2245),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3674),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3636),
.B(n_3637),
.Y(n_3967)
);

O2A1O1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3706),
.A2(n_2248),
.B(n_2249),
.C(n_2247),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3695),
.A2(n_2251),
.B(n_2250),
.Y(n_3969)
);

A2O1A1Ixp33_ASAP7_75t_L g3970 ( 
.A1(n_3763),
.A2(n_2257),
.B(n_2258),
.C(n_2256),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3703),
.A2(n_2261),
.B(n_2259),
.Y(n_3971)
);

INVxp33_ASAP7_75t_SL g3972 ( 
.A(n_3638),
.Y(n_3972)
);

A2O1A1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_3766),
.A2(n_2264),
.B(n_2265),
.C(n_2262),
.Y(n_3973)
);

AOI21x1_ASAP7_75t_L g3974 ( 
.A1(n_3704),
.A2(n_191),
.B(n_190),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3619),
.B(n_2271),
.Y(n_3975)
);

AND2x4_ASAP7_75t_SL g3976 ( 
.A(n_3732),
.B(n_192),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3683),
.Y(n_3977)
);

AOI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3788),
.A2(n_2274),
.B1(n_2275),
.B2(n_2273),
.Y(n_3978)
);

INVx3_ASAP7_75t_L g3979 ( 
.A(n_3785),
.Y(n_3979)
);

AOI21xp33_ASAP7_75t_L g3980 ( 
.A1(n_3691),
.A2(n_2280),
.B(n_2277),
.Y(n_3980)
);

AND2x2_ASAP7_75t_SL g3981 ( 
.A(n_3594),
.B(n_1),
.Y(n_3981)
);

BUFx3_ASAP7_75t_L g3982 ( 
.A(n_3671),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3707),
.A2(n_3708),
.B(n_3578),
.Y(n_3983)
);

A2O1A1Ixp33_ASAP7_75t_L g3984 ( 
.A1(n_3819),
.A2(n_2288),
.B(n_2289),
.C(n_2286),
.Y(n_3984)
);

O2A1O1Ixp33_ASAP7_75t_L g3985 ( 
.A1(n_3580),
.A2(n_2294),
.B(n_2296),
.C(n_2290),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3681),
.B(n_2298),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3711),
.B(n_2300),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3586),
.A2(n_2303),
.B(n_2302),
.Y(n_3988)
);

BUFx2_ASAP7_75t_L g3989 ( 
.A(n_3665),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3778),
.B(n_2307),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3590),
.A2(n_2310),
.B(n_2309),
.Y(n_3991)
);

BUFx3_ASAP7_75t_L g3992 ( 
.A(n_3613),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3644),
.B(n_2313),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3716),
.B(n_2316),
.Y(n_3994)
);

O2A1O1Ixp5_ASAP7_75t_L g3995 ( 
.A1(n_3611),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_3995)
);

INVx3_ASAP7_75t_L g3996 ( 
.A(n_3776),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3738),
.B(n_2317),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3548),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3551),
.Y(n_3999)
);

BUFx3_ASAP7_75t_L g4000 ( 
.A(n_3791),
.Y(n_4000)
);

CKINVDCx20_ASAP7_75t_R g4001 ( 
.A(n_3752),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_SL g4002 ( 
.A(n_3762),
.B(n_2327),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3562),
.B(n_2328),
.Y(n_4003)
);

NAND2x1p5_ASAP7_75t_L g4004 ( 
.A(n_3822),
.B(n_2),
.Y(n_4004)
);

A2O1A1Ixp33_ASAP7_75t_L g4005 ( 
.A1(n_3712),
.A2(n_2335),
.B(n_2338),
.C(n_2329),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3690),
.Y(n_4006)
);

AOI22xp5_ASAP7_75t_L g4007 ( 
.A1(n_3768),
.A2(n_2340),
.B1(n_2342),
.B2(n_2339),
.Y(n_4007)
);

OAI21xp33_ASAP7_75t_L g4008 ( 
.A1(n_3733),
.A2(n_2347),
.B(n_2343),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3553),
.Y(n_4009)
);

OAI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3761),
.A2(n_2351),
.B(n_2348),
.Y(n_4010)
);

O2A1O1Ixp33_ASAP7_75t_L g4011 ( 
.A1(n_3591),
.A2(n_2354),
.B(n_2355),
.C(n_2352),
.Y(n_4011)
);

AND2x4_ASAP7_75t_L g4012 ( 
.A(n_3730),
.B(n_2357),
.Y(n_4012)
);

INVx1_ASAP7_75t_SL g4013 ( 
.A(n_3774),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_L g4014 ( 
.A(n_3739),
.B(n_2367),
.Y(n_4014)
);

OAI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3625),
.A2(n_2375),
.B(n_2373),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3837),
.B(n_2378),
.Y(n_4016)
);

AOI22xp5_ASAP7_75t_L g4017 ( 
.A1(n_3784),
.A2(n_2383),
.B1(n_2384),
.B2(n_2382),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3759),
.B(n_2385),
.Y(n_4018)
);

AO21x1_ASAP7_75t_L g4019 ( 
.A1(n_3639),
.A2(n_3),
.B(n_4),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3561),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3579),
.Y(n_4021)
);

BUFx6f_ASAP7_75t_L g4022 ( 
.A(n_3748),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3592),
.Y(n_4023)
);

A2O1A1Ixp33_ASAP7_75t_L g4024 ( 
.A1(n_3808),
.A2(n_2388),
.B(n_2389),
.C(n_2386),
.Y(n_4024)
);

OAI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3815),
.A2(n_2393),
.B(n_2392),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3651),
.B(n_2395),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_L g4027 ( 
.A(n_3692),
.B(n_2398),
.Y(n_4027)
);

AND2x4_ASAP7_75t_L g4028 ( 
.A(n_3757),
.B(n_2400),
.Y(n_4028)
);

BUFx12f_ASAP7_75t_L g4029 ( 
.A(n_3783),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3728),
.B(n_2406),
.Y(n_4030)
);

O2A1O1Ixp5_ASAP7_75t_L g4031 ( 
.A1(n_3722),
.A2(n_6),
.B(n_3),
.C(n_5),
.Y(n_4031)
);

NOR2xp33_ASAP7_75t_L g4032 ( 
.A(n_3731),
.B(n_2409),
.Y(n_4032)
);

NOR3xp33_ASAP7_75t_L g4033 ( 
.A(n_3547),
.B(n_3654),
.C(n_3641),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3740),
.B(n_2411),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3679),
.B(n_2412),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3725),
.B(n_2422),
.Y(n_4036)
);

INVx3_ASAP7_75t_L g4037 ( 
.A(n_3792),
.Y(n_4037)
);

BUFx2_ASAP7_75t_L g4038 ( 
.A(n_3700),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3772),
.B(n_2423),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3677),
.B(n_2424),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3663),
.B(n_2425),
.Y(n_4041)
);

OAI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3764),
.A2(n_2433),
.B(n_2430),
.Y(n_4042)
);

BUFx3_ASAP7_75t_L g4043 ( 
.A(n_3789),
.Y(n_4043)
);

OAI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3793),
.A2(n_2435),
.B(n_2434),
.Y(n_4044)
);

A2O1A1Ixp33_ASAP7_75t_L g4045 ( 
.A1(n_3557),
.A2(n_2437),
.B(n_2440),
.C(n_2436),
.Y(n_4045)
);

INVx5_ASAP7_75t_L g4046 ( 
.A(n_3783),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3620),
.B(n_2443),
.Y(n_4047)
);

AOI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_3737),
.A2(n_2445),
.B(n_2444),
.Y(n_4048)
);

OAI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3574),
.A2(n_2447),
.B1(n_2448),
.B2(n_2446),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3598),
.Y(n_4050)
);

AOI22xp5_ASAP7_75t_L g4051 ( 
.A1(n_3698),
.A2(n_3601),
.B1(n_3630),
.B2(n_3676),
.Y(n_4051)
);

BUFx2_ASAP7_75t_SL g4052 ( 
.A(n_3735),
.Y(n_4052)
);

OAI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3794),
.A2(n_2453),
.B(n_2451),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3600),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3749),
.A2(n_2455),
.B(n_2454),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3603),
.B(n_3745),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3605),
.B(n_2463),
.Y(n_4057)
);

AOI21xp5_ASAP7_75t_L g4058 ( 
.A1(n_3765),
.A2(n_2466),
.B(n_2465),
.Y(n_4058)
);

INVx2_ASAP7_75t_SL g4059 ( 
.A(n_3810),
.Y(n_4059)
);

BUFx6f_ASAP7_75t_L g4060 ( 
.A(n_3743),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_3576),
.A2(n_2470),
.B(n_2468),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3606),
.B(n_2472),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_3746),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3612),
.Y(n_4064)
);

OAI21xp33_ASAP7_75t_L g4065 ( 
.A1(n_3747),
.A2(n_2476),
.B(n_2473),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_L g4066 ( 
.A(n_3754),
.B(n_2478),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3614),
.B(n_2483),
.Y(n_4067)
);

BUFx6f_ASAP7_75t_L g4068 ( 
.A(n_3734),
.Y(n_4068)
);

OAI21x1_ASAP7_75t_L g4069 ( 
.A1(n_3771),
.A2(n_6),
.B(n_7),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3616),
.B(n_2486),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3627),
.Y(n_4071)
);

NAND3xp33_ASAP7_75t_L g4072 ( 
.A(n_3744),
.B(n_2492),
.C(n_2491),
.Y(n_4072)
);

INVx2_ASAP7_75t_L g4073 ( 
.A(n_3821),
.Y(n_4073)
);

O2A1O1Ixp33_ASAP7_75t_L g4074 ( 
.A1(n_3751),
.A2(n_2494),
.B(n_2495),
.C(n_2493),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_3566),
.B(n_2497),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3593),
.A2(n_2503),
.B(n_2501),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3828),
.B(n_2504),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_L g4078 ( 
.A(n_3827),
.B(n_2506),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3727),
.Y(n_4079)
);

OAI21xp33_ASAP7_75t_L g4080 ( 
.A1(n_3780),
.A2(n_3760),
.B(n_3753),
.Y(n_4080)
);

AND2x4_ASAP7_75t_L g4081 ( 
.A(n_3719),
.B(n_2507),
.Y(n_4081)
);

BUFx4f_ASAP7_75t_L g4082 ( 
.A(n_3769),
.Y(n_4082)
);

OAI22xp5_ASAP7_75t_SL g4083 ( 
.A1(n_3846),
.A2(n_3790),
.B1(n_3687),
.B2(n_3779),
.Y(n_4083)
);

INVx2_ASAP7_75t_L g4084 ( 
.A(n_3966),
.Y(n_4084)
);

NOR2x1_ASAP7_75t_L g4085 ( 
.A(n_3982),
.B(n_3609),
.Y(n_4085)
);

XOR2xp5_ASAP7_75t_L g4086 ( 
.A(n_3913),
.B(n_3781),
.Y(n_4086)
);

AOI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_3946),
.A2(n_3597),
.B(n_3582),
.Y(n_4087)
);

A2O1A1Ixp33_ASAP7_75t_L g4088 ( 
.A1(n_3900),
.A2(n_3723),
.B(n_3640),
.C(n_3583),
.Y(n_4088)
);

INVx2_ASAP7_75t_SL g4089 ( 
.A(n_3937),
.Y(n_4089)
);

CKINVDCx8_ASAP7_75t_R g4090 ( 
.A(n_3839),
.Y(n_4090)
);

NOR2xp33_ASAP7_75t_L g4091 ( 
.A(n_3947),
.B(n_3932),
.Y(n_4091)
);

BUFx2_ASAP7_75t_L g4092 ( 
.A(n_3851),
.Y(n_4092)
);

AOI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_3934),
.A2(n_3648),
.B(n_3680),
.Y(n_4093)
);

NAND2x1p5_ASAP7_75t_L g4094 ( 
.A(n_3863),
.B(n_3868),
.Y(n_4094)
);

INVx1_ASAP7_75t_SL g4095 ( 
.A(n_3895),
.Y(n_4095)
);

NOR2xp33_ASAP7_75t_L g4096 ( 
.A(n_3972),
.B(n_3775),
.Y(n_4096)
);

BUFx6f_ASAP7_75t_SL g4097 ( 
.A(n_3874),
.Y(n_4097)
);

BUFx6f_ASAP7_75t_L g4098 ( 
.A(n_3839),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_4016),
.B(n_3807),
.Y(n_4099)
);

CKINVDCx5p33_ASAP7_75t_R g4100 ( 
.A(n_4001),
.Y(n_4100)
);

AO32x1_ASAP7_75t_L g4101 ( 
.A1(n_3906),
.A2(n_3770),
.A3(n_3773),
.B1(n_3729),
.B2(n_3786),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3977),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_SL g4103 ( 
.A(n_4046),
.B(n_3589),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3845),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_3840),
.B(n_3670),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3873),
.Y(n_4106)
);

AOI22xp5_ASAP7_75t_L g4107 ( 
.A1(n_4030),
.A2(n_2512),
.B1(n_2515),
.B2(n_2511),
.Y(n_4107)
);

BUFx2_ASAP7_75t_L g4108 ( 
.A(n_3847),
.Y(n_4108)
);

BUFx6f_ASAP7_75t_L g4109 ( 
.A(n_3863),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3961),
.B(n_3967),
.Y(n_4110)
);

OAI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3844),
.A2(n_2522),
.B1(n_2526),
.B2(n_2520),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3850),
.Y(n_4112)
);

NAND2x1p5_ASAP7_75t_L g4113 ( 
.A(n_3868),
.B(n_7),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3909),
.Y(n_4114)
);

OA22x2_ASAP7_75t_L g4115 ( 
.A1(n_3882),
.A2(n_2529),
.B1(n_2532),
.B2(n_2527),
.Y(n_4115)
);

AOI22xp33_ASAP7_75t_SL g4116 ( 
.A1(n_3957),
.A2(n_2536),
.B1(n_2538),
.B2(n_2534),
.Y(n_4116)
);

BUFx6f_ASAP7_75t_L g4117 ( 
.A(n_3880),
.Y(n_4117)
);

A2O1A1Ixp33_ASAP7_75t_L g4118 ( 
.A1(n_4080),
.A2(n_2540),
.B(n_2541),
.C(n_2539),
.Y(n_4118)
);

OAI21x1_ASAP7_75t_L g4119 ( 
.A1(n_4069),
.A2(n_195),
.B(n_194),
.Y(n_4119)
);

AOI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_3983),
.A2(n_2544),
.B(n_2542),
.Y(n_4120)
);

BUFx2_ASAP7_75t_L g4121 ( 
.A(n_3979),
.Y(n_4121)
);

AOI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_3911),
.A2(n_3893),
.B(n_4002),
.Y(n_4122)
);

INVx3_ASAP7_75t_SL g4123 ( 
.A(n_3882),
.Y(n_4123)
);

NOR3xp33_ASAP7_75t_SL g4124 ( 
.A(n_3941),
.B(n_2549),
.C(n_2545),
.Y(n_4124)
);

NOR2xp33_ASAP7_75t_R g4125 ( 
.A(n_3855),
.B(n_2552),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_4032),
.B(n_2553),
.Y(n_4126)
);

AOI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_3981),
.A2(n_2559),
.B1(n_2560),
.B2(n_2554),
.Y(n_4127)
);

INVx3_ASAP7_75t_L g4128 ( 
.A(n_3880),
.Y(n_4128)
);

OAI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_3859),
.A2(n_3876),
.B1(n_3978),
.B2(n_3848),
.Y(n_4129)
);

AOI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_3892),
.A2(n_2564),
.B1(n_2565),
.B2(n_2561),
.Y(n_4130)
);

NOR2xp33_ASAP7_75t_L g4131 ( 
.A(n_3854),
.B(n_2566),
.Y(n_4131)
);

OAI21xp33_ASAP7_75t_L g4132 ( 
.A1(n_3897),
.A2(n_2570),
.B(n_2568),
.Y(n_4132)
);

HB1xp67_ASAP7_75t_L g4133 ( 
.A(n_3878),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3960),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_4038),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3887),
.B(n_2571),
.Y(n_4136)
);

AOI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_3928),
.A2(n_2576),
.B(n_2575),
.Y(n_4137)
);

INVx5_ASAP7_75t_L g4138 ( 
.A(n_4029),
.Y(n_4138)
);

CKINVDCx8_ASAP7_75t_R g4139 ( 
.A(n_4046),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3875),
.B(n_2577),
.Y(n_4140)
);

BUFx10_ASAP7_75t_L g4141 ( 
.A(n_3888),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_3898),
.B(n_2579),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3926),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3920),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4036),
.B(n_2582),
.Y(n_4145)
);

A2O1A1Ixp33_ASAP7_75t_L g4146 ( 
.A1(n_3862),
.A2(n_3849),
.B(n_3959),
.C(n_3963),
.Y(n_4146)
);

BUFx5_ASAP7_75t_L g4147 ( 
.A(n_3929),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3956),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_3989),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_3912),
.B(n_2584),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3987),
.B(n_2585),
.Y(n_4151)
);

INVx3_ASAP7_75t_SL g4152 ( 
.A(n_3888),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4006),
.Y(n_4153)
);

A2O1A1Ixp33_ASAP7_75t_L g4154 ( 
.A1(n_3968),
.A2(n_4014),
.B(n_3980),
.C(n_3881),
.Y(n_4154)
);

AOI22xp33_ASAP7_75t_L g4155 ( 
.A1(n_4028),
.A2(n_2587),
.B1(n_2590),
.B2(n_2586),
.Y(n_4155)
);

BUFx2_ASAP7_75t_L g4156 ( 
.A(n_3992),
.Y(n_4156)
);

AOI21xp5_ASAP7_75t_L g4157 ( 
.A1(n_3935),
.A2(n_3948),
.B(n_3945),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3964),
.B(n_2594),
.Y(n_4158)
);

NOR2xp33_ASAP7_75t_L g4159 ( 
.A(n_4051),
.B(n_2595),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3884),
.B(n_2596),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3870),
.B(n_3872),
.Y(n_4161)
);

BUFx3_ASAP7_75t_L g4162 ( 
.A(n_3910),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3877),
.B(n_2598),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3939),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3879),
.B(n_2599),
.Y(n_4165)
);

INVx1_ASAP7_75t_SL g4166 ( 
.A(n_4013),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3958),
.Y(n_4167)
);

AOI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_3860),
.A2(n_2607),
.B1(n_2608),
.B2(n_2605),
.Y(n_4168)
);

AOI221xp5_ASAP7_75t_L g4169 ( 
.A1(n_3915),
.A2(n_2612),
.B1(n_2613),
.B2(n_2611),
.C(n_2609),
.Y(n_4169)
);

AND2x4_ASAP7_75t_L g4170 ( 
.A(n_3922),
.B(n_2615),
.Y(n_4170)
);

NOR2xp33_ASAP7_75t_L g4171 ( 
.A(n_3894),
.B(n_2616),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_3951),
.A2(n_2619),
.B(n_2617),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_L g4173 ( 
.A(n_3864),
.B(n_2621),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4082),
.B(n_2623),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3841),
.B(n_2626),
.Y(n_4175)
);

OR2x6_ASAP7_75t_SL g4176 ( 
.A(n_3942),
.B(n_2627),
.Y(n_4176)
);

O2A1O1Ixp33_ASAP7_75t_SL g4177 ( 
.A1(n_3970),
.A2(n_197),
.B(n_198),
.C(n_196),
.Y(n_4177)
);

BUFx6f_ASAP7_75t_L g4178 ( 
.A(n_3910),
.Y(n_4178)
);

OAI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_4027),
.A2(n_2630),
.B1(n_2632),
.B2(n_2628),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3994),
.B(n_3986),
.Y(n_4180)
);

CKINVDCx10_ASAP7_75t_R g4181 ( 
.A(n_3930),
.Y(n_4181)
);

O2A1O1Ixp5_ASAP7_75t_L g4182 ( 
.A1(n_4075),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_4182)
);

NAND3xp33_ASAP7_75t_SL g4183 ( 
.A(n_4044),
.B(n_4053),
.C(n_4017),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4021),
.Y(n_4184)
);

AOI33xp33_ASAP7_75t_L g4185 ( 
.A1(n_3867),
.A2(n_2652),
.A3(n_2636),
.B1(n_2653),
.B2(n_2646),
.B3(n_2635),
.Y(n_4185)
);

A2O1A1Ixp33_ASAP7_75t_L g4186 ( 
.A1(n_3865),
.A2(n_2661),
.B(n_10),
.C(n_8),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_3856),
.B(n_199),
.Y(n_4187)
);

BUFx6f_ASAP7_75t_L g4188 ( 
.A(n_3943),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3918),
.B(n_11),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_3930),
.B(n_201),
.Y(n_4190)
);

OAI22xp5_ASAP7_75t_L g4191 ( 
.A1(n_3973),
.A2(n_202),
.B1(n_204),
.B2(n_201),
.Y(n_4191)
);

AOI21xp5_ASAP7_75t_L g4192 ( 
.A1(n_4024),
.A2(n_204),
.B(n_202),
.Y(n_4192)
);

INVxp67_ASAP7_75t_SL g4193 ( 
.A(n_4000),
.Y(n_4193)
);

CKINVDCx5p33_ASAP7_75t_R g4194 ( 
.A(n_3943),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_3949),
.B(n_205),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_4034),
.B(n_11),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4054),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3975),
.B(n_12),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_3962),
.B(n_12),
.Y(n_4199)
);

INVx1_ASAP7_75t_SL g4200 ( 
.A(n_3949),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_3858),
.A2(n_206),
.B(n_205),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_4026),
.B(n_206),
.Y(n_4202)
);

NOR2xp33_ASAP7_75t_L g4203 ( 
.A(n_4041),
.B(n_207),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_3853),
.Y(n_4204)
);

NOR2xp33_ASAP7_75t_L g4205 ( 
.A(n_3953),
.B(n_207),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_4040),
.B(n_13),
.Y(n_4206)
);

OAI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_4010),
.A2(n_209),
.B1(n_210),
.B2(n_208),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_3857),
.Y(n_4208)
);

INVx4_ASAP7_75t_L g4209 ( 
.A(n_3996),
.Y(n_4209)
);

BUFx4f_ASAP7_75t_L g4210 ( 
.A(n_3952),
.Y(n_4210)
);

BUFx12f_ASAP7_75t_L g4211 ( 
.A(n_3921),
.Y(n_4211)
);

O2A1O1Ixp33_ASAP7_75t_L g4212 ( 
.A1(n_4005),
.A2(n_4045),
.B(n_3984),
.C(n_4011),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_4068),
.B(n_208),
.Y(n_4213)
);

OAI22xp5_ASAP7_75t_SL g4214 ( 
.A1(n_4004),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4071),
.Y(n_4215)
);

OAI22xp5_ASAP7_75t_L g4216 ( 
.A1(n_3885),
.A2(n_210),
.B1(n_211),
.B2(n_209),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4039),
.B(n_13),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_4043),
.Y(n_4218)
);

BUFx12f_ASAP7_75t_L g4219 ( 
.A(n_4059),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_3990),
.B(n_14),
.Y(n_4220)
);

OAI22xp5_ASAP7_75t_L g4221 ( 
.A1(n_3890),
.A2(n_212),
.B1(n_213),
.B2(n_211),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3954),
.B(n_16),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_4008),
.B(n_212),
.Y(n_4223)
);

AOI21xp5_ASAP7_75t_L g4224 ( 
.A1(n_3908),
.A2(n_214),
.B(n_213),
.Y(n_4224)
);

AOI21xp5_ASAP7_75t_L g4225 ( 
.A1(n_3925),
.A2(n_215),
.B(n_214),
.Y(n_4225)
);

BUFx6f_ASAP7_75t_L g4226 ( 
.A(n_4022),
.Y(n_4226)
);

BUFx8_ASAP7_75t_L g4227 ( 
.A(n_4012),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_3869),
.A2(n_3917),
.B(n_3842),
.Y(n_4228)
);

A2O1A1Ixp33_ASAP7_75t_L g4229 ( 
.A1(n_3985),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_4068),
.B(n_215),
.Y(n_4230)
);

OAI22xp5_ASAP7_75t_L g4231 ( 
.A1(n_3904),
.A2(n_217),
.B1(n_218),
.B2(n_216),
.Y(n_4231)
);

NAND3xp33_ASAP7_75t_SL g4232 ( 
.A(n_4007),
.B(n_17),
.C(n_18),
.Y(n_4232)
);

O2A1O1Ixp33_ASAP7_75t_L g4233 ( 
.A1(n_3883),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_4233)
);

OAI22xp5_ASAP7_75t_L g4234 ( 
.A1(n_3907),
.A2(n_3923),
.B1(n_3871),
.B2(n_4072),
.Y(n_4234)
);

NOR2xp33_ASAP7_75t_R g4235 ( 
.A(n_3944),
.B(n_216),
.Y(n_4235)
);

OAI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4047),
.A2(n_218),
.B1(n_219),
.B2(n_217),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3861),
.Y(n_4237)
);

AND2x4_ASAP7_75t_L g4238 ( 
.A(n_4056),
.B(n_20),
.Y(n_4238)
);

INVx4_ASAP7_75t_L g4239 ( 
.A(n_4022),
.Y(n_4239)
);

OAI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_3899),
.A2(n_20),
.B(n_21),
.Y(n_4240)
);

AND2x4_ASAP7_75t_L g4241 ( 
.A(n_4037),
.B(n_20),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_3998),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_3976),
.B(n_219),
.Y(n_4243)
);

O2A1O1Ixp5_ASAP7_75t_L g4244 ( 
.A1(n_3940),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_4244)
);

O2A1O1Ixp5_ASAP7_75t_L g4245 ( 
.A1(n_3995),
.A2(n_24),
.B(n_21),
.C(n_23),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4081),
.B(n_23),
.Y(n_4246)
);

INVxp67_ASAP7_75t_L g4247 ( 
.A(n_4079),
.Y(n_4247)
);

BUFx2_ASAP7_75t_L g4248 ( 
.A(n_3997),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_3999),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4009),
.Y(n_4250)
);

NOR2x1_ASAP7_75t_L g4251 ( 
.A(n_4052),
.B(n_3903),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4020),
.Y(n_4252)
);

AND2x4_ASAP7_75t_L g4253 ( 
.A(n_4060),
.B(n_24),
.Y(n_4253)
);

INVx1_ASAP7_75t_SL g4254 ( 
.A(n_4063),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4023),
.Y(n_4255)
);

A2O1A1Ixp33_ASAP7_75t_L g4256 ( 
.A1(n_4074),
.A2(n_4031),
.B(n_4065),
.C(n_3927),
.Y(n_4256)
);

O2A1O1Ixp33_ASAP7_75t_L g4257 ( 
.A1(n_4049),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_4257)
);

NAND3xp33_ASAP7_75t_SL g4258 ( 
.A(n_4033),
.B(n_25),
.C(n_26),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4050),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4064),
.Y(n_4260)
);

AO32x2_ASAP7_75t_L g4261 ( 
.A1(n_3891),
.A2(n_27),
.A3(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_4261)
);

AOI22xp33_ASAP7_75t_L g4262 ( 
.A1(n_4042),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_4262)
);

AOI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_3924),
.A2(n_221),
.B(n_220),
.Y(n_4263)
);

NOR2xp33_ASAP7_75t_L g4264 ( 
.A(n_4066),
.B(n_221),
.Y(n_4264)
);

BUFx6f_ASAP7_75t_L g4265 ( 
.A(n_4073),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_3931),
.A2(n_223),
.B(n_222),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_3914),
.B(n_224),
.Y(n_4267)
);

HB1xp67_ASAP7_75t_L g4268 ( 
.A(n_4018),
.Y(n_4268)
);

INVxp33_ASAP7_75t_SL g4269 ( 
.A(n_3916),
.Y(n_4269)
);

AOI21x1_ASAP7_75t_L g4270 ( 
.A1(n_3974),
.A2(n_30),
.B(n_31),
.Y(n_4270)
);

NOR2xp67_ASAP7_75t_L g4271 ( 
.A(n_3886),
.B(n_30),
.Y(n_4271)
);

AOI22xp5_ASAP7_75t_L g4272 ( 
.A1(n_3993),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_3933),
.B(n_32),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4035),
.B(n_225),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_L g4275 ( 
.A(n_4003),
.B(n_226),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4057),
.Y(n_4276)
);

NOR2xp33_ASAP7_75t_R g4277 ( 
.A(n_3896),
.B(n_226),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_4019),
.B(n_227),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4062),
.Y(n_4279)
);

AOI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_3936),
.A2(n_228),
.B(n_227),
.Y(n_4280)
);

BUFx2_ASAP7_75t_L g4281 ( 
.A(n_3905),
.Y(n_4281)
);

BUFx6f_ASAP7_75t_L g4282 ( 
.A(n_3919),
.Y(n_4282)
);

NOR2xp33_ASAP7_75t_L g4283 ( 
.A(n_3938),
.B(n_228),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4067),
.B(n_34),
.Y(n_4284)
);

AOI221xp5_ASAP7_75t_L g4285 ( 
.A1(n_3965),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_4285)
);

A2O1A1Ixp33_ASAP7_75t_L g4286 ( 
.A1(n_3950),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_4286)
);

CKINVDCx5p33_ASAP7_75t_R g4287 ( 
.A(n_4076),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_3955),
.A2(n_3889),
.B(n_3969),
.Y(n_4288)
);

AOI33xp33_ASAP7_75t_L g4289 ( 
.A1(n_4048),
.A2(n_41),
.A3(n_43),
.B1(n_39),
.B2(n_40),
.B3(n_42),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_4078),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4070),
.Y(n_4291)
);

CKINVDCx16_ASAP7_75t_R g4292 ( 
.A(n_4015),
.Y(n_4292)
);

OR2x6_ASAP7_75t_L g4293 ( 
.A(n_3988),
.B(n_41),
.Y(n_4293)
);

INVx3_ASAP7_75t_L g4294 ( 
.A(n_4077),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_R g4295 ( 
.A(n_3991),
.B(n_229),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_4025),
.Y(n_4296)
);

CKINVDCx5p33_ASAP7_75t_R g4297 ( 
.A(n_4055),
.Y(n_4297)
);

A2O1A1Ixp33_ASAP7_75t_SL g4298 ( 
.A1(n_3971),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_4298)
);

O2A1O1Ixp5_ASAP7_75t_SL g4299 ( 
.A1(n_3901),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_3902),
.Y(n_4300)
);

A2O1A1Ixp33_ASAP7_75t_L g4301 ( 
.A1(n_4058),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4061),
.A2(n_233),
.B(n_231),
.Y(n_4302)
);

OA22x2_ASAP7_75t_L g4303 ( 
.A1(n_3866),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_4303)
);

BUFx2_ASAP7_75t_L g4304 ( 
.A(n_3851),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_SL g4305 ( 
.A(n_3846),
.B(n_233),
.Y(n_4305)
);

A2O1A1Ixp33_ASAP7_75t_L g4306 ( 
.A1(n_3846),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_4306)
);

INVx3_ASAP7_75t_L g4307 ( 
.A(n_3863),
.Y(n_4307)
);

NOR2xp33_ASAP7_75t_L g4308 ( 
.A(n_3846),
.B(n_234),
.Y(n_4308)
);

CKINVDCx8_ASAP7_75t_R g4309 ( 
.A(n_3913),
.Y(n_4309)
);

AOI22xp5_ASAP7_75t_L g4310 ( 
.A1(n_3846),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_3846),
.B(n_50),
.Y(n_4311)
);

INVx8_ASAP7_75t_L g4312 ( 
.A(n_4029),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3966),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_4016),
.B(n_235),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3966),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4016),
.B(n_236),
.Y(n_4316)
);

BUFx12f_ASAP7_75t_L g4317 ( 
.A(n_3913),
.Y(n_4317)
);

BUFx2_ASAP7_75t_L g4318 ( 
.A(n_3851),
.Y(n_4318)
);

INVx4_ASAP7_75t_L g4319 ( 
.A(n_3863),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_3846),
.B(n_52),
.Y(n_4320)
);

INVx4_ASAP7_75t_L g4321 ( 
.A(n_3863),
.Y(n_4321)
);

OR2x6_ASAP7_75t_L g4322 ( 
.A(n_3839),
.B(n_52),
.Y(n_4322)
);

BUFx2_ASAP7_75t_L g4323 ( 
.A(n_3851),
.Y(n_4323)
);

O2A1O1Ixp33_ASAP7_75t_L g4324 ( 
.A1(n_3843),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_4324)
);

OAI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_3846),
.A2(n_237),
.B1(n_238),
.B2(n_236),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_3846),
.B(n_53),
.Y(n_4326)
);

HB1xp67_ASAP7_75t_L g4327 ( 
.A(n_3847),
.Y(n_4327)
);

BUFx2_ASAP7_75t_L g4328 ( 
.A(n_3851),
.Y(n_4328)
);

CKINVDCx16_ASAP7_75t_R g4329 ( 
.A(n_4001),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_SL g4330 ( 
.A(n_3846),
.B(n_237),
.Y(n_4330)
);

O2A1O1Ixp5_ASAP7_75t_L g4331 ( 
.A1(n_3852),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_3846),
.A2(n_239),
.B1(n_240),
.B2(n_238),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4313),
.Y(n_4333)
);

AOI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4091),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_4334)
);

AOI21xp33_ASAP7_75t_L g4335 ( 
.A1(n_4159),
.A2(n_57),
.B(n_58),
.Y(n_4335)
);

AOI21xp5_ASAP7_75t_L g4336 ( 
.A1(n_4183),
.A2(n_240),
.B(n_239),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4110),
.B(n_58),
.Y(n_4337)
);

BUFx6f_ASAP7_75t_L g4338 ( 
.A(n_4090),
.Y(n_4338)
);

AO32x2_ASAP7_75t_L g4339 ( 
.A1(n_4083),
.A2(n_61),
.A3(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_4339)
);

O2A1O1Ixp33_ASAP7_75t_L g4340 ( 
.A1(n_4308),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4314),
.B(n_242),
.Y(n_4341)
);

AO22x2_ASAP7_75t_L g4342 ( 
.A1(n_4129),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_SL g4343 ( 
.A(n_4292),
.B(n_243),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4157),
.A2(n_244),
.B(n_243),
.Y(n_4344)
);

AND2x4_ASAP7_75t_L g4345 ( 
.A(n_4089),
.B(n_245),
.Y(n_4345)
);

NOR2xp33_ASAP7_75t_L g4346 ( 
.A(n_4269),
.B(n_248),
.Y(n_4346)
);

OAI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_4171),
.A2(n_4126),
.B(n_4146),
.Y(n_4347)
);

CKINVDCx16_ASAP7_75t_R g4348 ( 
.A(n_4329),
.Y(n_4348)
);

OAI21x1_ASAP7_75t_SL g4349 ( 
.A1(n_4311),
.A2(n_64),
.B(n_65),
.Y(n_4349)
);

AOI21xp5_ASAP7_75t_SL g4350 ( 
.A1(n_4088),
.A2(n_66),
.B(n_67),
.Y(n_4350)
);

AO31x2_ASAP7_75t_L g4351 ( 
.A1(n_4281),
.A2(n_69),
.A3(n_67),
.B(n_68),
.Y(n_4351)
);

NOR2xp33_ASAP7_75t_L g4352 ( 
.A(n_4096),
.B(n_249),
.Y(n_4352)
);

AO32x2_ASAP7_75t_L g4353 ( 
.A1(n_4325),
.A2(n_69),
.A3(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_4353)
);

CKINVDCx5p33_ASAP7_75t_R g4354 ( 
.A(n_4100),
.Y(n_4354)
);

INVx3_ASAP7_75t_L g4355 ( 
.A(n_4139),
.Y(n_4355)
);

A2O1A1Ixp33_ASAP7_75t_L g4356 ( 
.A1(n_4264),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4095),
.B(n_72),
.Y(n_4357)
);

OAI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_4158),
.A2(n_4326),
.B(n_4320),
.Y(n_4358)
);

AOI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_4087),
.A2(n_251),
.B(n_250),
.Y(n_4359)
);

OA21x2_ASAP7_75t_L g4360 ( 
.A1(n_4331),
.A2(n_72),
.B(n_73),
.Y(n_4360)
);

AOI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_4122),
.A2(n_253),
.B(n_252),
.Y(n_4361)
);

AOI21xp5_ASAP7_75t_L g4362 ( 
.A1(n_4288),
.A2(n_255),
.B(n_254),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4084),
.Y(n_4363)
);

OAI21x1_ASAP7_75t_L g4364 ( 
.A1(n_4119),
.A2(n_256),
.B(n_255),
.Y(n_4364)
);

O2A1O1Ixp33_ASAP7_75t_SL g4365 ( 
.A1(n_4305),
.A2(n_257),
.B(n_258),
.C(n_256),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4133),
.B(n_73),
.Y(n_4366)
);

AOI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_4228),
.A2(n_260),
.B(n_257),
.Y(n_4367)
);

AOI21xp5_ASAP7_75t_L g4368 ( 
.A1(n_4161),
.A2(n_261),
.B(n_260),
.Y(n_4368)
);

OAI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_4151),
.A2(n_74),
.B(n_75),
.Y(n_4369)
);

AOI21x1_ASAP7_75t_SL g4370 ( 
.A1(n_4273),
.A2(n_75),
.B(n_76),
.Y(n_4370)
);

NAND3xp33_ASAP7_75t_L g4371 ( 
.A(n_4205),
.B(n_75),
.C(n_76),
.Y(n_4371)
);

OAI22x1_ASAP7_75t_L g4372 ( 
.A1(n_4123),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_4372)
);

OAI21x1_ASAP7_75t_L g4373 ( 
.A1(n_4270),
.A2(n_262),
.B(n_261),
.Y(n_4373)
);

AOI211x1_ASAP7_75t_L g4374 ( 
.A1(n_4220),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4315),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4102),
.Y(n_4376)
);

NAND2x1p5_ASAP7_75t_L g4377 ( 
.A(n_4210),
.B(n_263),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4108),
.B(n_78),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4327),
.B(n_79),
.Y(n_4379)
);

AOI21x1_ASAP7_75t_L g4380 ( 
.A1(n_4296),
.A2(n_79),
.B(n_80),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4268),
.B(n_80),
.Y(n_4381)
);

NAND2xp33_ASAP7_75t_R g4382 ( 
.A(n_4125),
.B(n_81),
.Y(n_4382)
);

BUFx6f_ASAP7_75t_SL g4383 ( 
.A(n_4098),
.Y(n_4383)
);

O2A1O1Ixp5_ASAP7_75t_SL g4384 ( 
.A1(n_4278),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_4384)
);

OAI21x1_ASAP7_75t_L g4385 ( 
.A1(n_4300),
.A2(n_265),
.B(n_264),
.Y(n_4385)
);

OAI21x1_ASAP7_75t_L g4386 ( 
.A1(n_4299),
.A2(n_4192),
.B(n_4148),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4180),
.B(n_81),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4290),
.B(n_82),
.Y(n_4388)
);

OAI21xp5_ASAP7_75t_L g4389 ( 
.A1(n_4160),
.A2(n_82),
.B(n_83),
.Y(n_4389)
);

NAND3xp33_ASAP7_75t_L g4390 ( 
.A(n_4223),
.B(n_83),
.C(n_84),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4104),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4276),
.B(n_85),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4291),
.B(n_85),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_SL g4394 ( 
.A1(n_4154),
.A2(n_85),
.B(n_86),
.Y(n_4394)
);

BUFx2_ASAP7_75t_L g4395 ( 
.A(n_4092),
.Y(n_4395)
);

O2A1O1Ixp5_ASAP7_75t_L g4396 ( 
.A1(n_4330),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_4396)
);

AO32x2_ASAP7_75t_L g4397 ( 
.A1(n_4332),
.A2(n_89),
.A3(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_4397)
);

INVx2_ASAP7_75t_SL g4398 ( 
.A(n_4098),
.Y(n_4398)
);

BUFx6f_ASAP7_75t_L g4399 ( 
.A(n_4152),
.Y(n_4399)
);

INVx5_ASAP7_75t_L g4400 ( 
.A(n_4312),
.Y(n_4400)
);

OAI21x1_ASAP7_75t_L g4401 ( 
.A1(n_4143),
.A2(n_266),
.B(n_264),
.Y(n_4401)
);

OAI21x1_ASAP7_75t_L g4402 ( 
.A1(n_4153),
.A2(n_267),
.B(n_266),
.Y(n_4402)
);

NOR2xp33_ASAP7_75t_L g4403 ( 
.A(n_4176),
.B(n_267),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4112),
.Y(n_4404)
);

BUFx12f_ASAP7_75t_L g4405 ( 
.A(n_4194),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4135),
.B(n_88),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_4279),
.B(n_89),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4294),
.B(n_89),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4316),
.B(n_269),
.Y(n_4409)
);

AO31x2_ASAP7_75t_L g4410 ( 
.A1(n_4256),
.A2(n_92),
.A3(n_90),
.B(n_91),
.Y(n_4410)
);

NAND3xp33_ASAP7_75t_SL g4411 ( 
.A(n_4295),
.B(n_90),
.C(n_92),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4140),
.A2(n_92),
.B(n_93),
.Y(n_4412)
);

AO31x2_ASAP7_75t_L g4413 ( 
.A1(n_4186),
.A2(n_95),
.A3(n_93),
.B(n_94),
.Y(n_4413)
);

OAI21x1_ASAP7_75t_L g4414 ( 
.A1(n_4134),
.A2(n_273),
.B(n_272),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4184),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_4166),
.B(n_93),
.Y(n_4416)
);

OA21x2_ASAP7_75t_L g4417 ( 
.A1(n_4244),
.A2(n_94),
.B(n_95),
.Y(n_4417)
);

BUFx12f_ASAP7_75t_L g4418 ( 
.A(n_4317),
.Y(n_4418)
);

OAI21x1_ASAP7_75t_L g4419 ( 
.A1(n_4245),
.A2(n_277),
.B(n_275),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4197),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4099),
.B(n_94),
.Y(n_4421)
);

AOI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_4234),
.A2(n_278),
.B(n_277),
.Y(n_4422)
);

AND2x4_ASAP7_75t_L g4423 ( 
.A(n_4162),
.B(n_4138),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_4141),
.Y(n_4424)
);

AO32x2_ASAP7_75t_L g4425 ( 
.A1(n_4207),
.A2(n_97),
.A3(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_4425)
);

INVxp67_ASAP7_75t_SL g4426 ( 
.A(n_4147),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4304),
.B(n_96),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_4318),
.B(n_96),
.Y(n_4428)
);

NOR4xp25_ASAP7_75t_L g4429 ( 
.A(n_4258),
.B(n_4306),
.C(n_4232),
.D(n_4324),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4093),
.A2(n_280),
.B(n_279),
.Y(n_4430)
);

OA21x2_ASAP7_75t_L g4431 ( 
.A1(n_4240),
.A2(n_97),
.B(n_98),
.Y(n_4431)
);

AOI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_4224),
.A2(n_280),
.B(n_279),
.Y(n_4432)
);

OAI21xp5_ASAP7_75t_L g4433 ( 
.A1(n_4173),
.A2(n_99),
.B(n_100),
.Y(n_4433)
);

NOR2xp33_ASAP7_75t_L g4434 ( 
.A(n_4086),
.B(n_281),
.Y(n_4434)
);

AOI22x1_ASAP7_75t_L g4435 ( 
.A1(n_4225),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_4435)
);

AOI21xp5_ASAP7_75t_L g4436 ( 
.A1(n_4233),
.A2(n_4212),
.B(n_4101),
.Y(n_4436)
);

NOR2x1_ASAP7_75t_L g4437 ( 
.A(n_4251),
.B(n_100),
.Y(n_4437)
);

NOR2xp67_ASAP7_75t_L g4438 ( 
.A(n_4209),
.B(n_101),
.Y(n_4438)
);

BUFx6f_ASAP7_75t_L g4439 ( 
.A(n_4109),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4114),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4187),
.B(n_281),
.Y(n_4441)
);

NOR2xp33_ASAP7_75t_L g4442 ( 
.A(n_4149),
.B(n_282),
.Y(n_4442)
);

AOI21xp5_ASAP7_75t_L g4443 ( 
.A1(n_4101),
.A2(n_283),
.B(n_282),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4215),
.Y(n_4444)
);

NOR2xp33_ASAP7_75t_SL g4445 ( 
.A(n_4309),
.B(n_102),
.Y(n_4445)
);

OAI21x1_ASAP7_75t_L g4446 ( 
.A1(n_4302),
.A2(n_285),
.B(n_284),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4144),
.Y(n_4447)
);

BUFx6f_ASAP7_75t_L g4448 ( 
.A(n_4109),
.Y(n_4448)
);

AOI21x1_ASAP7_75t_L g4449 ( 
.A1(n_4120),
.A2(n_102),
.B(n_103),
.Y(n_4449)
);

NAND2x1p5_ASAP7_75t_L g4450 ( 
.A(n_4138),
.B(n_286),
.Y(n_4450)
);

AOI21x1_ASAP7_75t_L g4451 ( 
.A1(n_4103),
.A2(n_102),
.B(n_103),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4164),
.Y(n_4452)
);

BUFx3_ASAP7_75t_L g4453 ( 
.A(n_4218),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_SL g4454 ( 
.A(n_4147),
.B(n_289),
.Y(n_4454)
);

OAI21x1_ASAP7_75t_L g4455 ( 
.A1(n_4263),
.A2(n_292),
.B(n_291),
.Y(n_4455)
);

NAND3xp33_ASAP7_75t_L g4456 ( 
.A(n_4202),
.B(n_4203),
.C(n_4310),
.Y(n_4456)
);

BUFx2_ASAP7_75t_L g4457 ( 
.A(n_4323),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_SL g4458 ( 
.A(n_4147),
.B(n_291),
.Y(n_4458)
);

AOI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_4177),
.A2(n_293),
.B(n_292),
.Y(n_4459)
);

BUFx6f_ASAP7_75t_SL g4460 ( 
.A(n_4322),
.Y(n_4460)
);

OAI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4266),
.A2(n_295),
.B(n_294),
.Y(n_4461)
);

OAI21xp5_ASAP7_75t_L g4462 ( 
.A1(n_4118),
.A2(n_103),
.B(n_104),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4167),
.Y(n_4463)
);

OAI21x1_ASAP7_75t_L g4464 ( 
.A1(n_4280),
.A2(n_297),
.B(n_296),
.Y(n_4464)
);

AOI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_4201),
.A2(n_298),
.B(n_296),
.Y(n_4465)
);

AOI21x1_ASAP7_75t_L g4466 ( 
.A1(n_4271),
.A2(n_4199),
.B(n_4217),
.Y(n_4466)
);

OAI21x1_ASAP7_75t_L g4467 ( 
.A1(n_4182),
.A2(n_299),
.B(n_298),
.Y(n_4467)
);

BUFx2_ASAP7_75t_L g4468 ( 
.A(n_4328),
.Y(n_4468)
);

BUFx3_ASAP7_75t_L g4469 ( 
.A(n_4094),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4193),
.B(n_104),
.Y(n_4470)
);

OAI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_4107),
.A2(n_105),
.B(n_106),
.Y(n_4471)
);

AO21x2_ASAP7_75t_L g4472 ( 
.A1(n_4277),
.A2(n_105),
.B(n_106),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4105),
.B(n_4156),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4252),
.Y(n_4474)
);

NOR2xp67_ASAP7_75t_SL g4475 ( 
.A(n_4211),
.B(n_107),
.Y(n_4475)
);

AOI221x1_ASAP7_75t_L g4476 ( 
.A1(n_4191),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.C(n_110),
.Y(n_4476)
);

AO21x1_ASAP7_75t_L g4477 ( 
.A1(n_4257),
.A2(n_107),
.B(n_108),
.Y(n_4477)
);

AOI21xp5_ASAP7_75t_SL g4478 ( 
.A1(n_4229),
.A2(n_108),
.B(n_109),
.Y(n_4478)
);

AO31x2_ASAP7_75t_L g4479 ( 
.A1(n_4204),
.A2(n_111),
.A3(n_109),
.B(n_110),
.Y(n_4479)
);

OAI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4111),
.A2(n_110),
.B(n_111),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4255),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_SL g4482 ( 
.A(n_4147),
.B(n_4282),
.Y(n_4482)
);

BUFx6f_ASAP7_75t_L g4483 ( 
.A(n_4117),
.Y(n_4483)
);

AND2x4_ASAP7_75t_L g4484 ( 
.A(n_4319),
.B(n_300),
.Y(n_4484)
);

OA22x2_ASAP7_75t_L g4485 ( 
.A1(n_4322),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_4485)
);

AOI21xp5_ASAP7_75t_L g4486 ( 
.A1(n_4298),
.A2(n_302),
.B(n_301),
.Y(n_4486)
);

AOI21xp5_ASAP7_75t_L g4487 ( 
.A1(n_4189),
.A2(n_305),
.B(n_303),
.Y(n_4487)
);

CKINVDCx6p67_ASAP7_75t_R g4488 ( 
.A(n_4181),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_4198),
.A2(n_305),
.B(n_303),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4121),
.B(n_112),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_4208),
.Y(n_4491)
);

OAI21x1_ASAP7_75t_L g4492 ( 
.A1(n_4259),
.A2(n_307),
.B(n_306),
.Y(n_4492)
);

AOI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_4196),
.A2(n_310),
.B(n_309),
.Y(n_4493)
);

NAND2x1p5_ASAP7_75t_L g4494 ( 
.A(n_4321),
.B(n_4117),
.Y(n_4494)
);

AOI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_4206),
.A2(n_310),
.B(n_309),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4262),
.A2(n_4165),
.B(n_4163),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_4237),
.Y(n_4497)
);

AOI21xp33_ASAP7_75t_L g4498 ( 
.A1(n_4132),
.A2(n_113),
.B(n_114),
.Y(n_4498)
);

NAND3xp33_ASAP7_75t_L g4499 ( 
.A(n_4285),
.B(n_114),
.C(n_115),
.Y(n_4499)
);

INVxp67_ASAP7_75t_L g4500 ( 
.A(n_4106),
.Y(n_4500)
);

AO21x2_ASAP7_75t_L g4501 ( 
.A1(n_4137),
.A2(n_115),
.B(n_116),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4241),
.B(n_115),
.Y(n_4502)
);

AOI21xp5_ASAP7_75t_SL g4503 ( 
.A1(n_4286),
.A2(n_116),
.B(n_117),
.Y(n_4503)
);

OAI21x1_ASAP7_75t_L g4504 ( 
.A1(n_4242),
.A2(n_313),
.B(n_312),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4254),
.B(n_116),
.Y(n_4505)
);

AOI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_4297),
.A2(n_316),
.B(n_315),
.Y(n_4506)
);

AO31x2_ASAP7_75t_L g4507 ( 
.A1(n_4249),
.A2(n_4260),
.A3(n_4250),
.B(n_4301),
.Y(n_4507)
);

AOI21x1_ASAP7_75t_L g4508 ( 
.A1(n_4213),
.A2(n_117),
.B(n_118),
.Y(n_4508)
);

OAI21x1_ASAP7_75t_L g4509 ( 
.A1(n_4230),
.A2(n_316),
.B(n_315),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_4307),
.B(n_4239),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4274),
.B(n_117),
.Y(n_4511)
);

BUFx6f_ASAP7_75t_L g4512 ( 
.A(n_4178),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4267),
.B(n_317),
.Y(n_4513)
);

AOI22xp5_ASAP7_75t_L g4514 ( 
.A1(n_4303),
.A2(n_4275),
.B1(n_4214),
.B2(n_4283),
.Y(n_4514)
);

AOI21xp5_ASAP7_75t_L g4515 ( 
.A1(n_4293),
.A2(n_320),
.B(n_318),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4247),
.Y(n_4516)
);

AOI22xp5_ASAP7_75t_L g4517 ( 
.A1(n_4238),
.A2(n_4142),
.B1(n_4145),
.B2(n_4115),
.Y(n_4517)
);

NAND3x1_ASAP7_75t_L g4518 ( 
.A(n_4085),
.B(n_118),
.C(n_119),
.Y(n_4518)
);

NAND3xp33_ASAP7_75t_SL g4519 ( 
.A(n_4235),
.B(n_118),
.C(n_119),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4289),
.B(n_119),
.Y(n_4520)
);

AOI21xp5_ASAP7_75t_L g4521 ( 
.A1(n_4293),
.A2(n_322),
.B(n_321),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4200),
.B(n_120),
.Y(n_4522)
);

INVx3_ASAP7_75t_L g4523 ( 
.A(n_4188),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4265),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4265),
.Y(n_4525)
);

NAND2x1p5_ASAP7_75t_L g4526 ( 
.A(n_4188),
.B(n_323),
.Y(n_4526)
);

OAI22x1_ASAP7_75t_L g4527 ( 
.A1(n_4113),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_4527)
);

AOI221x1_ASAP7_75t_L g4528 ( 
.A1(n_4236),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_4528)
);

AOI22xp5_ASAP7_75t_L g4529 ( 
.A1(n_4116),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_4529)
);

AOI22xp33_ASAP7_75t_L g4530 ( 
.A1(n_4347),
.A2(n_4284),
.B1(n_4246),
.B2(n_4248),
.Y(n_4530)
);

INVxp67_ASAP7_75t_L g4531 ( 
.A(n_4473),
.Y(n_4531)
);

OAI21x1_ASAP7_75t_SL g4532 ( 
.A1(n_4471),
.A2(n_4221),
.B(n_4216),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4391),
.Y(n_4533)
);

CKINVDCx20_ASAP7_75t_R g4534 ( 
.A(n_4488),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4404),
.Y(n_4535)
);

INVxp67_ASAP7_75t_SL g4536 ( 
.A(n_4426),
.Y(n_4536)
);

AO31x2_ASAP7_75t_L g4537 ( 
.A1(n_4436),
.A2(n_4231),
.A3(n_4179),
.B(n_4172),
.Y(n_4537)
);

NOR2xp33_ASAP7_75t_L g4538 ( 
.A(n_4346),
.B(n_4128),
.Y(n_4538)
);

INVx3_ASAP7_75t_SL g4539 ( 
.A(n_4354),
.Y(n_4539)
);

O2A1O1Ixp33_ASAP7_75t_SL g4540 ( 
.A1(n_4356),
.A2(n_4195),
.B(n_4190),
.C(n_4222),
.Y(n_4540)
);

INVxp67_ASAP7_75t_L g4541 ( 
.A(n_4395),
.Y(n_4541)
);

AND2x4_ASAP7_75t_L g4542 ( 
.A(n_4457),
.B(n_4226),
.Y(n_4542)
);

INVx3_ASAP7_75t_L g4543 ( 
.A(n_4338),
.Y(n_4543)
);

OAI21x1_ASAP7_75t_L g4544 ( 
.A1(n_4367),
.A2(n_4386),
.B(n_4362),
.Y(n_4544)
);

OAI22xp33_ASAP7_75t_SL g4545 ( 
.A1(n_4514),
.A2(n_4127),
.B1(n_4272),
.B2(n_4287),
.Y(n_4545)
);

INVxp67_ASAP7_75t_L g4546 ( 
.A(n_4468),
.Y(n_4546)
);

OAI21x1_ASAP7_75t_L g4547 ( 
.A1(n_4385),
.A2(n_4175),
.B(n_4150),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4415),
.Y(n_4548)
);

AOI21x1_ASAP7_75t_L g4549 ( 
.A1(n_4466),
.A2(n_4136),
.B(n_4253),
.Y(n_4549)
);

BUFx4f_ASAP7_75t_SL g4550 ( 
.A(n_4418),
.Y(n_4550)
);

INVxp33_ASAP7_75t_SL g4551 ( 
.A(n_4453),
.Y(n_4551)
);

BUFx3_ASAP7_75t_L g4552 ( 
.A(n_4399),
.Y(n_4552)
);

NAND3xp33_ASAP7_75t_L g4553 ( 
.A(n_4456),
.B(n_4124),
.C(n_4185),
.Y(n_4553)
);

INVx4_ASAP7_75t_L g4554 ( 
.A(n_4400),
.Y(n_4554)
);

INVx1_ASAP7_75t_SL g4555 ( 
.A(n_4338),
.Y(n_4555)
);

BUFx3_ASAP7_75t_L g4556 ( 
.A(n_4399),
.Y(n_4556)
);

INVx4_ASAP7_75t_L g4557 ( 
.A(n_4405),
.Y(n_4557)
);

BUFx12f_ASAP7_75t_L g4558 ( 
.A(n_4439),
.Y(n_4558)
);

AND2x4_ASAP7_75t_L g4559 ( 
.A(n_4500),
.B(n_4226),
.Y(n_4559)
);

OA21x2_ASAP7_75t_L g4560 ( 
.A1(n_4443),
.A2(n_4131),
.B(n_4155),
.Y(n_4560)
);

OA21x2_ASAP7_75t_L g4561 ( 
.A1(n_4336),
.A2(n_4130),
.B(n_4169),
.Y(n_4561)
);

NAND2x1p5_ASAP7_75t_L g4562 ( 
.A(n_4355),
.B(n_4439),
.Y(n_4562)
);

OAI21x1_ASAP7_75t_L g4563 ( 
.A1(n_4359),
.A2(n_4243),
.B(n_4261),
.Y(n_4563)
);

OAI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_4422),
.A2(n_4168),
.B(n_4170),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4420),
.Y(n_4565)
);

INVx1_ASAP7_75t_SL g4566 ( 
.A(n_4448),
.Y(n_4566)
);

AO31x2_ASAP7_75t_L g4567 ( 
.A1(n_4476),
.A2(n_4261),
.A3(n_4227),
.B(n_125),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_L g4568 ( 
.A1(n_4361),
.A2(n_4174),
.B(n_4312),
.Y(n_4568)
);

OA21x2_ASAP7_75t_L g4569 ( 
.A1(n_4373),
.A2(n_4097),
.B(n_123),
.Y(n_4569)
);

CKINVDCx8_ASAP7_75t_R g4570 ( 
.A(n_4348),
.Y(n_4570)
);

AOI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4382),
.A2(n_4352),
.B1(n_4343),
.B2(n_4411),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_SL g4572 ( 
.A(n_4358),
.B(n_4219),
.Y(n_4572)
);

BUFx3_ASAP7_75t_L g4573 ( 
.A(n_4423),
.Y(n_4573)
);

BUFx5_ASAP7_75t_L g4574 ( 
.A(n_4524),
.Y(n_4574)
);

OAI21x1_ASAP7_75t_L g4575 ( 
.A1(n_4364),
.A2(n_124),
.B(n_126),
.Y(n_4575)
);

INVx2_ASAP7_75t_SL g4576 ( 
.A(n_4483),
.Y(n_4576)
);

OAI21x1_ASAP7_75t_L g4577 ( 
.A1(n_4446),
.A2(n_124),
.B(n_126),
.Y(n_4577)
);

OAI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_4394),
.A2(n_127),
.B(n_128),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4444),
.Y(n_4579)
);

AO31x2_ASAP7_75t_L g4580 ( 
.A1(n_4477),
.A2(n_4481),
.A3(n_4474),
.B(n_4375),
.Y(n_4580)
);

BUFx3_ASAP7_75t_L g4581 ( 
.A(n_4448),
.Y(n_4581)
);

AOI21xp5_ASAP7_75t_L g4582 ( 
.A1(n_4350),
.A2(n_325),
.B(n_324),
.Y(n_4582)
);

OAI21x1_ASAP7_75t_L g4583 ( 
.A1(n_4380),
.A2(n_127),
.B(n_128),
.Y(n_4583)
);

O2A1O1Ixp33_ASAP7_75t_L g4584 ( 
.A1(n_4335),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4333),
.Y(n_4585)
);

NAND2x1p5_ASAP7_75t_L g4586 ( 
.A(n_4512),
.B(n_4469),
.Y(n_4586)
);

OAI21x1_ASAP7_75t_L g4587 ( 
.A1(n_4455),
.A2(n_129),
.B(n_130),
.Y(n_4587)
);

OAI21x1_ASAP7_75t_L g4588 ( 
.A1(n_4461),
.A2(n_129),
.B(n_131),
.Y(n_4588)
);

NOR2xp33_ASAP7_75t_L g4589 ( 
.A(n_4442),
.B(n_324),
.Y(n_4589)
);

OAI21x1_ASAP7_75t_L g4590 ( 
.A1(n_4464),
.A2(n_131),
.B(n_132),
.Y(n_4590)
);

NAND2x1p5_ASAP7_75t_L g4591 ( 
.A(n_4512),
.B(n_325),
.Y(n_4591)
);

CKINVDCx5p33_ASAP7_75t_R g4592 ( 
.A(n_4383),
.Y(n_4592)
);

A2O1A1Ixp33_ASAP7_75t_L g4593 ( 
.A1(n_4496),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4363),
.Y(n_4594)
);

HB1xp67_ASAP7_75t_L g4595 ( 
.A(n_4410),
.Y(n_4595)
);

BUFx2_ASAP7_75t_L g4596 ( 
.A(n_4510),
.Y(n_4596)
);

OAI22xp33_ASAP7_75t_L g4597 ( 
.A1(n_4485),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_4597)
);

HB1xp67_ASAP7_75t_L g4598 ( 
.A(n_4482),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_4376),
.Y(n_4599)
);

OAI21x1_ASAP7_75t_SL g4600 ( 
.A1(n_4433),
.A2(n_327),
.B(n_326),
.Y(n_4600)
);

OAI211xp5_ASAP7_75t_L g4601 ( 
.A1(n_4340),
.A2(n_136),
.B(n_133),
.C(n_135),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4440),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4447),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4421),
.B(n_326),
.Y(n_4604)
);

OAI21x1_ASAP7_75t_L g4605 ( 
.A1(n_4419),
.A2(n_135),
.B(n_136),
.Y(n_4605)
);

OAI21xp5_ASAP7_75t_L g4606 ( 
.A1(n_4432),
.A2(n_136),
.B(n_137),
.Y(n_4606)
);

AO21x2_ASAP7_75t_L g4607 ( 
.A1(n_4459),
.A2(n_137),
.B(n_138),
.Y(n_4607)
);

CKINVDCx6p67_ASAP7_75t_R g4608 ( 
.A(n_4460),
.Y(n_4608)
);

AO21x2_ASAP7_75t_L g4609 ( 
.A1(n_4462),
.A2(n_137),
.B(n_138),
.Y(n_4609)
);

OA21x2_ASAP7_75t_L g4610 ( 
.A1(n_4492),
.A2(n_138),
.B(n_139),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4463),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4337),
.B(n_139),
.Y(n_4612)
);

OAI21x1_ASAP7_75t_L g4613 ( 
.A1(n_4344),
.A2(n_140),
.B(n_141),
.Y(n_4613)
);

INVx3_ASAP7_75t_L g4614 ( 
.A(n_4494),
.Y(n_4614)
);

OR2x6_ASAP7_75t_L g4615 ( 
.A(n_4515),
.B(n_140),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4452),
.Y(n_4616)
);

AOI21x1_ASAP7_75t_L g4617 ( 
.A1(n_4454),
.A2(n_142),
.B(n_143),
.Y(n_4617)
);

OAI21x1_ASAP7_75t_L g4618 ( 
.A1(n_4504),
.A2(n_4370),
.B(n_4401),
.Y(n_4618)
);

AOI22xp33_ASAP7_75t_SL g4619 ( 
.A1(n_4342),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_4619)
);

AND2x4_ASAP7_75t_L g4620 ( 
.A(n_4525),
.B(n_327),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4491),
.Y(n_4621)
);

AOI22xp33_ASAP7_75t_L g4622 ( 
.A1(n_4499),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_4622)
);

OAI21x1_ASAP7_75t_L g4623 ( 
.A1(n_4402),
.A2(n_144),
.B(n_145),
.Y(n_4623)
);

BUFx6f_ASAP7_75t_L g4624 ( 
.A(n_4398),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4516),
.Y(n_4625)
);

O2A1O1Ixp33_ASAP7_75t_L g4626 ( 
.A1(n_4519),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_4523),
.Y(n_4627)
);

BUFx2_ASAP7_75t_L g4628 ( 
.A(n_4424),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4497),
.Y(n_4629)
);

NOR2xp33_ASAP7_75t_SL g4630 ( 
.A(n_4475),
.B(n_147),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4507),
.Y(n_4631)
);

O2A1O1Ixp33_ASAP7_75t_L g4632 ( 
.A1(n_4369),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4513),
.B(n_151),
.Y(n_4633)
);

AOI21x1_ASAP7_75t_L g4634 ( 
.A1(n_4458),
.A2(n_152),
.B(n_153),
.Y(n_4634)
);

A2O1A1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4412),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_4635)
);

AOI21xp5_ASAP7_75t_L g4636 ( 
.A1(n_4430),
.A2(n_331),
.B(n_330),
.Y(n_4636)
);

AOI22xp33_ASAP7_75t_L g4637 ( 
.A1(n_4371),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_4637)
);

AOI21xp5_ASAP7_75t_L g4638 ( 
.A1(n_4465),
.A2(n_331),
.B(n_330),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4479),
.Y(n_4639)
);

INVx3_ASAP7_75t_L g4640 ( 
.A(n_4484),
.Y(n_4640)
);

NAND2x1p5_ASAP7_75t_L g4641 ( 
.A(n_4437),
.B(n_332),
.Y(n_4641)
);

OAI22xp5_ASAP7_75t_L g4642 ( 
.A1(n_4334),
.A2(n_333),
.B1(n_334),
.B2(n_332),
.Y(n_4642)
);

INVx1_ASAP7_75t_SL g4643 ( 
.A(n_4388),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4387),
.B(n_155),
.Y(n_4644)
);

AO21x2_ASAP7_75t_L g4645 ( 
.A1(n_4449),
.A2(n_156),
.B(n_158),
.Y(n_4645)
);

NOR2xp67_ASAP7_75t_L g4646 ( 
.A(n_4390),
.B(n_158),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4381),
.B(n_158),
.Y(n_4647)
);

OAI21x1_ASAP7_75t_L g4648 ( 
.A1(n_4414),
.A2(n_159),
.B(n_160),
.Y(n_4648)
);

OAI22xp5_ASAP7_75t_SL g4649 ( 
.A1(n_4403),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4479),
.Y(n_4650)
);

OR2x6_ASAP7_75t_L g4651 ( 
.A(n_4521),
.B(n_160),
.Y(n_4651)
);

INVx1_ASAP7_75t_SL g4652 ( 
.A(n_4441),
.Y(n_4652)
);

AOI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4478),
.A2(n_335),
.B(n_334),
.Y(n_4653)
);

AOI22xp33_ASAP7_75t_L g4654 ( 
.A1(n_4480),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_4654)
);

AOI22xp33_ASAP7_75t_L g4655 ( 
.A1(n_4389),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_4655)
);

AND2x4_ASAP7_75t_L g4656 ( 
.A(n_4507),
.B(n_336),
.Y(n_4656)
);

INVx4_ASAP7_75t_L g4657 ( 
.A(n_4377),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4351),
.Y(n_4658)
);

AOI22xp5_ASAP7_75t_L g4659 ( 
.A1(n_4445),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_SL g4660 ( 
.A(n_4429),
.B(n_337),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4341),
.B(n_338),
.Y(n_4661)
);

BUFx12f_ASAP7_75t_L g4662 ( 
.A(n_4345),
.Y(n_4662)
);

AO32x2_ASAP7_75t_L g4663 ( 
.A1(n_4339),
.A2(n_167),
.A3(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4531),
.B(n_4379),
.Y(n_4664)
);

BUFx2_ASAP7_75t_L g4665 ( 
.A(n_4541),
.Y(n_4665)
);

NOR2xp33_ASAP7_75t_L g4666 ( 
.A(n_4551),
.B(n_4434),
.Y(n_4666)
);

AOI221xp5_ASAP7_75t_L g4667 ( 
.A1(n_4597),
.A2(n_4372),
.B1(n_4487),
.B2(n_4493),
.C(n_4489),
.Y(n_4667)
);

HB1xp67_ASAP7_75t_L g4668 ( 
.A(n_4546),
.Y(n_4668)
);

INVx8_ASAP7_75t_L g4669 ( 
.A(n_4558),
.Y(n_4669)
);

AOI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4536),
.A2(n_4503),
.B(n_4365),
.Y(n_4670)
);

BUFx3_ASAP7_75t_L g4671 ( 
.A(n_4552),
.Y(n_4671)
);

BUFx2_ASAP7_75t_R g4672 ( 
.A(n_4570),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4625),
.B(n_4392),
.Y(n_4673)
);

AOI21xp5_ASAP7_75t_L g4674 ( 
.A1(n_4532),
.A2(n_4506),
.B(n_4431),
.Y(n_4674)
);

NAND2xp5_ASAP7_75t_L g4675 ( 
.A(n_4533),
.B(n_4393),
.Y(n_4675)
);

AND2x4_ASAP7_75t_L g4676 ( 
.A(n_4573),
.B(n_4438),
.Y(n_4676)
);

OR2x2_ASAP7_75t_L g4677 ( 
.A(n_4535),
.B(n_4378),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4652),
.B(n_4542),
.Y(n_4678)
);

AOI21x1_ASAP7_75t_L g4679 ( 
.A1(n_4549),
.A2(n_4451),
.B(n_4508),
.Y(n_4679)
);

AOI21x1_ASAP7_75t_L g4680 ( 
.A1(n_4572),
.A2(n_4470),
.B(n_4368),
.Y(n_4680)
);

BUFx10_ASAP7_75t_L g4681 ( 
.A(n_4592),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4596),
.B(n_4409),
.Y(n_4682)
);

OAI21x1_ASAP7_75t_L g4683 ( 
.A1(n_4544),
.A2(n_4435),
.B(n_4467),
.Y(n_4683)
);

AND2x4_ASAP7_75t_L g4684 ( 
.A(n_4556),
.B(n_4472),
.Y(n_4684)
);

OA21x2_ASAP7_75t_L g4685 ( 
.A1(n_4658),
.A2(n_4528),
.B(n_4495),
.Y(n_4685)
);

BUFx2_ASAP7_75t_R g4686 ( 
.A(n_4627),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4548),
.B(n_4407),
.Y(n_4687)
);

OAI21x1_ASAP7_75t_L g4688 ( 
.A1(n_4618),
.A2(n_4384),
.B(n_4486),
.Y(n_4688)
);

AO21x2_ASAP7_75t_L g4689 ( 
.A1(n_4639),
.A2(n_4349),
.B(n_4520),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4565),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_SL g4691 ( 
.A(n_4643),
.B(n_4517),
.Y(n_4691)
);

OA21x2_ASAP7_75t_L g4692 ( 
.A1(n_4650),
.A2(n_4366),
.B(n_4406),
.Y(n_4692)
);

AND2x4_ASAP7_75t_L g4693 ( 
.A(n_4598),
.B(n_4490),
.Y(n_4693)
);

AOI21xp5_ASAP7_75t_L g4694 ( 
.A1(n_4593),
.A2(n_4498),
.B(n_4396),
.Y(n_4694)
);

NAND2x1p5_ASAP7_75t_L g4695 ( 
.A(n_4554),
.B(n_4509),
.Y(n_4695)
);

BUFx12f_ASAP7_75t_L g4696 ( 
.A(n_4557),
.Y(n_4696)
);

OAI21x1_ASAP7_75t_L g4697 ( 
.A1(n_4631),
.A2(n_4360),
.B(n_4417),
.Y(n_4697)
);

NOR2xp33_ASAP7_75t_R g4698 ( 
.A(n_4534),
.B(n_4550),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_4539),
.Y(n_4699)
);

INVx8_ASAP7_75t_L g4700 ( 
.A(n_4662),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4579),
.Y(n_4701)
);

CKINVDCx5p33_ASAP7_75t_R g4702 ( 
.A(n_4608),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4559),
.B(n_4427),
.Y(n_4703)
);

BUFx3_ASAP7_75t_L g4704 ( 
.A(n_4628),
.Y(n_4704)
);

BUFx3_ASAP7_75t_L g4705 ( 
.A(n_4543),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_SL g4706 ( 
.A(n_4574),
.B(n_4374),
.Y(n_4706)
);

OR2x2_ASAP7_75t_L g4707 ( 
.A(n_4585),
.B(n_4603),
.Y(n_4707)
);

A2O1A1Ixp33_ASAP7_75t_L g4708 ( 
.A1(n_4632),
.A2(n_4529),
.B(n_4511),
.C(n_4408),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4616),
.Y(n_4709)
);

AO31x2_ASAP7_75t_L g4710 ( 
.A1(n_4635),
.A2(n_4527),
.A3(n_4357),
.B(n_4339),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4629),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4574),
.B(n_4428),
.Y(n_4712)
);

AO21x2_ASAP7_75t_L g4713 ( 
.A1(n_4595),
.A2(n_4416),
.B(n_4505),
.Y(n_4713)
);

OA21x2_ASAP7_75t_L g4714 ( 
.A1(n_4656),
.A2(n_4522),
.B(n_4502),
.Y(n_4714)
);

BUFx12f_ASAP7_75t_L g4715 ( 
.A(n_4624),
.Y(n_4715)
);

OAI21x1_ASAP7_75t_L g4716 ( 
.A1(n_4547),
.A2(n_4518),
.B(n_4526),
.Y(n_4716)
);

INVx2_ASAP7_75t_SL g4717 ( 
.A(n_4624),
.Y(n_4717)
);

INVx1_ASAP7_75t_SL g4718 ( 
.A(n_4555),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4594),
.Y(n_4719)
);

INVxp67_ASAP7_75t_SL g4720 ( 
.A(n_4599),
.Y(n_4720)
);

INVx2_ASAP7_75t_SL g4721 ( 
.A(n_4581),
.Y(n_4721)
);

INVx6_ASAP7_75t_L g4722 ( 
.A(n_4657),
.Y(n_4722)
);

OAI21x1_ASAP7_75t_L g4723 ( 
.A1(n_4623),
.A2(n_4450),
.B(n_4425),
.Y(n_4723)
);

NAND2x1p5_ASAP7_75t_L g4724 ( 
.A(n_4566),
.B(n_4353),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4580),
.B(n_4612),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4602),
.Y(n_4726)
);

AOI21xp5_ASAP7_75t_L g4727 ( 
.A1(n_4578),
.A2(n_4501),
.B(n_4425),
.Y(n_4727)
);

OR2x2_ASAP7_75t_L g4728 ( 
.A(n_4604),
.B(n_4413),
.Y(n_4728)
);

AOI21xp5_ASAP7_75t_L g4729 ( 
.A1(n_4582),
.A2(n_4397),
.B(n_4353),
.Y(n_4729)
);

INVx3_ASAP7_75t_L g4730 ( 
.A(n_4586),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4580),
.B(n_165),
.Y(n_4731)
);

AO31x2_ASAP7_75t_L g4732 ( 
.A1(n_4611),
.A2(n_4397),
.A3(n_168),
.B(n_166),
.Y(n_4732)
);

NAND2x1p5_ASAP7_75t_L g4733 ( 
.A(n_4614),
.B(n_340),
.Y(n_4733)
);

CKINVDCx20_ASAP7_75t_R g4734 ( 
.A(n_4576),
.Y(n_4734)
);

NOR2x1_ASAP7_75t_SL g4735 ( 
.A(n_4615),
.B(n_341),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4538),
.B(n_168),
.Y(n_4736)
);

OAI22xp5_ASAP7_75t_L g4737 ( 
.A1(n_4571),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_4737)
);

INVx4_ASAP7_75t_L g4738 ( 
.A(n_4640),
.Y(n_4738)
);

NOR2xp33_ASAP7_75t_L g4739 ( 
.A(n_4589),
.B(n_342),
.Y(n_4739)
);

OAI21xp5_ASAP7_75t_L g4740 ( 
.A1(n_4653),
.A2(n_4638),
.B(n_4636),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4621),
.Y(n_4741)
);

OR2x2_ASAP7_75t_L g4742 ( 
.A(n_4644),
.B(n_170),
.Y(n_4742)
);

BUFx8_ASAP7_75t_L g4743 ( 
.A(n_4661),
.Y(n_4743)
);

AOI22xp5_ASAP7_75t_L g4744 ( 
.A1(n_4630),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4583),
.Y(n_4745)
);

AO31x2_ASAP7_75t_L g4746 ( 
.A1(n_4642),
.A2(n_173),
.A3(n_171),
.B(n_172),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4663),
.Y(n_4747)
);

NOR2xp33_ASAP7_75t_L g4748 ( 
.A(n_4562),
.B(n_342),
.Y(n_4748)
);

NAND2x1p5_ASAP7_75t_L g4749 ( 
.A(n_4568),
.B(n_343),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4569),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4663),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4647),
.B(n_174),
.Y(n_4752)
);

OA21x2_ASAP7_75t_L g4753 ( 
.A1(n_4563),
.A2(n_174),
.B(n_175),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4645),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4537),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4633),
.B(n_176),
.Y(n_4756)
);

OAI21xp33_ASAP7_75t_L g4757 ( 
.A1(n_4660),
.A2(n_176),
.B(n_177),
.Y(n_4757)
);

AOI22xp5_ASAP7_75t_L g4758 ( 
.A1(n_4649),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_4758)
);

HB1xp67_ASAP7_75t_L g4759 ( 
.A(n_4537),
.Y(n_4759)
);

AO21x2_ASAP7_75t_L g4760 ( 
.A1(n_4646),
.A2(n_178),
.B(n_179),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4610),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4567),
.B(n_179),
.Y(n_4762)
);

BUFx12f_ASAP7_75t_L g4763 ( 
.A(n_4620),
.Y(n_4763)
);

NOR2x1_ASAP7_75t_SL g4764 ( 
.A(n_4615),
.B(n_344),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4567),
.B(n_180),
.Y(n_4765)
);

OAI21xp5_ASAP7_75t_L g4766 ( 
.A1(n_4601),
.A2(n_180),
.B(n_181),
.Y(n_4766)
);

AO22x2_ASAP7_75t_L g4767 ( 
.A1(n_4553),
.A2(n_183),
.B1(n_180),
.B2(n_182),
.Y(n_4767)
);

AOI21x1_ASAP7_75t_L g4768 ( 
.A1(n_4617),
.A2(n_182),
.B(n_183),
.Y(n_4768)
);

AO21x2_ASAP7_75t_L g4769 ( 
.A1(n_4600),
.A2(n_183),
.B(n_184),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4648),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4605),
.Y(n_4771)
);

BUFx2_ASAP7_75t_L g4772 ( 
.A(n_4651),
.Y(n_4772)
);

OR2x2_ASAP7_75t_L g4773 ( 
.A(n_4530),
.B(n_186),
.Y(n_4773)
);

INVx2_ASAP7_75t_SL g4774 ( 
.A(n_4591),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4619),
.B(n_186),
.Y(n_4775)
);

OAI21x1_ASAP7_75t_L g4776 ( 
.A1(n_4634),
.A2(n_186),
.B(n_187),
.Y(n_4776)
);

AOI22xp33_ASAP7_75t_L g4777 ( 
.A1(n_4545),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_4777)
);

OA21x2_ASAP7_75t_L g4778 ( 
.A1(n_4575),
.A2(n_187),
.B(n_188),
.Y(n_4778)
);

BUFx2_ASAP7_75t_L g4779 ( 
.A(n_4641),
.Y(n_4779)
);

AND2x4_ASAP7_75t_L g4780 ( 
.A(n_4564),
.B(n_345),
.Y(n_4780)
);

A2O1A1Ixp33_ASAP7_75t_L g4781 ( 
.A1(n_4626),
.A2(n_188),
.B(n_189),
.C(n_345),
.Y(n_4781)
);

NOR2x1_ASAP7_75t_L g4782 ( 
.A(n_4607),
.B(n_189),
.Y(n_4782)
);

HB1xp67_ASAP7_75t_L g4783 ( 
.A(n_4609),
.Y(n_4783)
);

AO21x2_ASAP7_75t_L g4784 ( 
.A1(n_4606),
.A2(n_4587),
.B(n_4577),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4659),
.B(n_346),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4588),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4560),
.B(n_348),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4707),
.Y(n_4788)
);

HB1xp67_ASAP7_75t_L g4789 ( 
.A(n_4668),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_4709),
.Y(n_4790)
);

INVx2_ASAP7_75t_L g4791 ( 
.A(n_4719),
.Y(n_4791)
);

INVx2_ASAP7_75t_SL g4792 ( 
.A(n_4671),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4690),
.Y(n_4793)
);

INVx3_ASAP7_75t_L g4794 ( 
.A(n_4715),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4665),
.B(n_4590),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4701),
.Y(n_4796)
);

HB1xp67_ASAP7_75t_L g4797 ( 
.A(n_4725),
.Y(n_4797)
);

INVxp67_ASAP7_75t_SL g4798 ( 
.A(n_4692),
.Y(n_4798)
);

AND2x4_ASAP7_75t_L g4799 ( 
.A(n_4704),
.B(n_4613),
.Y(n_4799)
);

INVx3_ASAP7_75t_L g4800 ( 
.A(n_4705),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4711),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4726),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_4677),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4761),
.Y(n_4804)
);

INVx2_ASAP7_75t_L g4805 ( 
.A(n_4741),
.Y(n_4805)
);

INVx2_ASAP7_75t_SL g4806 ( 
.A(n_4700),
.Y(n_4806)
);

HB1xp67_ASAP7_75t_L g4807 ( 
.A(n_4750),
.Y(n_4807)
);

AND2x2_ASAP7_75t_L g4808 ( 
.A(n_4678),
.B(n_4561),
.Y(n_4808)
);

BUFx2_ASAP7_75t_L g4809 ( 
.A(n_4693),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4754),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4682),
.B(n_4637),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4713),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4772),
.B(n_4655),
.Y(n_4813)
);

OA21x2_ASAP7_75t_L g4814 ( 
.A1(n_4731),
.A2(n_4654),
.B(n_4622),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4738),
.B(n_4584),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4687),
.Y(n_4816)
);

BUFx12f_ASAP7_75t_L g4817 ( 
.A(n_4702),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4720),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4675),
.Y(n_4819)
);

AO31x2_ASAP7_75t_L g4820 ( 
.A1(n_4747),
.A2(n_4540),
.A3(n_350),
.B(n_348),
.Y(n_4820)
);

OR2x2_ASAP7_75t_L g4821 ( 
.A(n_4728),
.B(n_349),
.Y(n_4821)
);

AND2x2_ASAP7_75t_L g4822 ( 
.A(n_4703),
.B(n_351),
.Y(n_4822)
);

HB1xp67_ASAP7_75t_L g4823 ( 
.A(n_4689),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4745),
.Y(n_4824)
);

BUFx2_ASAP7_75t_L g4825 ( 
.A(n_4712),
.Y(n_4825)
);

OR2x2_ASAP7_75t_L g4826 ( 
.A(n_4664),
.B(n_352),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4673),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4783),
.Y(n_4828)
);

AOI22xp33_ASAP7_75t_SL g4829 ( 
.A1(n_4724),
.A2(n_4727),
.B1(n_4780),
.B2(n_4751),
.Y(n_4829)
);

AOI22xp33_ASAP7_75t_L g4830 ( 
.A1(n_4729),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_4830)
);

AND2x2_ASAP7_75t_L g4831 ( 
.A(n_4721),
.B(n_353),
.Y(n_4831)
);

AND2x2_ASAP7_75t_L g4832 ( 
.A(n_4717),
.B(n_355),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4771),
.Y(n_4833)
);

AND2x2_ASAP7_75t_L g4834 ( 
.A(n_4718),
.B(n_4736),
.Y(n_4834)
);

BUFx6f_ASAP7_75t_L g4835 ( 
.A(n_4669),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4734),
.B(n_355),
.Y(n_4836)
);

INVx2_ASAP7_75t_L g4837 ( 
.A(n_4786),
.Y(n_4837)
);

OA21x2_ASAP7_75t_L g4838 ( 
.A1(n_4697),
.A2(n_4759),
.B(n_4755),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4787),
.B(n_356),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_4770),
.Y(n_4840)
);

HB1xp67_ASAP7_75t_L g4841 ( 
.A(n_4685),
.Y(n_4841)
);

INVxp67_ASAP7_75t_R g4842 ( 
.A(n_4672),
.Y(n_4842)
);

INVx3_ASAP7_75t_L g4843 ( 
.A(n_4676),
.Y(n_4843)
);

OR2x2_ASAP7_75t_L g4844 ( 
.A(n_4714),
.B(n_357),
.Y(n_4844)
);

INVx3_ASAP7_75t_L g4845 ( 
.A(n_4669),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4752),
.B(n_357),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4753),
.Y(n_4847)
);

HB1xp67_ASAP7_75t_L g4848 ( 
.A(n_4784),
.Y(n_4848)
);

BUFx3_ASAP7_75t_L g4849 ( 
.A(n_4696),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4732),
.Y(n_4850)
);

NOR2xp67_ASAP7_75t_L g4851 ( 
.A(n_4699),
.B(n_359),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4684),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4666),
.B(n_359),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4762),
.Y(n_4854)
);

INVx2_ASAP7_75t_SL g4855 ( 
.A(n_4700),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4765),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4778),
.Y(n_4857)
);

BUFx6f_ASAP7_75t_L g4858 ( 
.A(n_4763),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4680),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4679),
.Y(n_4860)
);

OAI21x1_ASAP7_75t_L g4861 ( 
.A1(n_4683),
.A2(n_360),
.B(n_361),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4706),
.Y(n_4862)
);

HB1xp67_ASAP7_75t_L g4863 ( 
.A(n_4723),
.Y(n_4863)
);

AOI21x1_ASAP7_75t_L g4864 ( 
.A1(n_4674),
.A2(n_362),
.B(n_363),
.Y(n_4864)
);

OR2x2_ASAP7_75t_L g4865 ( 
.A(n_4742),
.B(n_362),
.Y(n_4865)
);

AO21x2_ASAP7_75t_L g4866 ( 
.A1(n_4691),
.A2(n_364),
.B(n_366),
.Y(n_4866)
);

INVx2_ASAP7_75t_L g4867 ( 
.A(n_4749),
.Y(n_4867)
);

OAI21x1_ASAP7_75t_L g4868 ( 
.A1(n_4716),
.A2(n_364),
.B(n_368),
.Y(n_4868)
);

INVx3_ASAP7_75t_L g4869 ( 
.A(n_4722),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_4779),
.Y(n_4870)
);

INVx2_ASAP7_75t_L g4871 ( 
.A(n_4695),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4782),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4768),
.Y(n_4873)
);

INVx3_ASAP7_75t_L g4874 ( 
.A(n_4730),
.Y(n_4874)
);

HB1xp67_ASAP7_75t_L g4875 ( 
.A(n_4769),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4776),
.Y(n_4876)
);

INVx5_ASAP7_75t_L g4877 ( 
.A(n_4681),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4774),
.Y(n_4878)
);

OAI21x1_ASAP7_75t_L g4879 ( 
.A1(n_4670),
.A2(n_368),
.B(n_369),
.Y(n_4879)
);

AOI21x1_ASAP7_75t_L g4880 ( 
.A1(n_4767),
.A2(n_369),
.B(n_370),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4686),
.B(n_370),
.Y(n_4881)
);

BUFx6f_ASAP7_75t_L g4882 ( 
.A(n_4733),
.Y(n_4882)
);

OAI21x1_ASAP7_75t_L g4883 ( 
.A1(n_4688),
.A2(n_371),
.B(n_372),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4746),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4756),
.Y(n_4885)
);

AND2x4_ASAP7_75t_L g4886 ( 
.A(n_4735),
.B(n_372),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4710),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4710),
.Y(n_4888)
);

BUFx2_ASAP7_75t_L g4889 ( 
.A(n_4698),
.Y(n_4889)
);

OAI21xp5_ASAP7_75t_L g4890 ( 
.A1(n_4739),
.A2(n_373),
.B(n_375),
.Y(n_4890)
);

INVx2_ASAP7_75t_L g4891 ( 
.A(n_4760),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4773),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4764),
.B(n_376),
.Y(n_4893)
);

HB1xp67_ASAP7_75t_SL g4894 ( 
.A(n_4743),
.Y(n_4894)
);

OA21x2_ASAP7_75t_L g4895 ( 
.A1(n_4740),
.A2(n_377),
.B(n_378),
.Y(n_4895)
);

BUFx3_ASAP7_75t_L g4896 ( 
.A(n_4748),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4785),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4757),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4775),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4708),
.Y(n_4900)
);

OAI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4758),
.A2(n_377),
.B(n_379),
.Y(n_4901)
);

INVx3_ASAP7_75t_L g4902 ( 
.A(n_4667),
.Y(n_4902)
);

BUFx2_ASAP7_75t_L g4903 ( 
.A(n_4766),
.Y(n_4903)
);

OR2x2_ASAP7_75t_L g4904 ( 
.A(n_4737),
.B(n_379),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4744),
.B(n_380),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4777),
.B(n_380),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4781),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4694),
.B(n_381),
.Y(n_4908)
);

BUFx3_ASAP7_75t_L g4909 ( 
.A(n_4696),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4668),
.B(n_381),
.Y(n_4910)
);

HB1xp67_ASAP7_75t_L g4911 ( 
.A(n_4668),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4707),
.Y(n_4912)
);

INVx2_ASAP7_75t_L g4913 ( 
.A(n_4709),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4709),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4707),
.Y(n_4915)
);

BUFx12f_ASAP7_75t_L g4916 ( 
.A(n_4702),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4665),
.B(n_382),
.Y(n_4917)
);

AO21x2_ASAP7_75t_L g4918 ( 
.A1(n_4731),
.A2(n_382),
.B(n_383),
.Y(n_4918)
);

INVx2_ASAP7_75t_SL g4919 ( 
.A(n_4671),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4803),
.B(n_384),
.Y(n_4920)
);

BUFx3_ASAP7_75t_L g4921 ( 
.A(n_4817),
.Y(n_4921)
);

A2O1A1Ixp33_ASAP7_75t_L g4922 ( 
.A1(n_4902),
.A2(n_4903),
.B(n_4900),
.C(n_4908),
.Y(n_4922)
);

AOI21xp33_ASAP7_75t_L g4923 ( 
.A1(n_4887),
.A2(n_386),
.B(n_387),
.Y(n_4923)
);

INVx3_ASAP7_75t_L g4924 ( 
.A(n_4800),
.Y(n_4924)
);

INVx3_ASAP7_75t_L g4925 ( 
.A(n_4843),
.Y(n_4925)
);

AOI21x1_ASAP7_75t_L g4926 ( 
.A1(n_4841),
.A2(n_386),
.B(n_387),
.Y(n_4926)
);

OAI22xp5_ASAP7_75t_L g4927 ( 
.A1(n_4829),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4907),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_4928)
);

A2O1A1Ixp33_ASAP7_75t_L g4929 ( 
.A1(n_4890),
.A2(n_4901),
.B(n_4844),
.C(n_4851),
.Y(n_4929)
);

INVxp67_ASAP7_75t_L g4930 ( 
.A(n_4789),
.Y(n_4930)
);

INVx2_ASAP7_75t_SL g4931 ( 
.A(n_4877),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4804),
.Y(n_4932)
);

OAI22xp5_ASAP7_75t_L g4933 ( 
.A1(n_4830),
.A2(n_4898),
.B1(n_4904),
.B2(n_4862),
.Y(n_4933)
);

BUFx6f_ASAP7_75t_L g4934 ( 
.A(n_4835),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4825),
.B(n_391),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4854),
.B(n_392),
.Y(n_4936)
);

AOI22xp33_ASAP7_75t_L g4937 ( 
.A1(n_4892),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4911),
.B(n_393),
.Y(n_4938)
);

HB1xp67_ASAP7_75t_L g4939 ( 
.A(n_4828),
.Y(n_4939)
);

OAI22xp5_ASAP7_75t_L g4940 ( 
.A1(n_4897),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_4940)
);

AOI21x1_ASAP7_75t_L g4941 ( 
.A1(n_4823),
.A2(n_395),
.B(n_397),
.Y(n_4941)
);

AOI22xp33_ASAP7_75t_L g4942 ( 
.A1(n_4856),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4807),
.Y(n_4943)
);

INVx3_ASAP7_75t_L g4944 ( 
.A(n_4877),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4809),
.B(n_398),
.Y(n_4945)
);

AND2x2_ASAP7_75t_L g4946 ( 
.A(n_4870),
.B(n_399),
.Y(n_4946)
);

NOR2xp67_ASAP7_75t_SL g4947 ( 
.A(n_4858),
.B(n_400),
.Y(n_4947)
);

AO31x2_ASAP7_75t_L g4948 ( 
.A1(n_4812),
.A2(n_402),
.A3(n_400),
.B(n_401),
.Y(n_4948)
);

INVx1_ASAP7_75t_SL g4949 ( 
.A(n_4889),
.Y(n_4949)
);

AOI21xp5_ASAP7_75t_L g4950 ( 
.A1(n_4859),
.A2(n_401),
.B(n_402),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4810),
.Y(n_4951)
);

AOI22xp5_ASAP7_75t_L g4952 ( 
.A1(n_4815),
.A2(n_4808),
.B1(n_4905),
.B2(n_4814),
.Y(n_4952)
);

AOI22xp33_ASAP7_75t_L g4953 ( 
.A1(n_4899),
.A2(n_406),
.B1(n_403),
.B2(n_405),
.Y(n_4953)
);

OAI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4839),
.A2(n_407),
.B1(n_403),
.B2(n_405),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4819),
.B(n_407),
.Y(n_4955)
);

AOI21xp33_ASAP7_75t_L g4956 ( 
.A1(n_4888),
.A2(n_408),
.B(n_409),
.Y(n_4956)
);

AND2x4_ASAP7_75t_SL g4957 ( 
.A(n_4858),
.B(n_410),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4834),
.B(n_411),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4818),
.Y(n_4959)
);

AOI22xp33_ASAP7_75t_SL g4960 ( 
.A1(n_4875),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4960)
);

AOI221xp5_ASAP7_75t_L g4961 ( 
.A1(n_4872),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4793),
.Y(n_4962)
);

BUFx2_ASAP7_75t_L g4963 ( 
.A(n_4795),
.Y(n_4963)
);

HB1xp67_ASAP7_75t_L g4964 ( 
.A(n_4863),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4867),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_4965)
);

INVx2_ASAP7_75t_L g4966 ( 
.A(n_4840),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4827),
.B(n_421),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_4824),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_4837),
.Y(n_4969)
);

OAI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4879),
.A2(n_422),
.B(n_423),
.Y(n_4970)
);

INVx3_ASAP7_75t_L g4971 ( 
.A(n_4874),
.Y(n_4971)
);

OAI22xp33_ASAP7_75t_L g4972 ( 
.A1(n_4821),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_4972)
);

AOI22xp33_ASAP7_75t_L g4973 ( 
.A1(n_4891),
.A2(n_430),
.B1(n_427),
.B2(n_429),
.Y(n_4973)
);

INVxp67_ASAP7_75t_L g4974 ( 
.A(n_4797),
.Y(n_4974)
);

OAI21x1_ASAP7_75t_L g4975 ( 
.A1(n_4860),
.A2(n_430),
.B(n_431),
.Y(n_4975)
);

NAND3xp33_ASAP7_75t_L g4976 ( 
.A(n_4848),
.B(n_432),
.C(n_433),
.Y(n_4976)
);

HB1xp67_ASAP7_75t_L g4977 ( 
.A(n_4847),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4788),
.B(n_434),
.Y(n_4978)
);

AOI221xp5_ASAP7_75t_L g4979 ( 
.A1(n_4884),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.C(n_438),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4816),
.B(n_4912),
.Y(n_4980)
);

BUFx2_ASAP7_75t_L g4981 ( 
.A(n_4792),
.Y(n_4981)
);

AOI22xp5_ASAP7_75t_L g4982 ( 
.A1(n_4906),
.A2(n_439),
.B1(n_436),
.B2(n_438),
.Y(n_4982)
);

AOI22xp33_ASAP7_75t_SL g4983 ( 
.A1(n_4813),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4915),
.B(n_442),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4796),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4895),
.A2(n_444),
.B(n_446),
.Y(n_4986)
);

OAI22xp5_ASAP7_75t_L g4987 ( 
.A1(n_4910),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4790),
.Y(n_4988)
);

AOI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4918),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_4989)
);

OAI221xp5_ASAP7_75t_L g4990 ( 
.A1(n_4880),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.C(n_453),
.Y(n_4990)
);

AOI22xp33_ASAP7_75t_L g4991 ( 
.A1(n_4857),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4913),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4914),
.Y(n_4993)
);

OAI22xp33_ASAP7_75t_L g4994 ( 
.A1(n_4896),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_4994)
);

BUFx2_ASAP7_75t_L g4995 ( 
.A(n_4919),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4801),
.Y(n_4996)
);

OAI21xp5_ASAP7_75t_L g4997 ( 
.A1(n_4864),
.A2(n_457),
.B(n_458),
.Y(n_4997)
);

OR2x2_ASAP7_75t_L g4998 ( 
.A(n_4833),
.B(n_458),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4850),
.Y(n_4999)
);

OAI22xp33_ASAP7_75t_L g5000 ( 
.A1(n_4826),
.A2(n_4842),
.B1(n_4885),
.B2(n_4865),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_4838),
.Y(n_5001)
);

BUFx3_ASAP7_75t_L g5002 ( 
.A(n_4916),
.Y(n_5002)
);

OAI22xp5_ASAP7_75t_L g5003 ( 
.A1(n_4799),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_5003)
);

OAI211xp5_ASAP7_75t_SL g5004 ( 
.A1(n_4846),
.A2(n_463),
.B(n_461),
.C(n_462),
.Y(n_5004)
);

AOI22xp33_ASAP7_75t_L g5005 ( 
.A1(n_4876),
.A2(n_467),
.B1(n_463),
.B2(n_466),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_4802),
.Y(n_5006)
);

AND2x4_ASAP7_75t_SL g5007 ( 
.A(n_4835),
.B(n_468),
.Y(n_5007)
);

AOI22xp33_ASAP7_75t_SL g5008 ( 
.A1(n_4811),
.A2(n_4866),
.B1(n_4881),
.B2(n_4893),
.Y(n_5008)
);

AOI22xp33_ASAP7_75t_SL g5009 ( 
.A1(n_4873),
.A2(n_471),
.B1(n_468),
.B2(n_469),
.Y(n_5009)
);

NAND2xp5_ASAP7_75t_L g5010 ( 
.A(n_4871),
.B(n_469),
.Y(n_5010)
);

AOI22xp5_ASAP7_75t_L g5011 ( 
.A1(n_4852),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_5011)
);

BUFx6f_ASAP7_75t_L g5012 ( 
.A(n_4849),
.Y(n_5012)
);

CKINVDCx20_ASAP7_75t_R g5013 ( 
.A(n_4909),
.Y(n_5013)
);

OAI211xp5_ASAP7_75t_SL g5014 ( 
.A1(n_4794),
.A2(n_475),
.B(n_472),
.C(n_473),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4805),
.Y(n_5015)
);

INVx2_ASAP7_75t_L g5016 ( 
.A(n_4791),
.Y(n_5016)
);

AND2x2_ASAP7_75t_L g5017 ( 
.A(n_4878),
.B(n_476),
.Y(n_5017)
);

AOI22xp5_ASAP7_75t_L g5018 ( 
.A1(n_4886),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_5018)
);

AOI22xp33_ASAP7_75t_SL g5019 ( 
.A1(n_4917),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_5019)
);

OAI21x1_ASAP7_75t_L g5020 ( 
.A1(n_4883),
.A2(n_481),
.B(n_483),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4820),
.Y(n_5021)
);

BUFx6f_ASAP7_75t_L g5022 ( 
.A(n_4882),
.Y(n_5022)
);

OAI22xp5_ASAP7_75t_L g5023 ( 
.A1(n_4894),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_5023)
);

AOI22xp33_ASAP7_75t_SL g5024 ( 
.A1(n_4836),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_5024)
);

AOI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4868),
.A2(n_488),
.B(n_489),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4820),
.Y(n_5026)
);

OAI22xp33_ASAP7_75t_L g5027 ( 
.A1(n_4882),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_SL g5028 ( 
.A(n_4806),
.B(n_490),
.Y(n_5028)
);

OA21x2_ASAP7_75t_L g5029 ( 
.A1(n_4861),
.A2(n_491),
.B(n_492),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4831),
.B(n_493),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4822),
.Y(n_5031)
);

AOI22xp33_ASAP7_75t_L g5032 ( 
.A1(n_4853),
.A2(n_4832),
.B1(n_4869),
.B2(n_4855),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4845),
.Y(n_5033)
);

AOI22xp33_ASAP7_75t_L g5034 ( 
.A1(n_4903),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.Y(n_5034)
);

INVx2_ASAP7_75t_SL g5035 ( 
.A(n_4877),
.Y(n_5035)
);

OAI211xp5_ASAP7_75t_SL g5036 ( 
.A1(n_4902),
.A2(n_500),
.B(n_497),
.C(n_498),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4825),
.B(n_500),
.Y(n_5037)
);

OAI21x1_ASAP7_75t_SL g5038 ( 
.A1(n_4792),
.A2(n_501),
.B(n_502),
.Y(n_5038)
);

AO31x2_ASAP7_75t_L g5039 ( 
.A1(n_4812),
.A2(n_503),
.A3(n_501),
.B(n_502),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4908),
.A2(n_503),
.B(n_504),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4789),
.B(n_505),
.Y(n_5041)
);

AOI22xp33_ASAP7_75t_L g5042 ( 
.A1(n_4903),
.A2(n_508),
.B1(n_505),
.B2(n_506),
.Y(n_5042)
);

INVx2_ASAP7_75t_L g5043 ( 
.A(n_4862),
.Y(n_5043)
);

AOI22xp33_ASAP7_75t_L g5044 ( 
.A1(n_4903),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4789),
.B(n_512),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4804),
.Y(n_5046)
);

OAI22xp5_ASAP7_75t_L g5047 ( 
.A1(n_4903),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_5047)
);

OAI22xp5_ASAP7_75t_L g5048 ( 
.A1(n_4903),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4862),
.Y(n_5049)
);

INVx4_ASAP7_75t_L g5050 ( 
.A(n_4817),
.Y(n_5050)
);

OAI22xp33_ASAP7_75t_L g5051 ( 
.A1(n_4903),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_5051)
);

OA21x2_ASAP7_75t_L g5052 ( 
.A1(n_4798),
.A2(n_518),
.B(n_519),
.Y(n_5052)
);

OAI22xp5_ASAP7_75t_L g5053 ( 
.A1(n_4903),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_5053)
);

AOI22xp33_ASAP7_75t_SL g5054 ( 
.A1(n_4903),
.A2(n_526),
.B1(n_523),
.B2(n_524),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4862),
.Y(n_5055)
);

AO31x2_ASAP7_75t_L g5056 ( 
.A1(n_4812),
.A2(n_528),
.A3(n_524),
.B(n_527),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4804),
.Y(n_5057)
);

HB1xp67_ASAP7_75t_L g5058 ( 
.A(n_4841),
.Y(n_5058)
);

AO221x2_ASAP7_75t_L g5059 ( 
.A1(n_4910),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.C(n_534),
.Y(n_5059)
);

HB1xp67_ASAP7_75t_L g5060 ( 
.A(n_4841),
.Y(n_5060)
);

AOI22xp33_ASAP7_75t_SL g5061 ( 
.A1(n_4903),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_5061)
);

AND2x2_ASAP7_75t_L g5062 ( 
.A(n_4789),
.B(n_538),
.Y(n_5062)
);

INVx2_ASAP7_75t_L g5063 ( 
.A(n_5043),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4932),
.Y(n_5064)
);

AOI22xp33_ASAP7_75t_L g5065 ( 
.A1(n_5059),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_5046),
.Y(n_5066)
);

INVx2_ASAP7_75t_L g5067 ( 
.A(n_5049),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_4963),
.B(n_539),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_5057),
.Y(n_5069)
);

HB1xp67_ASAP7_75t_L g5070 ( 
.A(n_4977),
.Y(n_5070)
);

NOR2x1_ASAP7_75t_SL g5071 ( 
.A(n_4920),
.B(n_542),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4974),
.B(n_542),
.Y(n_5072)
);

AND2x2_ASAP7_75t_SL g5073 ( 
.A(n_4952),
.B(n_544),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_5055),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4951),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_4981),
.B(n_544),
.Y(n_5076)
);

AND2x2_ASAP7_75t_L g5077 ( 
.A(n_4995),
.B(n_546),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4999),
.Y(n_5078)
);

BUFx3_ASAP7_75t_L g5079 ( 
.A(n_5013),
.Y(n_5079)
);

NAND3xp33_ASAP7_75t_L g5080 ( 
.A(n_4922),
.B(n_546),
.C(n_547),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4930),
.B(n_549),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_4925),
.B(n_550),
.Y(n_5082)
);

OR2x2_ASAP7_75t_L g5083 ( 
.A(n_4980),
.B(n_551),
.Y(n_5083)
);

INVx2_ASAP7_75t_L g5084 ( 
.A(n_4943),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_4924),
.B(n_4971),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4962),
.Y(n_5086)
);

INVxp67_ASAP7_75t_L g5087 ( 
.A(n_4949),
.Y(n_5087)
);

AND2x4_ASAP7_75t_SL g5088 ( 
.A(n_5012),
.B(n_5050),
.Y(n_5088)
);

AOI22xp33_ASAP7_75t_L g5089 ( 
.A1(n_4927),
.A2(n_555),
.B1(n_552),
.B2(n_553),
.Y(n_5089)
);

INVx2_ASAP7_75t_L g5090 ( 
.A(n_4966),
.Y(n_5090)
);

BUFx2_ASAP7_75t_L g5091 ( 
.A(n_4931),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_4968),
.Y(n_5092)
);

AND2x2_ASAP7_75t_L g5093 ( 
.A(n_5033),
.B(n_560),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_4939),
.B(n_561),
.Y(n_5094)
);

AND2x2_ASAP7_75t_L g5095 ( 
.A(n_5035),
.B(n_5058),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_4969),
.Y(n_5096)
);

AND2x2_ASAP7_75t_L g5097 ( 
.A(n_5060),
.B(n_562),
.Y(n_5097)
);

AND2x2_ASAP7_75t_L g5098 ( 
.A(n_5031),
.B(n_563),
.Y(n_5098)
);

INVxp67_ASAP7_75t_L g5099 ( 
.A(n_4936),
.Y(n_5099)
);

HB1xp67_ASAP7_75t_L g5100 ( 
.A(n_5021),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_4985),
.Y(n_5101)
);

HB1xp67_ASAP7_75t_L g5102 ( 
.A(n_5026),
.Y(n_5102)
);

HB1xp67_ASAP7_75t_L g5103 ( 
.A(n_4964),
.Y(n_5103)
);

BUFx2_ASAP7_75t_L g5104 ( 
.A(n_4921),
.Y(n_5104)
);

INVx2_ASAP7_75t_L g5105 ( 
.A(n_5001),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4996),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4984),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_L g5108 ( 
.A(n_4935),
.B(n_564),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_5006),
.Y(n_5109)
);

AOI22xp33_ASAP7_75t_L g5110 ( 
.A1(n_5008),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_5032),
.B(n_565),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_5015),
.Y(n_5112)
);

AOI22xp33_ASAP7_75t_L g5113 ( 
.A1(n_5052),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_5113)
);

AND2x2_ASAP7_75t_L g5114 ( 
.A(n_4958),
.B(n_567),
.Y(n_5114)
);

AND2x2_ASAP7_75t_L g5115 ( 
.A(n_5041),
.B(n_568),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4959),
.Y(n_5116)
);

OAI22xp5_ASAP7_75t_L g5117 ( 
.A1(n_4976),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_5117)
);

INVx2_ASAP7_75t_L g5118 ( 
.A(n_4992),
.Y(n_5118)
);

AND2x2_ASAP7_75t_L g5119 ( 
.A(n_5045),
.B(n_5062),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_4998),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_4945),
.B(n_4978),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_5037),
.B(n_570),
.Y(n_5122)
);

AOI22xp33_ASAP7_75t_L g5123 ( 
.A1(n_4990),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4955),
.Y(n_5124)
);

AOI22xp5_ASAP7_75t_L g5125 ( 
.A1(n_4933),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.Y(n_5125)
);

BUFx2_ASAP7_75t_L g5126 ( 
.A(n_5002),
.Y(n_5126)
);

OR2x2_ASAP7_75t_L g5127 ( 
.A(n_4938),
.B(n_576),
.Y(n_5127)
);

OR2x2_ASAP7_75t_L g5128 ( 
.A(n_4967),
.B(n_577),
.Y(n_5128)
);

AND2x2_ASAP7_75t_L g5129 ( 
.A(n_4946),
.B(n_578),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_5016),
.Y(n_5130)
);

OR2x2_ASAP7_75t_L g5131 ( 
.A(n_4988),
.B(n_578),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_4993),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_5022),
.B(n_579),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5010),
.Y(n_5134)
);

INVxp67_ASAP7_75t_SL g5135 ( 
.A(n_5000),
.Y(n_5135)
);

CKINVDCx6p67_ASAP7_75t_R g5136 ( 
.A(n_5012),
.Y(n_5136)
);

OR2x2_ASAP7_75t_L g5137 ( 
.A(n_4929),
.B(n_580),
.Y(n_5137)
);

BUFx3_ASAP7_75t_L g5138 ( 
.A(n_4934),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4948),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_5022),
.B(n_580),
.Y(n_5140)
);

NAND2x1_ASAP7_75t_L g5141 ( 
.A(n_4934),
.B(n_581),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4948),
.Y(n_5142)
);

NOR2xp33_ASAP7_75t_L g5143 ( 
.A(n_5030),
.B(n_581),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_5039),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_5017),
.B(n_583),
.Y(n_5145)
);

AOI22xp33_ASAP7_75t_L g5146 ( 
.A1(n_4986),
.A2(n_586),
.B1(n_583),
.B2(n_584),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_5040),
.B(n_584),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_5056),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_4957),
.B(n_587),
.Y(n_5149)
);

INVx2_ASAP7_75t_SL g5150 ( 
.A(n_5007),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4941),
.Y(n_5151)
);

AND2x4_ASAP7_75t_L g5152 ( 
.A(n_4975),
.B(n_589),
.Y(n_5152)
);

HB1xp67_ASAP7_75t_L g5153 ( 
.A(n_4926),
.Y(n_5153)
);

AOI22xp33_ASAP7_75t_L g5154 ( 
.A1(n_4997),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_5029),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_5020),
.Y(n_5156)
);

INVx3_ASAP7_75t_L g5157 ( 
.A(n_5038),
.Y(n_5157)
);

BUFx6f_ASAP7_75t_L g5158 ( 
.A(n_5028),
.Y(n_5158)
);

HB1xp67_ASAP7_75t_L g5159 ( 
.A(n_5003),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4972),
.Y(n_5160)
);

INVx2_ASAP7_75t_SL g5161 ( 
.A(n_5011),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_5018),
.Y(n_5162)
);

INVx2_ASAP7_75t_L g5163 ( 
.A(n_4987),
.Y(n_5163)
);

AND2x4_ASAP7_75t_L g5164 ( 
.A(n_4970),
.B(n_593),
.Y(n_5164)
);

BUFx2_ASAP7_75t_L g5165 ( 
.A(n_5047),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_5024),
.B(n_593),
.Y(n_5166)
);

INVx2_ASAP7_75t_L g5167 ( 
.A(n_5048),
.Y(n_5167)
);

INVx2_ASAP7_75t_SL g5168 ( 
.A(n_5053),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_5019),
.B(n_594),
.Y(n_5169)
);

INVxp67_ASAP7_75t_SL g5170 ( 
.A(n_4950),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_4940),
.Y(n_5171)
);

AND2x4_ASAP7_75t_L g5172 ( 
.A(n_4982),
.B(n_596),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4954),
.Y(n_5173)
);

AND2x2_ASAP7_75t_L g5174 ( 
.A(n_4947),
.B(n_597),
.Y(n_5174)
);

AND2x2_ASAP7_75t_L g5175 ( 
.A(n_5023),
.B(n_598),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_5051),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4965),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_4989),
.B(n_4960),
.Y(n_5178)
);

OR2x2_ASAP7_75t_L g5179 ( 
.A(n_4937),
.B(n_598),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5025),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_5004),
.Y(n_5181)
);

NOR2xp33_ASAP7_75t_L g5182 ( 
.A(n_5014),
.B(n_599),
.Y(n_5182)
);

INVx2_ASAP7_75t_L g5183 ( 
.A(n_4923),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4956),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4994),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_4979),
.B(n_5054),
.Y(n_5186)
);

AND2x2_ASAP7_75t_L g5187 ( 
.A(n_5061),
.B(n_601),
.Y(n_5187)
);

OR2x2_ASAP7_75t_L g5188 ( 
.A(n_5034),
.B(n_601),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4973),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_4961),
.B(n_602),
.Y(n_5190)
);

HB1xp67_ASAP7_75t_L g5191 ( 
.A(n_4991),
.Y(n_5191)
);

BUFx3_ASAP7_75t_L g5192 ( 
.A(n_5027),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_5042),
.B(n_602),
.Y(n_5193)
);

BUFx2_ASAP7_75t_L g5194 ( 
.A(n_5009),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_4953),
.Y(n_5195)
);

OR2x2_ASAP7_75t_L g5196 ( 
.A(n_5044),
.B(n_603),
.Y(n_5196)
);

INVx2_ASAP7_75t_SL g5197 ( 
.A(n_4983),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_4942),
.B(n_606),
.Y(n_5198)
);

AOI22xp33_ASAP7_75t_L g5199 ( 
.A1(n_5036),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_5005),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4928),
.Y(n_5201)
);

HB1xp67_ASAP7_75t_L g5202 ( 
.A(n_4977),
.Y(n_5202)
);

BUFx2_ASAP7_75t_L g5203 ( 
.A(n_4944),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_4974),
.B(n_611),
.Y(n_5204)
);

OR2x2_ASAP7_75t_L g5205 ( 
.A(n_4974),
.B(n_611),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_4974),
.B(n_612),
.Y(n_5206)
);

AND2x2_ASAP7_75t_L g5207 ( 
.A(n_4963),
.B(n_612),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_4974),
.B(n_613),
.Y(n_5208)
);

INVx2_ASAP7_75t_L g5209 ( 
.A(n_5043),
.Y(n_5209)
);

NAND2xp5_ASAP7_75t_L g5210 ( 
.A(n_4974),
.B(n_614),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4932),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_4932),
.Y(n_5212)
);

NAND3xp33_ASAP7_75t_L g5213 ( 
.A(n_4922),
.B(n_615),
.C(n_616),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_4944),
.B(n_615),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_4963),
.B(n_616),
.Y(n_5215)
);

AND2x2_ASAP7_75t_L g5216 ( 
.A(n_4963),
.B(n_617),
.Y(n_5216)
);

NAND3xp33_ASAP7_75t_SL g5217 ( 
.A(n_4922),
.B(n_618),
.C(n_619),
.Y(n_5217)
);

OR2x2_ASAP7_75t_L g5218 ( 
.A(n_4974),
.B(n_618),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_L g5219 ( 
.A(n_4974),
.B(n_619),
.Y(n_5219)
);

BUFx6f_ASAP7_75t_L g5220 ( 
.A(n_5012),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_5043),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4932),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_5064),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5066),
.Y(n_5224)
);

INVxp67_ASAP7_75t_SL g5225 ( 
.A(n_5153),
.Y(n_5225)
);

AND2x2_ASAP7_75t_L g5226 ( 
.A(n_5091),
.B(n_5203),
.Y(n_5226)
);

AND2x2_ASAP7_75t_L g5227 ( 
.A(n_5095),
.B(n_621),
.Y(n_5227)
);

AND2x2_ASAP7_75t_L g5228 ( 
.A(n_5085),
.B(n_623),
.Y(n_5228)
);

OR2x2_ASAP7_75t_L g5229 ( 
.A(n_5124),
.B(n_5107),
.Y(n_5229)
);

AND2x2_ASAP7_75t_L g5230 ( 
.A(n_5119),
.B(n_624),
.Y(n_5230)
);

AND2x2_ASAP7_75t_L g5231 ( 
.A(n_5087),
.B(n_625),
.Y(n_5231)
);

AND2x2_ASAP7_75t_L g5232 ( 
.A(n_5121),
.B(n_5068),
.Y(n_5232)
);

OR2x2_ASAP7_75t_L g5233 ( 
.A(n_5120),
.B(n_5155),
.Y(n_5233)
);

AND2x4_ASAP7_75t_L g5234 ( 
.A(n_5104),
.B(n_626),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_5099),
.B(n_627),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_5139),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_5126),
.Y(n_5237)
);

AND2x4_ASAP7_75t_L g5238 ( 
.A(n_5138),
.B(n_628),
.Y(n_5238)
);

HB1xp67_ASAP7_75t_L g5239 ( 
.A(n_5151),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_5069),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_5075),
.Y(n_5241)
);

AND2x2_ASAP7_75t_L g5242 ( 
.A(n_5207),
.B(n_629),
.Y(n_5242)
);

AND2x2_ASAP7_75t_L g5243 ( 
.A(n_5215),
.B(n_630),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_5216),
.B(n_630),
.Y(n_5244)
);

HB1xp67_ASAP7_75t_L g5245 ( 
.A(n_5103),
.Y(n_5245)
);

AND2x4_ASAP7_75t_L g5246 ( 
.A(n_5134),
.B(n_631),
.Y(n_5246)
);

AND2x2_ASAP7_75t_L g5247 ( 
.A(n_5159),
.B(n_632),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5086),
.Y(n_5248)
);

AND2x2_ASAP7_75t_L g5249 ( 
.A(n_5163),
.B(n_632),
.Y(n_5249)
);

INVx2_ASAP7_75t_L g5250 ( 
.A(n_5142),
.Y(n_5250)
);

AND2x2_ASAP7_75t_L g5251 ( 
.A(n_5173),
.B(n_633),
.Y(n_5251)
);

AND2x2_ASAP7_75t_L g5252 ( 
.A(n_5171),
.B(n_633),
.Y(n_5252)
);

AND2x2_ASAP7_75t_L g5253 ( 
.A(n_5097),
.B(n_5070),
.Y(n_5253)
);

NAND2x1p5_ASAP7_75t_L g5254 ( 
.A(n_5141),
.B(n_635),
.Y(n_5254)
);

OR2x2_ASAP7_75t_L g5255 ( 
.A(n_5101),
.B(n_636),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_5144),
.Y(n_5256)
);

AND2x2_ASAP7_75t_L g5257 ( 
.A(n_5202),
.B(n_636),
.Y(n_5257)
);

INVx3_ASAP7_75t_L g5258 ( 
.A(n_5079),
.Y(n_5258)
);

AND2x4_ASAP7_75t_L g5259 ( 
.A(n_5098),
.B(n_637),
.Y(n_5259)
);

AND2x2_ASAP7_75t_L g5260 ( 
.A(n_5156),
.B(n_637),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5106),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_L g5262 ( 
.A(n_5180),
.B(n_639),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_L g5263 ( 
.A(n_5165),
.B(n_640),
.Y(n_5263)
);

AND2x2_ASAP7_75t_L g5264 ( 
.A(n_5135),
.B(n_640),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_5170),
.B(n_641),
.Y(n_5265)
);

NAND2xp5_ASAP7_75t_L g5266 ( 
.A(n_5183),
.B(n_642),
.Y(n_5266)
);

NOR2xp33_ASAP7_75t_L g5267 ( 
.A(n_5157),
.B(n_643),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_5211),
.Y(n_5268)
);

OR2x2_ASAP7_75t_L g5269 ( 
.A(n_5212),
.B(n_643),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_5184),
.B(n_644),
.Y(n_5270)
);

HB1xp67_ASAP7_75t_L g5271 ( 
.A(n_5078),
.Y(n_5271)
);

INVx2_ASAP7_75t_L g5272 ( 
.A(n_5105),
.Y(n_5272)
);

INVx2_ASAP7_75t_L g5273 ( 
.A(n_5063),
.Y(n_5273)
);

AND2x2_ASAP7_75t_L g5274 ( 
.A(n_5093),
.B(n_5167),
.Y(n_5274)
);

NOR2x1_ASAP7_75t_L g5275 ( 
.A(n_5083),
.B(n_645),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_5222),
.B(n_646),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_5100),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5076),
.B(n_646),
.Y(n_5278)
);

AND2x2_ASAP7_75t_L g5279 ( 
.A(n_5077),
.B(n_647),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_SL g5280 ( 
.A(n_5158),
.B(n_648),
.Y(n_5280)
);

INVxp67_ASAP7_75t_L g5281 ( 
.A(n_5137),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5102),
.Y(n_5282)
);

HB1xp67_ASAP7_75t_L g5283 ( 
.A(n_5185),
.Y(n_5283)
);

NOR2xp33_ASAP7_75t_L g5284 ( 
.A(n_5181),
.B(n_651),
.Y(n_5284)
);

OR2x2_ASAP7_75t_L g5285 ( 
.A(n_5160),
.B(n_651),
.Y(n_5285)
);

AND2x2_ASAP7_75t_L g5286 ( 
.A(n_5168),
.B(n_652),
.Y(n_5286)
);

BUFx2_ASAP7_75t_L g5287 ( 
.A(n_5214),
.Y(n_5287)
);

AND2x2_ASAP7_75t_L g5288 ( 
.A(n_5082),
.B(n_5177),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_5094),
.B(n_653),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_5131),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_5176),
.B(n_653),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5132),
.Y(n_5292)
);

NOR2xp67_ASAP7_75t_L g5293 ( 
.A(n_5080),
.B(n_654),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5205),
.Y(n_5294)
);

OR2x2_ASAP7_75t_L g5295 ( 
.A(n_5218),
.B(n_654),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5067),
.Y(n_5296)
);

NOR2xp33_ASAP7_75t_SL g5297 ( 
.A(n_5213),
.B(n_655),
.Y(n_5297)
);

AND2x2_ASAP7_75t_L g5298 ( 
.A(n_5115),
.B(n_656),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_5074),
.Y(n_5299)
);

INVx2_ASAP7_75t_L g5300 ( 
.A(n_5209),
.Y(n_5300)
);

NOR2x1_ASAP7_75t_SL g5301 ( 
.A(n_5158),
.B(n_657),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_5221),
.Y(n_5302)
);

AND2x2_ASAP7_75t_L g5303 ( 
.A(n_5071),
.B(n_657),
.Y(n_5303)
);

AND2x4_ASAP7_75t_L g5304 ( 
.A(n_5150),
.B(n_658),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_5162),
.B(n_659),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_5072),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_5096),
.Y(n_5307)
);

NAND2xp5_ASAP7_75t_SL g5308 ( 
.A(n_5204),
.B(n_5206),
.Y(n_5308)
);

INVxp67_ASAP7_75t_L g5309 ( 
.A(n_5191),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5208),
.Y(n_5310)
);

AND2x4_ASAP7_75t_SL g5311 ( 
.A(n_5133),
.B(n_659),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_5210),
.Y(n_5312)
);

OR2x2_ASAP7_75t_L g5313 ( 
.A(n_5200),
.B(n_5219),
.Y(n_5313)
);

BUFx2_ASAP7_75t_SL g5314 ( 
.A(n_5114),
.Y(n_5314)
);

INVx2_ASAP7_75t_L g5315 ( 
.A(n_5118),
.Y(n_5315)
);

INVxp67_ASAP7_75t_SL g5316 ( 
.A(n_5192),
.Y(n_5316)
);

AND2x4_ASAP7_75t_SL g5317 ( 
.A(n_5140),
.B(n_660),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_5081),
.B(n_660),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5109),
.Y(n_5319)
);

NAND2xp5_ASAP7_75t_L g5320 ( 
.A(n_5127),
.B(n_661),
.Y(n_5320)
);

INVxp67_ASAP7_75t_L g5321 ( 
.A(n_5194),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_5112),
.Y(n_5322)
);

AND2x2_ASAP7_75t_L g5323 ( 
.A(n_5111),
.B(n_5129),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_5201),
.B(n_661),
.Y(n_5324)
);

NAND3xp33_ASAP7_75t_SL g5325 ( 
.A(n_5110),
.B(n_663),
.C(n_664),
.Y(n_5325)
);

AND2x2_ASAP7_75t_SL g5326 ( 
.A(n_5164),
.B(n_663),
.Y(n_5326)
);

OAI221xp5_ASAP7_75t_SL g5327 ( 
.A1(n_5065),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.C(n_667),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_5189),
.B(n_668),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_5128),
.B(n_669),
.Y(n_5329)
);

AND2x4_ASAP7_75t_L g5330 ( 
.A(n_5152),
.B(n_669),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5116),
.Y(n_5331)
);

AND2x4_ASAP7_75t_SL g5332 ( 
.A(n_5145),
.B(n_670),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_5195),
.Y(n_5333)
);

HB1xp67_ASAP7_75t_L g5334 ( 
.A(n_5108),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_5161),
.B(n_671),
.Y(n_5335)
);

AND2x2_ASAP7_75t_L g5336 ( 
.A(n_5143),
.B(n_5122),
.Y(n_5336)
);

AND2x2_ASAP7_75t_L g5337 ( 
.A(n_5175),
.B(n_672),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5090),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5092),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5130),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_5174),
.B(n_672),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5125),
.B(n_673),
.Y(n_5342)
);

INVx4_ASAP7_75t_L g5343 ( 
.A(n_5149),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_SL g5344 ( 
.A(n_5172),
.B(n_674),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_5147),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5178),
.Y(n_5346)
);

AND2x2_ASAP7_75t_L g5347 ( 
.A(n_5197),
.B(n_675),
.Y(n_5347)
);

INVx2_ASAP7_75t_L g5348 ( 
.A(n_5186),
.Y(n_5348)
);

INVx2_ASAP7_75t_L g5349 ( 
.A(n_5169),
.Y(n_5349)
);

AND2x2_ASAP7_75t_L g5350 ( 
.A(n_5166),
.B(n_676),
.Y(n_5350)
);

AND2x2_ASAP7_75t_L g5351 ( 
.A(n_5187),
.B(n_677),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5190),
.Y(n_5352)
);

AND2x2_ASAP7_75t_L g5353 ( 
.A(n_5182),
.B(n_678),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5198),
.Y(n_5354)
);

HB1xp67_ASAP7_75t_L g5355 ( 
.A(n_5117),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_5113),
.B(n_680),
.Y(n_5356)
);

AND2x4_ASAP7_75t_SL g5357 ( 
.A(n_5193),
.B(n_681),
.Y(n_5357)
);

NAND2xp5_ASAP7_75t_L g5358 ( 
.A(n_5217),
.B(n_682),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_5179),
.Y(n_5359)
);

AND2x4_ASAP7_75t_L g5360 ( 
.A(n_5188),
.B(n_682),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5196),
.Y(n_5361)
);

AND2x2_ASAP7_75t_L g5362 ( 
.A(n_5154),
.B(n_683),
.Y(n_5362)
);

AND2x2_ASAP7_75t_L g5363 ( 
.A(n_5123),
.B(n_5089),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5146),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_5199),
.Y(n_5365)
);

NOR2xp33_ASAP7_75t_L g5366 ( 
.A(n_5136),
.B(n_683),
.Y(n_5366)
);

INVx2_ASAP7_75t_L g5367 ( 
.A(n_5148),
.Y(n_5367)
);

INVxp67_ASAP7_75t_SL g5368 ( 
.A(n_5153),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_5064),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_5064),
.Y(n_5370)
);

AND2x2_ASAP7_75t_L g5371 ( 
.A(n_5091),
.B(n_684),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5099),
.B(n_685),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_SL g5373 ( 
.A(n_5087),
.B(n_686),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_5099),
.B(n_687),
.Y(n_5374)
);

INVxp67_ASAP7_75t_L g5375 ( 
.A(n_5091),
.Y(n_5375)
);

AND2x2_ASAP7_75t_L g5376 ( 
.A(n_5091),
.B(n_687),
.Y(n_5376)
);

AND2x2_ASAP7_75t_L g5377 ( 
.A(n_5091),
.B(n_688),
.Y(n_5377)
);

NOR2x1_ASAP7_75t_L g5378 ( 
.A(n_5104),
.B(n_689),
.Y(n_5378)
);

AND2x2_ASAP7_75t_L g5379 ( 
.A(n_5091),
.B(n_689),
.Y(n_5379)
);

NOR3xp33_ASAP7_75t_L g5380 ( 
.A(n_5217),
.B(n_690),
.C(n_691),
.Y(n_5380)
);

AND2x2_ASAP7_75t_L g5381 ( 
.A(n_5091),
.B(n_691),
.Y(n_5381)
);

AND2x2_ASAP7_75t_L g5382 ( 
.A(n_5091),
.B(n_692),
.Y(n_5382)
);

AND2x2_ASAP7_75t_L g5383 ( 
.A(n_5091),
.B(n_692),
.Y(n_5383)
);

AND2x4_ASAP7_75t_SL g5384 ( 
.A(n_5136),
.B(n_693),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5148),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_5099),
.B(n_693),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_5064),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_5099),
.B(n_694),
.Y(n_5388)
);

HB1xp67_ASAP7_75t_L g5389 ( 
.A(n_5153),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_5064),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5091),
.B(n_695),
.Y(n_5391)
);

INVx2_ASAP7_75t_SL g5392 ( 
.A(n_5088),
.Y(n_5392)
);

OR2x2_ASAP7_75t_L g5393 ( 
.A(n_5084),
.B(n_696),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_5148),
.Y(n_5394)
);

AND2x2_ASAP7_75t_SL g5395 ( 
.A(n_5073),
.B(n_696),
.Y(n_5395)
);

INVx4_ASAP7_75t_L g5396 ( 
.A(n_5220),
.Y(n_5396)
);

AND2x2_ASAP7_75t_L g5397 ( 
.A(n_5091),
.B(n_697),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5064),
.Y(n_5398)
);

INVx2_ASAP7_75t_L g5399 ( 
.A(n_5148),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_5148),
.Y(n_5400)
);

OR2x6_ASAP7_75t_SL g5401 ( 
.A(n_5137),
.B(n_697),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_L g5402 ( 
.A(n_5099),
.B(n_700),
.Y(n_5402)
);

HB1xp67_ASAP7_75t_L g5403 ( 
.A(n_5153),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5099),
.B(n_701),
.Y(n_5404)
);

AND2x2_ASAP7_75t_L g5405 ( 
.A(n_5091),
.B(n_702),
.Y(n_5405)
);

AND2x2_ASAP7_75t_L g5406 ( 
.A(n_5091),
.B(n_702),
.Y(n_5406)
);

AND2x2_ASAP7_75t_L g5407 ( 
.A(n_5091),
.B(n_703),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5064),
.Y(n_5408)
);

INVx2_ASAP7_75t_L g5409 ( 
.A(n_5148),
.Y(n_5409)
);

AND2x2_ASAP7_75t_L g5410 ( 
.A(n_5091),
.B(n_704),
.Y(n_5410)
);

INVx2_ASAP7_75t_L g5411 ( 
.A(n_5148),
.Y(n_5411)
);

INVx2_ASAP7_75t_SL g5412 ( 
.A(n_5258),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5271),
.Y(n_5413)
);

HB1xp67_ASAP7_75t_L g5414 ( 
.A(n_5237),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5229),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5233),
.Y(n_5416)
);

OAI221xp5_ASAP7_75t_L g5417 ( 
.A1(n_5348),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.C(n_708),
.Y(n_5417)
);

AO21x2_ASAP7_75t_L g5418 ( 
.A1(n_5225),
.A2(n_705),
.B(n_708),
.Y(n_5418)
);

NAND4xp25_ASAP7_75t_L g5419 ( 
.A(n_5375),
.B(n_711),
.C(n_709),
.D(n_710),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_5223),
.Y(n_5420)
);

AND2x2_ASAP7_75t_L g5421 ( 
.A(n_5232),
.B(n_5314),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_5287),
.Y(n_5422)
);

AND2x4_ASAP7_75t_L g5423 ( 
.A(n_5343),
.B(n_712),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5224),
.Y(n_5424)
);

AOI22xp33_ASAP7_75t_L g5425 ( 
.A1(n_5346),
.A2(n_715),
.B1(n_713),
.B2(n_714),
.Y(n_5425)
);

NAND2xp5_ASAP7_75t_L g5426 ( 
.A(n_5345),
.B(n_715),
.Y(n_5426)
);

INVx2_ASAP7_75t_SL g5427 ( 
.A(n_5384),
.Y(n_5427)
);

OAI22xp5_ASAP7_75t_L g5428 ( 
.A1(n_5321),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_5428)
);

OAI211xp5_ASAP7_75t_SL g5429 ( 
.A1(n_5355),
.A2(n_718),
.B(n_716),
.C(n_717),
.Y(n_5429)
);

AND2x2_ASAP7_75t_L g5430 ( 
.A(n_5253),
.B(n_719),
.Y(n_5430)
);

INVx4_ASAP7_75t_L g5431 ( 
.A(n_5234),
.Y(n_5431)
);

OAI31xp33_ASAP7_75t_L g5432 ( 
.A1(n_5281),
.A2(n_722),
.A3(n_720),
.B(n_721),
.Y(n_5432)
);

NOR3xp33_ASAP7_75t_SL g5433 ( 
.A(n_5368),
.B(n_721),
.C(n_722),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_L g5434 ( 
.A(n_5334),
.B(n_5264),
.Y(n_5434)
);

INVxp67_ASAP7_75t_L g5435 ( 
.A(n_5401),
.Y(n_5435)
);

AOI22xp5_ASAP7_75t_L g5436 ( 
.A1(n_5297),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_5436)
);

AOI22xp5_ASAP7_75t_L g5437 ( 
.A1(n_5395),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_5437)
);

AND2x2_ASAP7_75t_L g5438 ( 
.A(n_5226),
.B(n_726),
.Y(n_5438)
);

OAI33xp33_ASAP7_75t_L g5439 ( 
.A1(n_5309),
.A2(n_729),
.A3(n_731),
.B1(n_727),
.B2(n_728),
.B3(n_730),
.Y(n_5439)
);

INVx3_ASAP7_75t_L g5440 ( 
.A(n_5396),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5240),
.Y(n_5441)
);

NAND2xp5_ASAP7_75t_L g5442 ( 
.A(n_5247),
.B(n_727),
.Y(n_5442)
);

NAND3x1_ASAP7_75t_L g5443 ( 
.A(n_5263),
.B(n_728),
.C(n_729),
.Y(n_5443)
);

OAI321xp33_ASAP7_75t_L g5444 ( 
.A1(n_5327),
.A2(n_734),
.A3(n_736),
.B1(n_732),
.B2(n_733),
.C(n_735),
.Y(n_5444)
);

AND2x2_ASAP7_75t_L g5445 ( 
.A(n_5306),
.B(n_732),
.Y(n_5445)
);

AOI33xp33_ASAP7_75t_L g5446 ( 
.A1(n_5352),
.A2(n_1716),
.A3(n_1714),
.B1(n_1717),
.B2(n_1715),
.B3(n_1713),
.Y(n_5446)
);

NAND2xp33_ASAP7_75t_R g5447 ( 
.A(n_5358),
.B(n_734),
.Y(n_5447)
);

BUFx2_ASAP7_75t_L g5448 ( 
.A(n_5392),
.Y(n_5448)
);

NAND3xp33_ASAP7_75t_L g5449 ( 
.A(n_5380),
.B(n_736),
.C(n_737),
.Y(n_5449)
);

OR2x2_ASAP7_75t_L g5450 ( 
.A(n_5313),
.B(n_5283),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5310),
.B(n_738),
.Y(n_5451)
);

BUFx3_ASAP7_75t_L g5452 ( 
.A(n_5332),
.Y(n_5452)
);

INVx2_ASAP7_75t_L g5453 ( 
.A(n_5393),
.Y(n_5453)
);

AND2x4_ASAP7_75t_L g5454 ( 
.A(n_5274),
.B(n_5288),
.Y(n_5454)
);

AND2x2_ASAP7_75t_L g5455 ( 
.A(n_5312),
.B(n_740),
.Y(n_5455)
);

INVx3_ASAP7_75t_L g5456 ( 
.A(n_5304),
.Y(n_5456)
);

INVx3_ASAP7_75t_L g5457 ( 
.A(n_5238),
.Y(n_5457)
);

AND2x2_ASAP7_75t_L g5458 ( 
.A(n_5227),
.B(n_741),
.Y(n_5458)
);

AOI211x1_ASAP7_75t_L g5459 ( 
.A1(n_5373),
.A2(n_744),
.B(n_742),
.C(n_743),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5241),
.Y(n_5460)
);

OR2x2_ASAP7_75t_L g5461 ( 
.A(n_5245),
.B(n_1708),
.Y(n_5461)
);

BUFx2_ASAP7_75t_L g5462 ( 
.A(n_5378),
.Y(n_5462)
);

AND2x2_ASAP7_75t_L g5463 ( 
.A(n_5230),
.B(n_742),
.Y(n_5463)
);

INVxp67_ASAP7_75t_L g5464 ( 
.A(n_5316),
.Y(n_5464)
);

HB1xp67_ASAP7_75t_L g5465 ( 
.A(n_5389),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5248),
.Y(n_5466)
);

OAI221xp5_ASAP7_75t_L g5467 ( 
.A1(n_5293),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.C(n_746),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_L g5468 ( 
.A(n_5354),
.B(n_745),
.Y(n_5468)
);

INVxp67_ASAP7_75t_SL g5469 ( 
.A(n_5275),
.Y(n_5469)
);

AOI221xp5_ASAP7_75t_L g5470 ( 
.A1(n_5403),
.A2(n_748),
.B1(n_746),
.B2(n_747),
.C(n_749),
.Y(n_5470)
);

OAI33xp33_ASAP7_75t_L g5471 ( 
.A1(n_5277),
.A2(n_5282),
.A3(n_5365),
.B1(n_5265),
.B2(n_5364),
.B3(n_5342),
.Y(n_5471)
);

AND2x2_ASAP7_75t_L g5472 ( 
.A(n_5294),
.B(n_748),
.Y(n_5472)
);

OAI211xp5_ASAP7_75t_SL g5473 ( 
.A1(n_5308),
.A2(n_752),
.B(n_750),
.C(n_751),
.Y(n_5473)
);

HB1xp67_ASAP7_75t_L g5474 ( 
.A(n_5239),
.Y(n_5474)
);

INVx2_ASAP7_75t_L g5475 ( 
.A(n_5367),
.Y(n_5475)
);

NOR2x1_ASAP7_75t_SL g5476 ( 
.A(n_5255),
.B(n_750),
.Y(n_5476)
);

AOI221xp5_ASAP7_75t_L g5477 ( 
.A1(n_5333),
.A2(n_755),
.B1(n_753),
.B2(n_754),
.C(n_756),
.Y(n_5477)
);

INVx2_ASAP7_75t_L g5478 ( 
.A(n_5385),
.Y(n_5478)
);

AO21x2_ASAP7_75t_L g5479 ( 
.A1(n_5328),
.A2(n_757),
.B(n_758),
.Y(n_5479)
);

OR2x2_ASAP7_75t_L g5480 ( 
.A(n_5290),
.B(n_1711),
.Y(n_5480)
);

BUFx2_ASAP7_75t_L g5481 ( 
.A(n_5371),
.Y(n_5481)
);

INVx2_ASAP7_75t_L g5482 ( 
.A(n_5394),
.Y(n_5482)
);

INVxp67_ASAP7_75t_L g5483 ( 
.A(n_5267),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5261),
.Y(n_5484)
);

OR2x2_ASAP7_75t_L g5485 ( 
.A(n_5276),
.B(n_1712),
.Y(n_5485)
);

NOR2xp33_ASAP7_75t_L g5486 ( 
.A(n_5336),
.B(n_5266),
.Y(n_5486)
);

HB1xp67_ASAP7_75t_L g5487 ( 
.A(n_5268),
.Y(n_5487)
);

OR2x2_ASAP7_75t_L g5488 ( 
.A(n_5262),
.B(n_1712),
.Y(n_5488)
);

AND2x2_ASAP7_75t_L g5489 ( 
.A(n_5376),
.B(n_759),
.Y(n_5489)
);

AND2x4_ASAP7_75t_L g5490 ( 
.A(n_5377),
.B(n_760),
.Y(n_5490)
);

AND2x2_ASAP7_75t_L g5491 ( 
.A(n_5379),
.B(n_761),
.Y(n_5491)
);

AND2x4_ASAP7_75t_L g5492 ( 
.A(n_5381),
.B(n_761),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_5369),
.Y(n_5493)
);

AND2x4_ASAP7_75t_L g5494 ( 
.A(n_5382),
.B(n_5383),
.Y(n_5494)
);

INVx2_ASAP7_75t_L g5495 ( 
.A(n_5399),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5251),
.B(n_763),
.Y(n_5496)
);

AOI22xp33_ASAP7_75t_SL g5497 ( 
.A1(n_5326),
.A2(n_766),
.B1(n_763),
.B2(n_764),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5370),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_5400),
.Y(n_5499)
);

AND2x2_ASAP7_75t_L g5500 ( 
.A(n_5391),
.B(n_767),
.Y(n_5500)
);

INVx4_ASAP7_75t_L g5501 ( 
.A(n_5278),
.Y(n_5501)
);

HB1xp67_ASAP7_75t_L g5502 ( 
.A(n_5387),
.Y(n_5502)
);

BUFx2_ASAP7_75t_L g5503 ( 
.A(n_5397),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5252),
.B(n_768),
.Y(n_5504)
);

AOI31xp33_ASAP7_75t_L g5505 ( 
.A1(n_5254),
.A2(n_780),
.A3(n_788),
.B(n_769),
.Y(n_5505)
);

OAI221xp5_ASAP7_75t_SL g5506 ( 
.A1(n_5356),
.A2(n_5353),
.B1(n_5363),
.B2(n_5270),
.C(n_5303),
.Y(n_5506)
);

OR2x2_ASAP7_75t_L g5507 ( 
.A(n_5390),
.B(n_1704),
.Y(n_5507)
);

INVx2_ASAP7_75t_L g5508 ( 
.A(n_5409),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5398),
.Y(n_5509)
);

NAND3xp33_ASAP7_75t_L g5510 ( 
.A(n_5284),
.B(n_772),
.C(n_773),
.Y(n_5510)
);

AND2x2_ASAP7_75t_L g5511 ( 
.A(n_5405),
.B(n_775),
.Y(n_5511)
);

AOI33xp33_ASAP7_75t_L g5512 ( 
.A1(n_5231),
.A2(n_5286),
.A3(n_5359),
.B1(n_5337),
.B2(n_5361),
.B3(n_5362),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5411),
.Y(n_5513)
);

INVxp67_ASAP7_75t_L g5514 ( 
.A(n_5285),
.Y(n_5514)
);

AND2x2_ASAP7_75t_L g5515 ( 
.A(n_5406),
.B(n_5407),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5408),
.Y(n_5516)
);

INVx2_ASAP7_75t_L g5517 ( 
.A(n_5236),
.Y(n_5517)
);

OAI221xp5_ASAP7_75t_SL g5518 ( 
.A1(n_5351),
.A2(n_779),
.B1(n_777),
.B2(n_778),
.C(n_781),
.Y(n_5518)
);

INVx1_ASAP7_75t_SL g5519 ( 
.A(n_5311),
.Y(n_5519)
);

AND2x2_ASAP7_75t_L g5520 ( 
.A(n_5410),
.B(n_782),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5250),
.Y(n_5521)
);

AOI22xp33_ASAP7_75t_L g5522 ( 
.A1(n_5272),
.A2(n_5349),
.B1(n_5325),
.B2(n_5300),
.Y(n_5522)
);

INVx1_ASAP7_75t_SL g5523 ( 
.A(n_5317),
.Y(n_5523)
);

HB1xp67_ASAP7_75t_L g5524 ( 
.A(n_5269),
.Y(n_5524)
);

NAND2xp5_ASAP7_75t_L g5525 ( 
.A(n_5257),
.B(n_5249),
.Y(n_5525)
);

AND2x2_ASAP7_75t_L g5526 ( 
.A(n_5228),
.B(n_783),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_5256),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_5260),
.B(n_785),
.Y(n_5528)
);

OAI33xp33_ASAP7_75t_L g5529 ( 
.A1(n_5324),
.A2(n_5335),
.A3(n_5344),
.B1(n_5331),
.B2(n_5322),
.B3(n_5319),
.Y(n_5529)
);

AOI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_5323),
.A2(n_789),
.B1(n_786),
.B2(n_787),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5291),
.B(n_790),
.Y(n_5531)
);

INVx3_ASAP7_75t_L g5532 ( 
.A(n_5246),
.Y(n_5532)
);

INVx2_ASAP7_75t_L g5533 ( 
.A(n_5307),
.Y(n_5533)
);

NAND4xp25_ASAP7_75t_L g5534 ( 
.A(n_5366),
.B(n_794),
.C(n_792),
.D(n_793),
.Y(n_5534)
);

NAND3xp33_ASAP7_75t_L g5535 ( 
.A(n_5280),
.B(n_793),
.C(n_796),
.Y(n_5535)
);

NOR3xp33_ASAP7_75t_L g5536 ( 
.A(n_5235),
.B(n_796),
.C(n_797),
.Y(n_5536)
);

INVxp67_ASAP7_75t_L g5537 ( 
.A(n_5301),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5292),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_5372),
.Y(n_5539)
);

OAI33xp33_ASAP7_75t_L g5540 ( 
.A1(n_5318),
.A2(n_802),
.A3(n_804),
.B1(n_797),
.B2(n_801),
.B3(n_803),
.Y(n_5540)
);

OAI321xp33_ASAP7_75t_L g5541 ( 
.A1(n_5347),
.A2(n_805),
.A3(n_807),
.B1(n_803),
.B2(n_804),
.C(n_806),
.Y(n_5541)
);

OAI33xp33_ASAP7_75t_L g5542 ( 
.A1(n_5289),
.A2(n_810),
.A3(n_812),
.B1(n_808),
.B2(n_809),
.B3(n_811),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_5501),
.B(n_5279),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5487),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_5469),
.B(n_5350),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_L g5546 ( 
.A(n_5524),
.B(n_5242),
.Y(n_5546)
);

INVx1_ASAP7_75t_SL g5547 ( 
.A(n_5481),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_5502),
.Y(n_5548)
);

INVx2_ASAP7_75t_L g5549 ( 
.A(n_5454),
.Y(n_5549)
);

AND2x4_ASAP7_75t_L g5550 ( 
.A(n_5431),
.B(n_5298),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_5421),
.B(n_5243),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5426),
.Y(n_5552)
);

OR2x2_ASAP7_75t_L g5553 ( 
.A(n_5450),
.B(n_5374),
.Y(n_5553)
);

AND2x2_ASAP7_75t_L g5554 ( 
.A(n_5503),
.B(n_5244),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_5515),
.B(n_5341),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5465),
.Y(n_5556)
);

AOI22xp33_ASAP7_75t_L g5557 ( 
.A1(n_5471),
.A2(n_5273),
.B1(n_5299),
.B2(n_5296),
.Y(n_5557)
);

AND2x2_ASAP7_75t_L g5558 ( 
.A(n_5448),
.B(n_5330),
.Y(n_5558)
);

HB1xp67_ASAP7_75t_L g5559 ( 
.A(n_5414),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5461),
.Y(n_5560)
);

INVx5_ASAP7_75t_SL g5561 ( 
.A(n_5423),
.Y(n_5561)
);

NOR2xp33_ASAP7_75t_L g5562 ( 
.A(n_5462),
.B(n_5329),
.Y(n_5562)
);

AND2x2_ASAP7_75t_L g5563 ( 
.A(n_5494),
.B(n_5295),
.Y(n_5563)
);

NOR2x1_ASAP7_75t_R g5564 ( 
.A(n_5452),
.B(n_5320),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5521),
.Y(n_5565)
);

AND2x2_ASAP7_75t_L g5566 ( 
.A(n_5412),
.B(n_5259),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_5456),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5476),
.Y(n_5568)
);

INVxp67_ASAP7_75t_SL g5569 ( 
.A(n_5435),
.Y(n_5569)
);

HB1xp67_ASAP7_75t_L g5570 ( 
.A(n_5464),
.Y(n_5570)
);

HB1xp67_ASAP7_75t_L g5571 ( 
.A(n_5422),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_5527),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_5420),
.Y(n_5573)
);

OR2x2_ASAP7_75t_L g5574 ( 
.A(n_5434),
.B(n_5386),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5424),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_5486),
.B(n_5388),
.Y(n_5576)
);

AND2x2_ASAP7_75t_L g5577 ( 
.A(n_5440),
.B(n_5402),
.Y(n_5577)
);

INVxp67_ASAP7_75t_L g5578 ( 
.A(n_5447),
.Y(n_5578)
);

OR2x2_ASAP7_75t_L g5579 ( 
.A(n_5415),
.B(n_5404),
.Y(n_5579)
);

AND2x2_ASAP7_75t_L g5580 ( 
.A(n_5457),
.B(n_5438),
.Y(n_5580)
);

HB1xp67_ASAP7_75t_L g5581 ( 
.A(n_5418),
.Y(n_5581)
);

AND2x4_ASAP7_75t_L g5582 ( 
.A(n_5427),
.B(n_5532),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5441),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5512),
.B(n_5305),
.Y(n_5584)
);

AND2x2_ASAP7_75t_L g5585 ( 
.A(n_5430),
.B(n_5360),
.Y(n_5585)
);

HB1xp67_ASAP7_75t_L g5586 ( 
.A(n_5474),
.Y(n_5586)
);

NOR2x1_ASAP7_75t_L g5587 ( 
.A(n_5419),
.B(n_5302),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5460),
.Y(n_5588)
);

NAND2xp5_ASAP7_75t_L g5589 ( 
.A(n_5479),
.B(n_5357),
.Y(n_5589)
);

OR2x2_ASAP7_75t_L g5590 ( 
.A(n_5539),
.B(n_5416),
.Y(n_5590)
);

INVx6_ASAP7_75t_L g5591 ( 
.A(n_5490),
.Y(n_5591)
);

NAND3xp33_ASAP7_75t_L g5592 ( 
.A(n_5433),
.B(n_5339),
.C(n_5338),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5466),
.Y(n_5593)
);

CKINVDCx16_ASAP7_75t_R g5594 ( 
.A(n_5492),
.Y(n_5594)
);

OR2x2_ASAP7_75t_L g5595 ( 
.A(n_5413),
.B(n_5340),
.Y(n_5595)
);

AND2x4_ASAP7_75t_L g5596 ( 
.A(n_5519),
.B(n_5315),
.Y(n_5596)
);

AND2x4_ASAP7_75t_L g5597 ( 
.A(n_5523),
.B(n_809),
.Y(n_5597)
);

INVx2_ASAP7_75t_L g5598 ( 
.A(n_5480),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5484),
.Y(n_5599)
);

NAND2xp5_ASAP7_75t_L g5600 ( 
.A(n_5445),
.B(n_810),
.Y(n_5600)
);

INVx3_ASAP7_75t_L g5601 ( 
.A(n_5526),
.Y(n_5601)
);

OR2x2_ASAP7_75t_L g5602 ( 
.A(n_5468),
.B(n_812),
.Y(n_5602)
);

INVx3_ASAP7_75t_L g5603 ( 
.A(n_5458),
.Y(n_5603)
);

INVx1_ASAP7_75t_SL g5604 ( 
.A(n_5463),
.Y(n_5604)
);

OR2x2_ASAP7_75t_L g5605 ( 
.A(n_5525),
.B(n_813),
.Y(n_5605)
);

INVxp33_ASAP7_75t_SL g5606 ( 
.A(n_5489),
.Y(n_5606)
);

NAND2xp5_ASAP7_75t_L g5607 ( 
.A(n_5451),
.B(n_814),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_5493),
.Y(n_5608)
);

INVx1_ASAP7_75t_SL g5609 ( 
.A(n_5491),
.Y(n_5609)
);

NAND3xp33_ASAP7_75t_L g5610 ( 
.A(n_5459),
.B(n_815),
.C(n_817),
.Y(n_5610)
);

NAND3xp33_ASAP7_75t_L g5611 ( 
.A(n_5470),
.B(n_815),
.C(n_817),
.Y(n_5611)
);

OAI21xp5_ASAP7_75t_L g5612 ( 
.A1(n_5443),
.A2(n_818),
.B(n_819),
.Y(n_5612)
);

AND2x2_ASAP7_75t_L g5613 ( 
.A(n_5472),
.B(n_818),
.Y(n_5613)
);

OR2x2_ASAP7_75t_L g5614 ( 
.A(n_5507),
.B(n_5538),
.Y(n_5614)
);

NOR2xp33_ASAP7_75t_L g5615 ( 
.A(n_5529),
.B(n_819),
.Y(n_5615)
);

AND2x2_ASAP7_75t_L g5616 ( 
.A(n_5483),
.B(n_820),
.Y(n_5616)
);

NAND2xp5_ASAP7_75t_L g5617 ( 
.A(n_5455),
.B(n_820),
.Y(n_5617)
);

NAND2x1p5_ASAP7_75t_L g5618 ( 
.A(n_5500),
.B(n_821),
.Y(n_5618)
);

OAI221xp5_ASAP7_75t_SL g5619 ( 
.A1(n_5446),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.C(n_824),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_5536),
.B(n_822),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5498),
.Y(n_5621)
);

AND2x2_ASAP7_75t_L g5622 ( 
.A(n_5511),
.B(n_825),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5514),
.B(n_826),
.Y(n_5623)
);

AND2x4_ASAP7_75t_L g5624 ( 
.A(n_5520),
.B(n_827),
.Y(n_5624)
);

AND2x4_ASAP7_75t_L g5625 ( 
.A(n_5537),
.B(n_828),
.Y(n_5625)
);

AND2x2_ASAP7_75t_L g5626 ( 
.A(n_5509),
.B(n_830),
.Y(n_5626)
);

NAND2xp5_ASAP7_75t_L g5627 ( 
.A(n_5530),
.B(n_831),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5516),
.Y(n_5628)
);

OR2x2_ASAP7_75t_L g5629 ( 
.A(n_5488),
.B(n_832),
.Y(n_5629)
);

AND2x2_ASAP7_75t_L g5630 ( 
.A(n_5442),
.B(n_5485),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5517),
.Y(n_5631)
);

OAI33xp33_ASAP7_75t_L g5632 ( 
.A1(n_5428),
.A2(n_834),
.A3(n_836),
.B1(n_832),
.B2(n_833),
.B3(n_835),
.Y(n_5632)
);

NOR2x1_ASAP7_75t_L g5633 ( 
.A(n_5534),
.B(n_834),
.Y(n_5633)
);

AND2x2_ASAP7_75t_L g5634 ( 
.A(n_5496),
.B(n_836),
.Y(n_5634)
);

AND2x2_ASAP7_75t_L g5635 ( 
.A(n_5543),
.B(n_5522),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5559),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_5609),
.B(n_5604),
.Y(n_5637)
);

AND2x2_ASAP7_75t_L g5638 ( 
.A(n_5551),
.B(n_5504),
.Y(n_5638)
);

OAI22xp5_ASAP7_75t_L g5639 ( 
.A1(n_5606),
.A2(n_5506),
.B1(n_5437),
.B2(n_5436),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5586),
.Y(n_5640)
);

NAND2xp5_ASAP7_75t_L g5641 ( 
.A(n_5554),
.B(n_5432),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_5630),
.B(n_5531),
.Y(n_5642)
);

AND2x2_ASAP7_75t_L g5643 ( 
.A(n_5558),
.B(n_5528),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5570),
.Y(n_5644)
);

INVx1_ASAP7_75t_SL g5645 ( 
.A(n_5591),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_L g5646 ( 
.A(n_5601),
.B(n_5603),
.Y(n_5646)
);

NAND2xp5_ASAP7_75t_L g5647 ( 
.A(n_5569),
.B(n_5555),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5623),
.Y(n_5648)
);

OR2x2_ASAP7_75t_L g5649 ( 
.A(n_5547),
.B(n_5449),
.Y(n_5649)
);

INVx1_ASAP7_75t_SL g5650 ( 
.A(n_5591),
.Y(n_5650)
);

OR2x2_ASAP7_75t_L g5651 ( 
.A(n_5546),
.B(n_5510),
.Y(n_5651)
);

INVx3_ASAP7_75t_L g5652 ( 
.A(n_5550),
.Y(n_5652)
);

AND2x2_ASAP7_75t_L g5653 ( 
.A(n_5561),
.B(n_5453),
.Y(n_5653)
);

OR2x2_ASAP7_75t_L g5654 ( 
.A(n_5556),
.B(n_5518),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_5590),
.Y(n_5655)
);

AOI21xp5_ASAP7_75t_SL g5656 ( 
.A1(n_5578),
.A2(n_5505),
.B(n_5535),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5616),
.Y(n_5657)
);

INVx2_ASAP7_75t_L g5658 ( 
.A(n_5618),
.Y(n_5658)
);

AND2x2_ASAP7_75t_L g5659 ( 
.A(n_5561),
.B(n_5497),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_5594),
.Y(n_5660)
);

NAND2xp5_ASAP7_75t_L g5661 ( 
.A(n_5581),
.B(n_5615),
.Y(n_5661)
);

AOI21xp5_ASAP7_75t_L g5662 ( 
.A1(n_5612),
.A2(n_5444),
.B(n_5439),
.Y(n_5662)
);

OR2x2_ASAP7_75t_L g5663 ( 
.A(n_5545),
.B(n_5533),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5629),
.Y(n_5664)
);

NAND3xp33_ASAP7_75t_L g5665 ( 
.A(n_5619),
.B(n_5633),
.C(n_5562),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5571),
.Y(n_5666)
);

OAI21xp5_ASAP7_75t_L g5667 ( 
.A1(n_5587),
.A2(n_5429),
.B(n_5541),
.Y(n_5667)
);

AOI22xp33_ASAP7_75t_L g5668 ( 
.A1(n_5598),
.A2(n_5540),
.B1(n_5542),
.B2(n_5482),
.Y(n_5668)
);

HB1xp67_ASAP7_75t_L g5669 ( 
.A(n_5596),
.Y(n_5669)
);

INVx2_ASAP7_75t_L g5670 ( 
.A(n_5585),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5595),
.Y(n_5671)
);

AND2x2_ASAP7_75t_L g5672 ( 
.A(n_5580),
.B(n_5425),
.Y(n_5672)
);

OAI21xp5_ASAP7_75t_L g5673 ( 
.A1(n_5610),
.A2(n_5467),
.B(n_5473),
.Y(n_5673)
);

HB1xp67_ASAP7_75t_L g5674 ( 
.A(n_5582),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5560),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5573),
.Y(n_5676)
);

OR2x2_ASAP7_75t_L g5677 ( 
.A(n_5614),
.B(n_5579),
.Y(n_5677)
);

OR2x2_ASAP7_75t_L g5678 ( 
.A(n_5553),
.B(n_5417),
.Y(n_5678)
);

NAND2xp5_ASAP7_75t_L g5679 ( 
.A(n_5626),
.B(n_5477),
.Y(n_5679)
);

OR2x2_ASAP7_75t_L g5680 ( 
.A(n_5584),
.B(n_5576),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5575),
.Y(n_5681)
);

INVxp67_ASAP7_75t_L g5682 ( 
.A(n_5597),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5583),
.Y(n_5683)
);

AND2x2_ASAP7_75t_L g5684 ( 
.A(n_5566),
.B(n_5513),
.Y(n_5684)
);

NAND4xp25_ASAP7_75t_L g5685 ( 
.A(n_5544),
.B(n_5478),
.C(n_5495),
.D(n_5475),
.Y(n_5685)
);

OR2x6_ASAP7_75t_L g5686 ( 
.A(n_5625),
.B(n_5605),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5588),
.Y(n_5687)
);

OR2x2_ASAP7_75t_L g5688 ( 
.A(n_5574),
.B(n_5499),
.Y(n_5688)
);

INVx2_ASAP7_75t_L g5689 ( 
.A(n_5568),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5593),
.Y(n_5690)
);

OR2x2_ASAP7_75t_L g5691 ( 
.A(n_5552),
.B(n_5508),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5599),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5608),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5621),
.Y(n_5694)
);

INVx1_ASAP7_75t_SL g5695 ( 
.A(n_5622),
.Y(n_5695)
);

AND2x2_ASAP7_75t_L g5696 ( 
.A(n_5577),
.B(n_838),
.Y(n_5696)
);

NAND2xp5_ASAP7_75t_L g5697 ( 
.A(n_5563),
.B(n_838),
.Y(n_5697)
);

AND2x2_ASAP7_75t_L g5698 ( 
.A(n_5549),
.B(n_839),
.Y(n_5698)
);

OR2x2_ASAP7_75t_L g5699 ( 
.A(n_5548),
.B(n_840),
.Y(n_5699)
);

INVxp67_ASAP7_75t_L g5700 ( 
.A(n_5589),
.Y(n_5700)
);

OR2x2_ASAP7_75t_L g5701 ( 
.A(n_5567),
.B(n_840),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5624),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5628),
.Y(n_5703)
);

OR2x2_ASAP7_75t_L g5704 ( 
.A(n_5565),
.B(n_841),
.Y(n_5704)
);

NAND3xp33_ASAP7_75t_L g5705 ( 
.A(n_5611),
.B(n_841),
.C(n_842),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_SL g5706 ( 
.A(n_5592),
.B(n_843),
.Y(n_5706)
);

NAND2x1p5_ASAP7_75t_L g5707 ( 
.A(n_5613),
.B(n_844),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5572),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5634),
.B(n_844),
.Y(n_5709)
);

NAND2xp33_ASAP7_75t_SL g5710 ( 
.A(n_5620),
.B(n_846),
.Y(n_5710)
);

OR2x2_ASAP7_75t_L g5711 ( 
.A(n_5602),
.B(n_846),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5631),
.Y(n_5712)
);

OR2x2_ASAP7_75t_L g5713 ( 
.A(n_5600),
.B(n_5607),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5617),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_5627),
.Y(n_5715)
);

AND2x4_ASAP7_75t_L g5716 ( 
.A(n_5557),
.B(n_848),
.Y(n_5716)
);

NAND3xp33_ASAP7_75t_L g5717 ( 
.A(n_5632),
.B(n_848),
.C(n_850),
.Y(n_5717)
);

INVxp67_ASAP7_75t_L g5718 ( 
.A(n_5564),
.Y(n_5718)
);

NAND2xp5_ASAP7_75t_L g5719 ( 
.A(n_5609),
.B(n_853),
.Y(n_5719)
);

INVxp67_ASAP7_75t_L g5720 ( 
.A(n_5674),
.Y(n_5720)
);

INVx2_ASAP7_75t_L g5721 ( 
.A(n_5707),
.Y(n_5721)
);

BUFx2_ASAP7_75t_L g5722 ( 
.A(n_5660),
.Y(n_5722)
);

OAI32xp33_ASAP7_75t_L g5723 ( 
.A1(n_5661),
.A2(n_856),
.A3(n_854),
.B1(n_855),
.B2(n_858),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5666),
.Y(n_5724)
);

INVx2_ASAP7_75t_L g5725 ( 
.A(n_5686),
.Y(n_5725)
);

AND2x2_ASAP7_75t_L g5726 ( 
.A(n_5638),
.B(n_860),
.Y(n_5726)
);

INVx2_ASAP7_75t_SL g5727 ( 
.A(n_5653),
.Y(n_5727)
);

AOI21xp33_ASAP7_75t_SL g5728 ( 
.A1(n_5718),
.A2(n_873),
.B(n_863),
.Y(n_5728)
);

NOR2xp33_ASAP7_75t_SL g5729 ( 
.A(n_5695),
.B(n_5682),
.Y(n_5729)
);

AOI32xp33_ASAP7_75t_L g5730 ( 
.A1(n_5716),
.A2(n_867),
.A3(n_864),
.B1(n_865),
.B2(n_868),
.Y(n_5730)
);

NAND2x1_ASAP7_75t_SL g5731 ( 
.A(n_5659),
.B(n_5643),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5711),
.Y(n_5732)
);

HB1xp67_ASAP7_75t_L g5733 ( 
.A(n_5645),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5719),
.Y(n_5734)
);

NOR2xp33_ASAP7_75t_L g5735 ( 
.A(n_5652),
.B(n_864),
.Y(n_5735)
);

NOR2xp33_ASAP7_75t_L g5736 ( 
.A(n_5642),
.B(n_867),
.Y(n_5736)
);

A2O1A1Ixp33_ASAP7_75t_L g5737 ( 
.A1(n_5662),
.A2(n_5665),
.B(n_5717),
.C(n_5673),
.Y(n_5737)
);

OR2x2_ASAP7_75t_L g5738 ( 
.A(n_5647),
.B(n_5637),
.Y(n_5738)
);

OAI21xp33_ASAP7_75t_SL g5739 ( 
.A1(n_5655),
.A2(n_868),
.B(n_869),
.Y(n_5739)
);

NOR3xp33_ASAP7_75t_L g5740 ( 
.A(n_5700),
.B(n_869),
.C(n_871),
.Y(n_5740)
);

NAND2x1p5_ASAP7_75t_L g5741 ( 
.A(n_5650),
.B(n_876),
.Y(n_5741)
);

O2A1O1Ixp5_ASAP7_75t_L g5742 ( 
.A1(n_5706),
.A2(n_878),
.B(n_875),
.C(n_877),
.Y(n_5742)
);

NOR2xp33_ASAP7_75t_L g5743 ( 
.A(n_5713),
.B(n_877),
.Y(n_5743)
);

OAI22xp5_ASAP7_75t_L g5744 ( 
.A1(n_5654),
.A2(n_880),
.B1(n_878),
.B2(n_879),
.Y(n_5744)
);

AOI221xp5_ASAP7_75t_L g5745 ( 
.A1(n_5715),
.A2(n_884),
.B1(n_882),
.B2(n_883),
.C(n_885),
.Y(n_5745)
);

AOI22xp5_ASAP7_75t_L g5746 ( 
.A1(n_5710),
.A2(n_5668),
.B1(n_5679),
.B2(n_5705),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5636),
.Y(n_5747)
);

OAI21xp33_ASAP7_75t_L g5748 ( 
.A1(n_5635),
.A2(n_885),
.B(n_886),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5688),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5640),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_5664),
.Y(n_5751)
);

INVx2_ASAP7_75t_L g5752 ( 
.A(n_5696),
.Y(n_5752)
);

NAND3xp33_ASAP7_75t_L g5753 ( 
.A(n_5639),
.B(n_886),
.C(n_887),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5709),
.Y(n_5754)
);

AOI22xp33_ASAP7_75t_SL g5755 ( 
.A1(n_5641),
.A2(n_889),
.B1(n_887),
.B2(n_888),
.Y(n_5755)
);

AND2x4_ASAP7_75t_L g5756 ( 
.A(n_5670),
.B(n_5684),
.Y(n_5756)
);

OAI21xp33_ASAP7_75t_SL g5757 ( 
.A1(n_5644),
.A2(n_5671),
.B(n_5649),
.Y(n_5757)
);

NOR2xp33_ASAP7_75t_L g5758 ( 
.A(n_5701),
.B(n_890),
.Y(n_5758)
);

INVx3_ASAP7_75t_L g5759 ( 
.A(n_5689),
.Y(n_5759)
);

INVx2_ASAP7_75t_L g5760 ( 
.A(n_5702),
.Y(n_5760)
);

NAND2xp5_ASAP7_75t_L g5761 ( 
.A(n_5657),
.B(n_891),
.Y(n_5761)
);

OAI22xp5_ASAP7_75t_L g5762 ( 
.A1(n_5651),
.A2(n_893),
.B1(n_891),
.B2(n_892),
.Y(n_5762)
);

NOR2xp33_ASAP7_75t_L g5763 ( 
.A(n_5697),
.B(n_892),
.Y(n_5763)
);

NOR2xp33_ASAP7_75t_L g5764 ( 
.A(n_5704),
.B(n_893),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5714),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5691),
.Y(n_5766)
);

NAND3xp33_ASAP7_75t_L g5767 ( 
.A(n_5656),
.B(n_894),
.C(n_895),
.Y(n_5767)
);

NOR2xp67_ASAP7_75t_L g5768 ( 
.A(n_5685),
.B(n_894),
.Y(n_5768)
);

NAND2xp5_ASAP7_75t_L g5769 ( 
.A(n_5698),
.B(n_895),
.Y(n_5769)
);

AOI22xp33_ASAP7_75t_L g5770 ( 
.A1(n_5680),
.A2(n_898),
.B1(n_896),
.B2(n_897),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5699),
.Y(n_5771)
);

OAI21xp33_ASAP7_75t_L g5772 ( 
.A1(n_5646),
.A2(n_899),
.B(n_900),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_5658),
.Y(n_5773)
);

OR2x2_ASAP7_75t_L g5774 ( 
.A(n_5663),
.B(n_901),
.Y(n_5774)
);

AOI21xp33_ASAP7_75t_L g5775 ( 
.A1(n_5678),
.A2(n_903),
.B(n_904),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5648),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5675),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5676),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5672),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5681),
.Y(n_5780)
);

OAI21xp5_ASAP7_75t_L g5781 ( 
.A1(n_5712),
.A2(n_906),
.B(n_905),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5683),
.Y(n_5782)
);

INVx3_ASAP7_75t_L g5783 ( 
.A(n_5708),
.Y(n_5783)
);

AOI211xp5_ASAP7_75t_L g5784 ( 
.A1(n_5687),
.A2(n_909),
.B(n_907),
.C(n_908),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5690),
.Y(n_5785)
);

AND2x2_ASAP7_75t_L g5786 ( 
.A(n_5692),
.B(n_912),
.Y(n_5786)
);

INVx2_ASAP7_75t_L g5787 ( 
.A(n_5693),
.Y(n_5787)
);

OA21x2_ASAP7_75t_L g5788 ( 
.A1(n_5694),
.A2(n_912),
.B(n_913),
.Y(n_5788)
);

AND2x2_ASAP7_75t_L g5789 ( 
.A(n_5703),
.B(n_916),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5677),
.Y(n_5790)
);

AOI221xp5_ASAP7_75t_L g5791 ( 
.A1(n_5716),
.A2(n_921),
.B1(n_918),
.B2(n_920),
.C(n_922),
.Y(n_5791)
);

INVx1_ASAP7_75t_SL g5792 ( 
.A(n_5669),
.Y(n_5792)
);

OAI211xp5_ASAP7_75t_SL g5793 ( 
.A1(n_5680),
.A2(n_925),
.B(n_922),
.C(n_924),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_5677),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5677),
.Y(n_5795)
);

O2A1O1Ixp33_ASAP7_75t_L g5796 ( 
.A1(n_5667),
.A2(n_927),
.B(n_924),
.C(n_926),
.Y(n_5796)
);

NOR2xp33_ASAP7_75t_SL g5797 ( 
.A(n_5733),
.B(n_5792),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5788),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5788),
.Y(n_5799)
);

NAND2xp5_ASAP7_75t_L g5800 ( 
.A(n_5726),
.B(n_929),
.Y(n_5800)
);

AND2x2_ASAP7_75t_L g5801 ( 
.A(n_5722),
.B(n_930),
.Y(n_5801)
);

OAI22xp5_ASAP7_75t_L g5802 ( 
.A1(n_5767),
.A2(n_933),
.B1(n_931),
.B2(n_932),
.Y(n_5802)
);

AOI21xp5_ASAP7_75t_L g5803 ( 
.A1(n_5737),
.A2(n_932),
.B(n_933),
.Y(n_5803)
);

OAI21xp5_ASAP7_75t_L g5804 ( 
.A1(n_5731),
.A2(n_934),
.B(n_935),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_5790),
.Y(n_5805)
);

NOR2xp33_ASAP7_75t_L g5806 ( 
.A(n_5728),
.B(n_936),
.Y(n_5806)
);

OAI21xp33_ASAP7_75t_L g5807 ( 
.A1(n_5729),
.A2(n_937),
.B(n_939),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5794),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5795),
.Y(n_5809)
);

AOI211xp5_ASAP7_75t_L g5810 ( 
.A1(n_5753),
.A2(n_945),
.B(n_943),
.C(n_944),
.Y(n_5810)
);

NAND3xp33_ASAP7_75t_L g5811 ( 
.A(n_5720),
.B(n_943),
.C(n_944),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5774),
.Y(n_5812)
);

OAI22xp5_ASAP7_75t_L g5813 ( 
.A1(n_5727),
.A2(n_5738),
.B1(n_5756),
.B2(n_5755),
.Y(n_5813)
);

OR2x2_ASAP7_75t_L g5814 ( 
.A(n_5766),
.B(n_5749),
.Y(n_5814)
);

NAND2xp5_ASAP7_75t_L g5815 ( 
.A(n_5752),
.B(n_946),
.Y(n_5815)
);

NAND2xp5_ASAP7_75t_L g5816 ( 
.A(n_5743),
.B(n_947),
.Y(n_5816)
);

OAI22xp33_ASAP7_75t_L g5817 ( 
.A1(n_5779),
.A2(n_951),
.B1(n_949),
.B2(n_950),
.Y(n_5817)
);

NAND2xp5_ASAP7_75t_L g5818 ( 
.A(n_5736),
.B(n_950),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_5786),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_5732),
.B(n_952),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5789),
.Y(n_5821)
);

OAI221xp5_ASAP7_75t_L g5822 ( 
.A1(n_5742),
.A2(n_955),
.B1(n_953),
.B2(n_954),
.C(n_956),
.Y(n_5822)
);

NAND2x1_ASAP7_75t_L g5823 ( 
.A(n_5783),
.B(n_956),
.Y(n_5823)
);

AOI22xp5_ASAP7_75t_L g5824 ( 
.A1(n_5734),
.A2(n_959),
.B1(n_957),
.B2(n_958),
.Y(n_5824)
);

OAI22xp5_ASAP7_75t_L g5825 ( 
.A1(n_5770),
.A2(n_962),
.B1(n_959),
.B2(n_960),
.Y(n_5825)
);

OAI33xp33_ASAP7_75t_L g5826 ( 
.A1(n_5747),
.A2(n_967),
.A3(n_970),
.B1(n_963),
.B2(n_966),
.B3(n_969),
.Y(n_5826)
);

AND2x2_ASAP7_75t_L g5827 ( 
.A(n_5735),
.B(n_5751),
.Y(n_5827)
);

AOI221xp5_ASAP7_75t_L g5828 ( 
.A1(n_5723),
.A2(n_974),
.B1(n_976),
.B2(n_973),
.C(n_975),
.Y(n_5828)
);

NAND2xp5_ASAP7_75t_L g5829 ( 
.A(n_5764),
.B(n_972),
.Y(n_5829)
);

AOI22x1_ASAP7_75t_L g5830 ( 
.A1(n_5750),
.A2(n_981),
.B1(n_979),
.B2(n_980),
.Y(n_5830)
);

AOI221xp5_ASAP7_75t_SL g5831 ( 
.A1(n_5724),
.A2(n_5777),
.B1(n_5765),
.B2(n_5776),
.C(n_5778),
.Y(n_5831)
);

OAI21xp5_ASAP7_75t_L g5832 ( 
.A1(n_5796),
.A2(n_5740),
.B(n_5744),
.Y(n_5832)
);

OAI321xp33_ASAP7_75t_L g5833 ( 
.A1(n_5725),
.A2(n_985),
.A3(n_987),
.B1(n_988),
.B2(n_984),
.C(n_986),
.Y(n_5833)
);

NAND2xp5_ASAP7_75t_L g5834 ( 
.A(n_5758),
.B(n_986),
.Y(n_5834)
);

OA21x2_ASAP7_75t_L g5835 ( 
.A1(n_5775),
.A2(n_987),
.B(n_988),
.Y(n_5835)
);

NAND2xp5_ASAP7_75t_L g5836 ( 
.A(n_5763),
.B(n_989),
.Y(n_5836)
);

AOI22xp5_ASAP7_75t_L g5837 ( 
.A1(n_5721),
.A2(n_991),
.B1(n_989),
.B2(n_990),
.Y(n_5837)
);

AOI22xp5_ASAP7_75t_L g5838 ( 
.A1(n_5773),
.A2(n_5754),
.B1(n_5771),
.B2(n_5748),
.Y(n_5838)
);

OR2x2_ASAP7_75t_L g5839 ( 
.A(n_5761),
.B(n_5787),
.Y(n_5839)
);

OAI32xp33_ASAP7_75t_L g5840 ( 
.A1(n_5793),
.A2(n_994),
.A3(n_992),
.B1(n_993),
.B2(n_997),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5760),
.Y(n_5841)
);

O2A1O1Ixp33_ASAP7_75t_SL g5842 ( 
.A1(n_5780),
.A2(n_994),
.B(n_992),
.C(n_993),
.Y(n_5842)
);

AND2x2_ASAP7_75t_L g5843 ( 
.A(n_5781),
.B(n_997),
.Y(n_5843)
);

AOI22xp5_ASAP7_75t_L g5844 ( 
.A1(n_5759),
.A2(n_1000),
.B1(n_998),
.B2(n_999),
.Y(n_5844)
);

OR2x2_ASAP7_75t_L g5845 ( 
.A(n_5782),
.B(n_5785),
.Y(n_5845)
);

NAND2xp5_ASAP7_75t_L g5846 ( 
.A(n_5730),
.B(n_1001),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5769),
.Y(n_5847)
);

AND2x2_ASAP7_75t_L g5848 ( 
.A(n_5772),
.B(n_1003),
.Y(n_5848)
);

AOI21xp5_ASAP7_75t_L g5849 ( 
.A1(n_5762),
.A2(n_1003),
.B(n_1004),
.Y(n_5849)
);

NAND2xp5_ASAP7_75t_L g5850 ( 
.A(n_5784),
.B(n_1004),
.Y(n_5850)
);

NAND2xp5_ASAP7_75t_L g5851 ( 
.A(n_5791),
.B(n_1005),
.Y(n_5851)
);

NAND2xp5_ASAP7_75t_L g5852 ( 
.A(n_5745),
.B(n_1005),
.Y(n_5852)
);

AND2x2_ASAP7_75t_L g5853 ( 
.A(n_5733),
.B(n_1006),
.Y(n_5853)
);

OA21x2_ASAP7_75t_L g5854 ( 
.A1(n_5767),
.A2(n_1008),
.B(n_1009),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5733),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5733),
.Y(n_5856)
);

NAND2xp5_ASAP7_75t_L g5857 ( 
.A(n_5726),
.B(n_1012),
.Y(n_5857)
);

INVx1_ASAP7_75t_L g5858 ( 
.A(n_5733),
.Y(n_5858)
);

NAND2xp5_ASAP7_75t_L g5859 ( 
.A(n_5726),
.B(n_1013),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5733),
.Y(n_5860)
);

AOI222xp33_ASAP7_75t_L g5861 ( 
.A1(n_5757),
.A2(n_1017),
.B1(n_1020),
.B2(n_1014),
.C1(n_1016),
.C2(n_1019),
.Y(n_5861)
);

OAI22xp5_ASAP7_75t_L g5862 ( 
.A1(n_5792),
.A2(n_1022),
.B1(n_1016),
.B2(n_1021),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5733),
.Y(n_5863)
);

A2O1A1Ixp33_ASAP7_75t_L g5864 ( 
.A1(n_5739),
.A2(n_1710),
.B(n_1023),
.C(n_1021),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5733),
.Y(n_5865)
);

OAI21xp5_ASAP7_75t_L g5866 ( 
.A1(n_5757),
.A2(n_1024),
.B(n_1025),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5733),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5733),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5733),
.Y(n_5869)
);

AOI21xp33_ASAP7_75t_SL g5870 ( 
.A1(n_5733),
.A2(n_1028),
.B(n_1029),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_L g5871 ( 
.A(n_5726),
.B(n_1036),
.Y(n_5871)
);

OR2x2_ASAP7_75t_L g5872 ( 
.A(n_5792),
.B(n_1036),
.Y(n_5872)
);

AOI22xp33_ASAP7_75t_L g5873 ( 
.A1(n_5768),
.A2(n_1039),
.B1(n_1037),
.B2(n_1038),
.Y(n_5873)
);

INVxp67_ASAP7_75t_L g5874 ( 
.A(n_5729),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5733),
.Y(n_5875)
);

NOR3xp33_ASAP7_75t_L g5876 ( 
.A(n_5757),
.B(n_1037),
.C(n_1039),
.Y(n_5876)
);

NOR2xp33_ASAP7_75t_L g5877 ( 
.A(n_5741),
.B(n_1040),
.Y(n_5877)
);

A2O1A1Ixp33_ASAP7_75t_L g5878 ( 
.A1(n_5739),
.A2(n_1696),
.B(n_1697),
.C(n_1695),
.Y(n_5878)
);

AOI222xp33_ASAP7_75t_L g5879 ( 
.A1(n_5757),
.A2(n_1045),
.B1(n_1047),
.B2(n_1043),
.C1(n_1044),
.C2(n_1046),
.Y(n_5879)
);

AOI22xp5_ASAP7_75t_L g5880 ( 
.A1(n_5746),
.A2(n_1049),
.B1(n_1047),
.B2(n_1048),
.Y(n_5880)
);

OAI21xp5_ASAP7_75t_SL g5881 ( 
.A1(n_5792),
.A2(n_1050),
.B(n_1051),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_L g5882 ( 
.A(n_5726),
.B(n_1054),
.Y(n_5882)
);

AOI21xp5_ASAP7_75t_L g5883 ( 
.A1(n_5757),
.A2(n_1055),
.B(n_1057),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_5726),
.B(n_1058),
.Y(n_5884)
);

NAND2x1_ASAP7_75t_SL g5885 ( 
.A(n_5733),
.B(n_1059),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5733),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5733),
.Y(n_5887)
);

OA21x2_ASAP7_75t_L g5888 ( 
.A1(n_5767),
.A2(n_1061),
.B(n_1062),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_5733),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5733),
.Y(n_5890)
);

NAND2xp33_ASAP7_75t_SL g5891 ( 
.A(n_5731),
.B(n_1062),
.Y(n_5891)
);

INVx1_ASAP7_75t_SL g5892 ( 
.A(n_5731),
.Y(n_5892)
);

AOI322xp5_ASAP7_75t_L g5893 ( 
.A1(n_5746),
.A2(n_1070),
.A3(n_1069),
.B1(n_1066),
.B2(n_1064),
.C1(n_1065),
.C2(n_1067),
.Y(n_5893)
);

OAI21xp5_ASAP7_75t_L g5894 ( 
.A1(n_5883),
.A2(n_1064),
.B(n_1065),
.Y(n_5894)
);

OAI32xp33_ASAP7_75t_L g5895 ( 
.A1(n_5876),
.A2(n_1070),
.A3(n_1066),
.B1(n_1069),
.B2(n_1071),
.Y(n_5895)
);

AOI21xp33_ASAP7_75t_L g5896 ( 
.A1(n_5892),
.A2(n_5799),
.B(n_5798),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5801),
.Y(n_5897)
);

NOR2xp33_ASAP7_75t_L g5898 ( 
.A(n_5874),
.B(n_1071),
.Y(n_5898)
);

INVxp67_ASAP7_75t_SL g5899 ( 
.A(n_5885),
.Y(n_5899)
);

INVx1_ASAP7_75t_SL g5900 ( 
.A(n_5891),
.Y(n_5900)
);

INVxp67_ASAP7_75t_L g5901 ( 
.A(n_5797),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5853),
.Y(n_5902)
);

NAND2xp5_ASAP7_75t_L g5903 ( 
.A(n_5864),
.B(n_1079),
.Y(n_5903)
);

A2O1A1Ixp33_ASAP7_75t_L g5904 ( 
.A1(n_5803),
.A2(n_1083),
.B(n_1080),
.C(n_1082),
.Y(n_5904)
);

OAI21xp5_ASAP7_75t_L g5905 ( 
.A1(n_5866),
.A2(n_5804),
.B(n_5861),
.Y(n_5905)
);

CKINVDCx14_ASAP7_75t_R g5906 ( 
.A(n_5813),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5855),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5856),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5858),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5860),
.Y(n_5910)
);

NAND2x1_ASAP7_75t_L g5911 ( 
.A(n_5863),
.B(n_1084),
.Y(n_5911)
);

AOI21xp5_ASAP7_75t_L g5912 ( 
.A1(n_5842),
.A2(n_1086),
.B(n_1087),
.Y(n_5912)
);

O2A1O1Ixp33_ASAP7_75t_L g5913 ( 
.A1(n_5879),
.A2(n_1089),
.B(n_1087),
.C(n_1088),
.Y(n_5913)
);

OAI31xp33_ASAP7_75t_L g5914 ( 
.A1(n_5878),
.A2(n_1093),
.A3(n_1090),
.B(n_1092),
.Y(n_5914)
);

NAND2xp5_ASAP7_75t_L g5915 ( 
.A(n_5870),
.B(n_5881),
.Y(n_5915)
);

HB1xp67_ASAP7_75t_L g5916 ( 
.A(n_5823),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5865),
.Y(n_5917)
);

NAND2x1_ASAP7_75t_L g5918 ( 
.A(n_5867),
.B(n_1094),
.Y(n_5918)
);

AND2x4_ASAP7_75t_L g5919 ( 
.A(n_5868),
.B(n_1094),
.Y(n_5919)
);

NOR3xp33_ASAP7_75t_L g5920 ( 
.A(n_5841),
.B(n_1706),
.C(n_1096),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_5869),
.Y(n_5921)
);

AND2x4_ASAP7_75t_L g5922 ( 
.A(n_5875),
.B(n_1097),
.Y(n_5922)
);

AOI22xp5_ASAP7_75t_L g5923 ( 
.A1(n_5812),
.A2(n_1100),
.B1(n_1098),
.B2(n_1099),
.Y(n_5923)
);

INVxp67_ASAP7_75t_SL g5924 ( 
.A(n_5877),
.Y(n_5924)
);

INVx2_ASAP7_75t_L g5925 ( 
.A(n_5830),
.Y(n_5925)
);

XNOR2xp5_ASAP7_75t_L g5926 ( 
.A(n_5838),
.B(n_1104),
.Y(n_5926)
);

AOI221xp5_ASAP7_75t_L g5927 ( 
.A1(n_5832),
.A2(n_1107),
.B1(n_1105),
.B2(n_1106),
.C(n_1108),
.Y(n_5927)
);

NOR2xp33_ASAP7_75t_L g5928 ( 
.A(n_5826),
.B(n_1111),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5886),
.Y(n_5929)
);

NAND2xp33_ASAP7_75t_L g5930 ( 
.A(n_5887),
.B(n_5889),
.Y(n_5930)
);

INVx1_ASAP7_75t_SL g5931 ( 
.A(n_5872),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5819),
.B(n_1113),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5890),
.Y(n_5933)
);

NAND2xp5_ASAP7_75t_L g5934 ( 
.A(n_5821),
.B(n_1119),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5800),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5857),
.Y(n_5936)
);

INVx1_ASAP7_75t_SL g5937 ( 
.A(n_5814),
.Y(n_5937)
);

INVxp67_ASAP7_75t_L g5938 ( 
.A(n_5806),
.Y(n_5938)
);

INVx1_ASAP7_75t_L g5939 ( 
.A(n_5859),
.Y(n_5939)
);

OAI32xp33_ASAP7_75t_L g5940 ( 
.A1(n_5845),
.A2(n_1125),
.A3(n_1123),
.B1(n_1124),
.B2(n_1126),
.Y(n_5940)
);

CKINVDCx5p33_ASAP7_75t_R g5941 ( 
.A(n_5871),
.Y(n_5941)
);

INVxp67_ASAP7_75t_L g5942 ( 
.A(n_5882),
.Y(n_5942)
);

AND2x2_ASAP7_75t_L g5943 ( 
.A(n_5827),
.B(n_5805),
.Y(n_5943)
);

INVx3_ASAP7_75t_L g5944 ( 
.A(n_5839),
.Y(n_5944)
);

AND2x2_ASAP7_75t_L g5945 ( 
.A(n_5808),
.B(n_1127),
.Y(n_5945)
);

NAND2xp5_ASAP7_75t_L g5946 ( 
.A(n_5893),
.B(n_1129),
.Y(n_5946)
);

NOR2xp33_ASAP7_75t_L g5947 ( 
.A(n_5807),
.B(n_1130),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5884),
.Y(n_5948)
);

AOI222xp33_ASAP7_75t_L g5949 ( 
.A1(n_5809),
.A2(n_5847),
.B1(n_5873),
.B2(n_5822),
.C1(n_5828),
.C2(n_5802),
.Y(n_5949)
);

AND2x2_ASAP7_75t_L g5950 ( 
.A(n_5831),
.B(n_1130),
.Y(n_5950)
);

INVxp67_ASAP7_75t_L g5951 ( 
.A(n_5854),
.Y(n_5951)
);

NAND2xp5_ASAP7_75t_L g5952 ( 
.A(n_5843),
.B(n_1135),
.Y(n_5952)
);

OA21x2_ASAP7_75t_L g5953 ( 
.A1(n_5820),
.A2(n_1136),
.B(n_1137),
.Y(n_5953)
);

OAI221xp5_ASAP7_75t_L g5954 ( 
.A1(n_5854),
.A2(n_1140),
.B1(n_1138),
.B2(n_1139),
.C(n_1141),
.Y(n_5954)
);

INVx1_ASAP7_75t_L g5955 ( 
.A(n_5836),
.Y(n_5955)
);

NAND2xp5_ASAP7_75t_L g5956 ( 
.A(n_5810),
.B(n_1138),
.Y(n_5956)
);

AOI222xp33_ASAP7_75t_L g5957 ( 
.A1(n_5840),
.A2(n_5833),
.B1(n_5852),
.B2(n_5850),
.C1(n_5851),
.C2(n_5825),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5829),
.Y(n_5958)
);

AOI21xp33_ASAP7_75t_SL g5959 ( 
.A1(n_5888),
.A2(n_1144),
.B(n_1143),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5834),
.Y(n_5960)
);

OR2x2_ASAP7_75t_L g5961 ( 
.A(n_5815),
.B(n_1145),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5816),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5818),
.Y(n_5963)
);

INVx2_ASAP7_75t_L g5964 ( 
.A(n_5835),
.Y(n_5964)
);

HB1xp67_ASAP7_75t_L g5965 ( 
.A(n_5848),
.Y(n_5965)
);

NAND2xp5_ASAP7_75t_L g5966 ( 
.A(n_5899),
.B(n_5849),
.Y(n_5966)
);

NAND2xp5_ASAP7_75t_SL g5967 ( 
.A(n_5901),
.B(n_5880),
.Y(n_5967)
);

AOI22xp33_ASAP7_75t_L g5968 ( 
.A1(n_5964),
.A2(n_5811),
.B1(n_5846),
.B2(n_5862),
.Y(n_5968)
);

O2A1O1Ixp33_ASAP7_75t_L g5969 ( 
.A1(n_5951),
.A2(n_5817),
.B(n_5824),
.C(n_5844),
.Y(n_5969)
);

OAI21xp33_ASAP7_75t_L g5970 ( 
.A1(n_5906),
.A2(n_5837),
.B(n_1147),
.Y(n_5970)
);

NAND3xp33_ASAP7_75t_SL g5971 ( 
.A(n_5937),
.B(n_1148),
.C(n_1149),
.Y(n_5971)
);

XNOR2xp5_ASAP7_75t_L g5972 ( 
.A(n_5926),
.B(n_5941),
.Y(n_5972)
);

NAND2xp33_ASAP7_75t_L g5973 ( 
.A(n_5916),
.B(n_1149),
.Y(n_5973)
);

NOR3xp33_ASAP7_75t_L g5974 ( 
.A(n_5944),
.B(n_1150),
.C(n_1151),
.Y(n_5974)
);

AOI33xp33_ASAP7_75t_L g5975 ( 
.A1(n_5907),
.A2(n_1154),
.A3(n_1156),
.B1(n_1152),
.B2(n_1153),
.B3(n_1155),
.Y(n_5975)
);

AOI21xp5_ASAP7_75t_L g5976 ( 
.A1(n_5930),
.A2(n_1156),
.B(n_1153),
.Y(n_5976)
);

INVx1_ASAP7_75t_SL g5977 ( 
.A(n_5943),
.Y(n_5977)
);

AOI221xp5_ASAP7_75t_L g5978 ( 
.A1(n_5905),
.A2(n_1170),
.B1(n_1179),
.B2(n_1162),
.C(n_1157),
.Y(n_5978)
);

NAND4xp25_ASAP7_75t_L g5979 ( 
.A(n_5949),
.B(n_1702),
.C(n_1162),
.D(n_1160),
.Y(n_5979)
);

AOI21xp5_ASAP7_75t_L g5980 ( 
.A1(n_5911),
.A2(n_1163),
.B(n_1161),
.Y(n_5980)
);

AOI211xp5_ASAP7_75t_SL g5981 ( 
.A1(n_5950),
.A2(n_5909),
.B(n_5910),
.C(n_5908),
.Y(n_5981)
);

NAND3xp33_ASAP7_75t_L g5982 ( 
.A(n_5959),
.B(n_1160),
.C(n_1161),
.Y(n_5982)
);

OAI22xp5_ASAP7_75t_L g5983 ( 
.A1(n_5925),
.A2(n_1166),
.B1(n_1164),
.B2(n_1165),
.Y(n_5983)
);

OAI221xp5_ASAP7_75t_SL g5984 ( 
.A1(n_5931),
.A2(n_1693),
.B1(n_1694),
.B2(n_1691),
.C(n_1690),
.Y(n_5984)
);

OA211x2_ASAP7_75t_L g5985 ( 
.A1(n_5918),
.A2(n_1168),
.B(n_1166),
.C(n_1167),
.Y(n_5985)
);

HB1xp67_ASAP7_75t_L g5986 ( 
.A(n_5915),
.Y(n_5986)
);

AOI211xp5_ASAP7_75t_L g5987 ( 
.A1(n_5917),
.A2(n_1696),
.B(n_1697),
.C(n_1695),
.Y(n_5987)
);

AOI222xp33_ASAP7_75t_L g5988 ( 
.A1(n_5938),
.A2(n_1173),
.B1(n_1176),
.B2(n_1171),
.C1(n_1172),
.C2(n_1175),
.Y(n_5988)
);

OAI21xp5_ASAP7_75t_L g5989 ( 
.A1(n_5912),
.A2(n_1172),
.B(n_1173),
.Y(n_5989)
);

AOI221xp5_ASAP7_75t_SL g5990 ( 
.A1(n_5921),
.A2(n_1177),
.B1(n_1175),
.B2(n_1176),
.C(n_1179),
.Y(n_5990)
);

OAI221xp5_ASAP7_75t_L g5991 ( 
.A1(n_5897),
.A2(n_1183),
.B1(n_1177),
.B2(n_1182),
.C(n_1184),
.Y(n_5991)
);

NOR2xp33_ASAP7_75t_SL g5992 ( 
.A(n_5902),
.B(n_1186),
.Y(n_5992)
);

O2A1O1Ixp33_ASAP7_75t_L g5993 ( 
.A1(n_5954),
.A2(n_1190),
.B(n_1187),
.C(n_1189),
.Y(n_5993)
);

AOI21xp5_ASAP7_75t_L g5994 ( 
.A1(n_5946),
.A2(n_1193),
.B(n_1192),
.Y(n_5994)
);

AOI22xp33_ASAP7_75t_L g5995 ( 
.A1(n_5965),
.A2(n_1197),
.B1(n_1194),
.B2(n_1195),
.Y(n_5995)
);

OAI21xp33_ASAP7_75t_SL g5996 ( 
.A1(n_5929),
.A2(n_1198),
.B(n_1199),
.Y(n_5996)
);

AOI221x1_ASAP7_75t_L g5997 ( 
.A1(n_5933),
.A2(n_1202),
.B1(n_1200),
.B2(n_1201),
.C(n_1203),
.Y(n_5997)
);

NAND3xp33_ASAP7_75t_SL g5998 ( 
.A(n_5957),
.B(n_1200),
.C(n_1203),
.Y(n_5998)
);

OAI211xp5_ASAP7_75t_L g5999 ( 
.A1(n_5924),
.A2(n_1210),
.B(n_1207),
.C(n_1208),
.Y(n_5999)
);

AOI21xp33_ASAP7_75t_L g6000 ( 
.A1(n_5942),
.A2(n_1208),
.B(n_1211),
.Y(n_6000)
);

AOI22xp5_ASAP7_75t_L g6001 ( 
.A1(n_5928),
.A2(n_1221),
.B1(n_1228),
.B2(n_1213),
.Y(n_6001)
);

INVx1_ASAP7_75t_L g6002 ( 
.A(n_5953),
.Y(n_6002)
);

AOI22xp33_ASAP7_75t_SL g6003 ( 
.A1(n_5955),
.A2(n_5963),
.B1(n_5960),
.B2(n_5962),
.Y(n_6003)
);

AOI211xp5_ASAP7_75t_L g6004 ( 
.A1(n_5898),
.A2(n_1218),
.B(n_1214),
.C(n_1217),
.Y(n_6004)
);

OAI31xp33_ASAP7_75t_L g6005 ( 
.A1(n_5904),
.A2(n_1221),
.A3(n_1219),
.B(n_1220),
.Y(n_6005)
);

NAND2xp5_ASAP7_75t_L g6006 ( 
.A(n_5919),
.B(n_1220),
.Y(n_6006)
);

AOI322xp5_ASAP7_75t_L g6007 ( 
.A1(n_5958),
.A2(n_1227),
.A3(n_1226),
.B1(n_1224),
.B2(n_1222),
.C1(n_1223),
.C2(n_1225),
.Y(n_6007)
);

NAND4xp25_ASAP7_75t_L g6008 ( 
.A(n_5935),
.B(n_5939),
.C(n_5948),
.D(n_5936),
.Y(n_6008)
);

NOR2xp33_ASAP7_75t_L g6009 ( 
.A(n_5895),
.B(n_1229),
.Y(n_6009)
);

OAI221xp5_ASAP7_75t_L g6010 ( 
.A1(n_5894),
.A2(n_1232),
.B1(n_1230),
.B2(n_1231),
.C(n_1233),
.Y(n_6010)
);

AOI221xp5_ASAP7_75t_L g6011 ( 
.A1(n_5913),
.A2(n_1248),
.B1(n_1254),
.B2(n_1240),
.C(n_1234),
.Y(n_6011)
);

NAND2xp5_ASAP7_75t_L g6012 ( 
.A(n_5922),
.B(n_1237),
.Y(n_6012)
);

AOI211xp5_ASAP7_75t_SL g6013 ( 
.A1(n_5932),
.A2(n_1239),
.B(n_1237),
.C(n_1238),
.Y(n_6013)
);

OAI21xp5_ASAP7_75t_SL g6014 ( 
.A1(n_5934),
.A2(n_1238),
.B(n_1239),
.Y(n_6014)
);

AOI32xp33_ASAP7_75t_L g6015 ( 
.A1(n_5947),
.A2(n_1244),
.A3(n_1242),
.B1(n_1243),
.B2(n_1245),
.Y(n_6015)
);

AOI222xp33_ASAP7_75t_L g6016 ( 
.A1(n_5903),
.A2(n_1245),
.B1(n_1247),
.B2(n_1242),
.C1(n_1243),
.C2(n_1246),
.Y(n_6016)
);

NAND2xp5_ASAP7_75t_L g6017 ( 
.A(n_5945),
.B(n_1246),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5961),
.Y(n_6018)
);

AND4x1_ASAP7_75t_L g6019 ( 
.A(n_5927),
.B(n_1250),
.C(n_1251),
.D(n_1249),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5952),
.Y(n_6020)
);

AOI222xp33_ASAP7_75t_L g6021 ( 
.A1(n_5956),
.A2(n_1251),
.B1(n_1253),
.B2(n_1248),
.C1(n_1249),
.C2(n_1252),
.Y(n_6021)
);

AOI211xp5_ASAP7_75t_L g6022 ( 
.A1(n_5940),
.A2(n_1690),
.B(n_1694),
.C(n_1689),
.Y(n_6022)
);

NAND2xp5_ASAP7_75t_L g6023 ( 
.A(n_5920),
.B(n_5914),
.Y(n_6023)
);

OAI21xp5_ASAP7_75t_SL g6024 ( 
.A1(n_5923),
.A2(n_1255),
.B(n_1257),
.Y(n_6024)
);

INVxp67_ASAP7_75t_SL g6025 ( 
.A(n_5901),
.Y(n_6025)
);

O2A1O1Ixp33_ASAP7_75t_L g6026 ( 
.A1(n_5951),
.A2(n_1263),
.B(n_1261),
.C(n_1262),
.Y(n_6026)
);

NAND2xp5_ASAP7_75t_SL g6027 ( 
.A(n_5901),
.B(n_1264),
.Y(n_6027)
);

NAND2xp5_ASAP7_75t_L g6028 ( 
.A(n_5899),
.B(n_1265),
.Y(n_6028)
);

NAND3xp33_ASAP7_75t_SL g6029 ( 
.A(n_5900),
.B(n_1265),
.C(n_1266),
.Y(n_6029)
);

AO211x2_ASAP7_75t_L g6030 ( 
.A1(n_5905),
.A2(n_1269),
.B(n_1266),
.C(n_1268),
.Y(n_6030)
);

AOI221x1_ASAP7_75t_L g6031 ( 
.A1(n_5896),
.A2(n_1270),
.B1(n_1268),
.B2(n_1269),
.C(n_1271),
.Y(n_6031)
);

NOR3xp33_ASAP7_75t_L g6032 ( 
.A(n_5944),
.B(n_1271),
.C(n_1273),
.Y(n_6032)
);

OAI221xp5_ASAP7_75t_L g6033 ( 
.A1(n_5896),
.A2(n_1277),
.B1(n_1275),
.B2(n_1276),
.C(n_1278),
.Y(n_6033)
);

NAND2xp5_ASAP7_75t_L g6034 ( 
.A(n_5899),
.B(n_1279),
.Y(n_6034)
);

NAND4xp25_ASAP7_75t_L g6035 ( 
.A(n_5901),
.B(n_1687),
.C(n_1688),
.D(n_1685),
.Y(n_6035)
);

NOR4xp25_ASAP7_75t_L g6036 ( 
.A(n_5896),
.B(n_1283),
.C(n_1280),
.D(n_1281),
.Y(n_6036)
);

NOR3xp33_ASAP7_75t_L g6037 ( 
.A(n_5944),
.B(n_1284),
.C(n_1285),
.Y(n_6037)
);

OAI221xp5_ASAP7_75t_L g6038 ( 
.A1(n_5896),
.A2(n_1288),
.B1(n_1285),
.B2(n_1286),
.C(n_1290),
.Y(n_6038)
);

NAND2xp5_ASAP7_75t_SL g6039 ( 
.A(n_5901),
.B(n_1286),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5964),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5964),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5964),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5964),
.Y(n_6043)
);

OAI322xp33_ASAP7_75t_L g6044 ( 
.A1(n_5906),
.A2(n_1684),
.A3(n_1682),
.B1(n_1689),
.B2(n_1698),
.C1(n_1683),
.C2(n_1681),
.Y(n_6044)
);

OAI221xp5_ASAP7_75t_L g6045 ( 
.A1(n_5896),
.A2(n_1294),
.B1(n_1292),
.B2(n_1293),
.C(n_1295),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5977),
.B(n_1300),
.Y(n_6046)
);

OAI21xp33_ASAP7_75t_L g6047 ( 
.A1(n_6025),
.A2(n_1303),
.B(n_1304),
.Y(n_6047)
);

AOI21xp33_ASAP7_75t_L g6048 ( 
.A1(n_6002),
.A2(n_1676),
.B(n_1675),
.Y(n_6048)
);

AOI221x1_ASAP7_75t_L g6049 ( 
.A1(n_6040),
.A2(n_6041),
.B1(n_6043),
.B2(n_6042),
.C(n_5979),
.Y(n_6049)
);

A2O1A1Ixp33_ASAP7_75t_L g6050 ( 
.A1(n_5981),
.A2(n_1314),
.B(n_1312),
.C(n_1313),
.Y(n_6050)
);

AOI221x1_ASAP7_75t_L g6051 ( 
.A1(n_6008),
.A2(n_1316),
.B1(n_1314),
.B2(n_1315),
.C(n_1317),
.Y(n_6051)
);

AOI22xp5_ASAP7_75t_L g6052 ( 
.A1(n_6001),
.A2(n_1318),
.B1(n_1316),
.B2(n_1317),
.Y(n_6052)
);

INVx2_ASAP7_75t_L g6053 ( 
.A(n_6030),
.Y(n_6053)
);

AOI322xp5_ASAP7_75t_L g6054 ( 
.A1(n_5998),
.A2(n_1328),
.A3(n_1327),
.B1(n_1325),
.B2(n_1322),
.C1(n_1323),
.C2(n_1326),
.Y(n_6054)
);

NAND2xp5_ASAP7_75t_L g6055 ( 
.A(n_6013),
.B(n_1325),
.Y(n_6055)
);

INVxp67_ASAP7_75t_L g6056 ( 
.A(n_5992),
.Y(n_6056)
);

AOI221xp5_ASAP7_75t_L g6057 ( 
.A1(n_6036),
.A2(n_1331),
.B1(n_1329),
.B2(n_1330),
.C(n_1332),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_6017),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_6006),
.Y(n_6059)
);

AOI211xp5_ASAP7_75t_L g6060 ( 
.A1(n_5973),
.A2(n_1335),
.B(n_1333),
.C(n_1334),
.Y(n_6060)
);

OAI221xp5_ASAP7_75t_L g6061 ( 
.A1(n_5968),
.A2(n_1336),
.B1(n_1333),
.B2(n_1335),
.C(n_1337),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_L g6062 ( 
.A(n_5980),
.B(n_1336),
.Y(n_6062)
);

NAND2xp5_ASAP7_75t_L g6063 ( 
.A(n_5990),
.B(n_1337),
.Y(n_6063)
);

OAI22xp5_ASAP7_75t_L g6064 ( 
.A1(n_6033),
.A2(n_1341),
.B1(n_1339),
.B2(n_1340),
.Y(n_6064)
);

OAI21xp5_ASAP7_75t_L g6065 ( 
.A1(n_5996),
.A2(n_1339),
.B(n_1340),
.Y(n_6065)
);

OAI22xp33_ASAP7_75t_L g6066 ( 
.A1(n_5966),
.A2(n_1344),
.B1(n_1342),
.B2(n_1343),
.Y(n_6066)
);

AOI221xp5_ASAP7_75t_L g6067 ( 
.A1(n_5969),
.A2(n_1350),
.B1(n_1347),
.B2(n_1349),
.C(n_1351),
.Y(n_6067)
);

AOI211xp5_ASAP7_75t_L g6068 ( 
.A1(n_5967),
.A2(n_5976),
.B(n_5989),
.C(n_5986),
.Y(n_6068)
);

OAI21xp5_ASAP7_75t_SL g6069 ( 
.A1(n_6003),
.A2(n_1352),
.B(n_1353),
.Y(n_6069)
);

OAI22xp5_ASAP7_75t_L g6070 ( 
.A1(n_6038),
.A2(n_1356),
.B1(n_1354),
.B2(n_1355),
.Y(n_6070)
);

NOR2xp33_ASAP7_75t_SL g6071 ( 
.A(n_6044),
.B(n_1355),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_6012),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5975),
.Y(n_6073)
);

AOI21xp33_ASAP7_75t_L g6074 ( 
.A1(n_5970),
.A2(n_1671),
.B(n_1670),
.Y(n_6074)
);

OAI22xp5_ASAP7_75t_L g6075 ( 
.A1(n_6045),
.A2(n_1360),
.B1(n_1358),
.B2(n_1359),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_6018),
.Y(n_6076)
);

AOI221xp5_ASAP7_75t_L g6077 ( 
.A1(n_5994),
.A2(n_1365),
.B1(n_1363),
.B2(n_1364),
.C(n_1367),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_6031),
.B(n_1368),
.Y(n_6078)
);

NAND2xp33_ASAP7_75t_L g6079 ( 
.A(n_5974),
.B(n_1369),
.Y(n_6079)
);

O2A1O1Ixp33_ASAP7_75t_L g6080 ( 
.A1(n_6026),
.A2(n_6029),
.B(n_6034),
.C(n_6028),
.Y(n_6080)
);

AOI22xp5_ASAP7_75t_L g6081 ( 
.A1(n_5971),
.A2(n_1375),
.B1(n_1371),
.B2(n_1374),
.Y(n_6081)
);

HB1xp67_ASAP7_75t_L g6082 ( 
.A(n_5985),
.Y(n_6082)
);

INVx2_ASAP7_75t_L g6083 ( 
.A(n_5972),
.Y(n_6083)
);

NAND2xp33_ASAP7_75t_L g6084 ( 
.A(n_6032),
.B(n_1381),
.Y(n_6084)
);

AOI22xp5_ASAP7_75t_L g6085 ( 
.A1(n_6020),
.A2(n_1383),
.B1(n_1381),
.B2(n_1382),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_5997),
.B(n_1383),
.Y(n_6086)
);

OAI221xp5_ASAP7_75t_L g6087 ( 
.A1(n_6024),
.A2(n_1389),
.B1(n_1387),
.B2(n_1388),
.C(n_1390),
.Y(n_6087)
);

AOI21xp5_ASAP7_75t_L g6088 ( 
.A1(n_6027),
.A2(n_1387),
.B(n_1388),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5982),
.Y(n_6089)
);

OAI221xp5_ASAP7_75t_L g6090 ( 
.A1(n_6014),
.A2(n_1397),
.B1(n_1395),
.B2(n_1396),
.C(n_1398),
.Y(n_6090)
);

OR2x2_ASAP7_75t_L g6091 ( 
.A(n_6039),
.B(n_6035),
.Y(n_6091)
);

O2A1O1Ixp33_ASAP7_75t_L g6092 ( 
.A1(n_6037),
.A2(n_1403),
.B(n_1401),
.C(n_1402),
.Y(n_6092)
);

AOI21xp33_ASAP7_75t_L g6093 ( 
.A1(n_6023),
.A2(n_1673),
.B(n_1672),
.Y(n_6093)
);

AOI322xp5_ASAP7_75t_L g6094 ( 
.A1(n_6009),
.A2(n_1411),
.A3(n_1409),
.B1(n_1406),
.B2(n_1402),
.C1(n_1404),
.C2(n_1408),
.Y(n_6094)
);

INVx2_ASAP7_75t_L g6095 ( 
.A(n_6053),
.Y(n_6095)
);

O2A1O1Ixp33_ASAP7_75t_L g6096 ( 
.A1(n_6050),
.A2(n_5984),
.B(n_6021),
.C(n_5983),
.Y(n_6096)
);

OAI222xp33_ASAP7_75t_L g6097 ( 
.A1(n_6082),
.A2(n_6015),
.B1(n_6010),
.B2(n_5993),
.C1(n_5995),
.C2(n_5991),
.Y(n_6097)
);

OAI211xp5_ASAP7_75t_L g6098 ( 
.A1(n_6049),
.A2(n_6016),
.B(n_5988),
.C(n_5987),
.Y(n_6098)
);

OAI21xp33_ASAP7_75t_L g6099 ( 
.A1(n_6071),
.A2(n_6083),
.B(n_6069),
.Y(n_6099)
);

O2A1O1Ixp33_ASAP7_75t_L g6100 ( 
.A1(n_6086),
.A2(n_6000),
.B(n_5999),
.C(n_6004),
.Y(n_6100)
);

INVxp67_ASAP7_75t_L g6101 ( 
.A(n_6078),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_6055),
.Y(n_6102)
);

BUFx12f_ASAP7_75t_L g6103 ( 
.A(n_6046),
.Y(n_6103)
);

O2A1O1Ixp33_ASAP7_75t_SL g6104 ( 
.A1(n_6076),
.A2(n_6022),
.B(n_5978),
.C(n_6007),
.Y(n_6104)
);

AND2x2_ASAP7_75t_L g6105 ( 
.A(n_6073),
.B(n_6019),
.Y(n_6105)
);

AOI21xp5_ASAP7_75t_L g6106 ( 
.A1(n_6063),
.A2(n_6005),
.B(n_6011),
.Y(n_6106)
);

INVx2_ASAP7_75t_SL g6107 ( 
.A(n_6091),
.Y(n_6107)
);

AOI21xp5_ASAP7_75t_L g6108 ( 
.A1(n_6088),
.A2(n_6066),
.B(n_6047),
.Y(n_6108)
);

AOI221xp5_ASAP7_75t_L g6109 ( 
.A1(n_6080),
.A2(n_1414),
.B1(n_1412),
.B2(n_1413),
.C(n_1415),
.Y(n_6109)
);

O2A1O1Ixp33_ASAP7_75t_L g6110 ( 
.A1(n_6048),
.A2(n_1415),
.B(n_1412),
.C(n_1413),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_6062),
.Y(n_6111)
);

NAND2xp5_ASAP7_75t_L g6112 ( 
.A(n_6051),
.B(n_1416),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_6058),
.Y(n_6113)
);

INVxp67_ASAP7_75t_SL g6114 ( 
.A(n_6068),
.Y(n_6114)
);

NAND2xp5_ASAP7_75t_L g6115 ( 
.A(n_6054),
.B(n_1417),
.Y(n_6115)
);

OAI221xp5_ASAP7_75t_L g6116 ( 
.A1(n_6065),
.A2(n_1419),
.B1(n_1417),
.B2(n_1418),
.C(n_1420),
.Y(n_6116)
);

OAI21xp5_ASAP7_75t_L g6117 ( 
.A1(n_6056),
.A2(n_1418),
.B(n_1421),
.Y(n_6117)
);

CKINVDCx5p33_ASAP7_75t_R g6118 ( 
.A(n_6059),
.Y(n_6118)
);

OAI31xp33_ASAP7_75t_L g6119 ( 
.A1(n_6089),
.A2(n_1423),
.A3(n_1421),
.B(n_1422),
.Y(n_6119)
);

OAI21xp5_ASAP7_75t_SL g6120 ( 
.A1(n_6074),
.A2(n_1422),
.B(n_1423),
.Y(n_6120)
);

AOI221xp5_ASAP7_75t_L g6121 ( 
.A1(n_6072),
.A2(n_1429),
.B1(n_1426),
.B2(n_1427),
.C(n_1430),
.Y(n_6121)
);

OAI21xp5_ASAP7_75t_SL g6122 ( 
.A1(n_6067),
.A2(n_1431),
.B(n_1432),
.Y(n_6122)
);

AOI221xp5_ASAP7_75t_L g6123 ( 
.A1(n_6057),
.A2(n_1436),
.B1(n_1434),
.B2(n_1435),
.C(n_1437),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_6081),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_6060),
.B(n_1701),
.Y(n_6125)
);

O2A1O1Ixp33_ASAP7_75t_L g6126 ( 
.A1(n_6079),
.A2(n_1441),
.B(n_1439),
.C(n_1440),
.Y(n_6126)
);

AND2x2_ASAP7_75t_SL g6127 ( 
.A(n_6112),
.B(n_6084),
.Y(n_6127)
);

NOR4xp25_ASAP7_75t_L g6128 ( 
.A(n_6099),
.B(n_6093),
.C(n_6061),
.D(n_6092),
.Y(n_6128)
);

NOR3x1_ASAP7_75t_L g6129 ( 
.A(n_6114),
.B(n_6087),
.C(n_6090),
.Y(n_6129)
);

AOI22xp5_ASAP7_75t_SL g6130 ( 
.A1(n_6118),
.A2(n_6070),
.B1(n_6075),
.B2(n_6064),
.Y(n_6130)
);

INVx2_ASAP7_75t_L g6131 ( 
.A(n_6103),
.Y(n_6131)
);

OAI21xp5_ASAP7_75t_SL g6132 ( 
.A1(n_6098),
.A2(n_6097),
.B(n_6107),
.Y(n_6132)
);

INVx2_ASAP7_75t_SL g6133 ( 
.A(n_6105),
.Y(n_6133)
);

OAI21xp5_ASAP7_75t_L g6134 ( 
.A1(n_6096),
.A2(n_6094),
.B(n_6077),
.Y(n_6134)
);

INVx1_ASAP7_75t_L g6135 ( 
.A(n_6111),
.Y(n_6135)
);

NOR3xp33_ASAP7_75t_L g6136 ( 
.A(n_6101),
.B(n_6085),
.C(n_6052),
.Y(n_6136)
);

INVx2_ASAP7_75t_SL g6137 ( 
.A(n_6113),
.Y(n_6137)
);

OAI22xp5_ASAP7_75t_SL g6138 ( 
.A1(n_6116),
.A2(n_1444),
.B1(n_1442),
.B2(n_1443),
.Y(n_6138)
);

O2A1O1Ixp33_ASAP7_75t_L g6139 ( 
.A1(n_6102),
.A2(n_1445),
.B(n_1443),
.C(n_1444),
.Y(n_6139)
);

NAND5xp2_ASAP7_75t_L g6140 ( 
.A(n_6100),
.B(n_1448),
.C(n_1446),
.D(n_1447),
.E(n_1449),
.Y(n_6140)
);

AOI221xp5_ASAP7_75t_L g6141 ( 
.A1(n_6104),
.A2(n_1451),
.B1(n_1446),
.B2(n_1450),
.C(n_1452),
.Y(n_6141)
);

AOI22xp5_ASAP7_75t_L g6142 ( 
.A1(n_6095),
.A2(n_1453),
.B1(n_1450),
.B2(n_1452),
.Y(n_6142)
);

AOI211xp5_ASAP7_75t_L g6143 ( 
.A1(n_6108),
.A2(n_1457),
.B(n_1455),
.C(n_1456),
.Y(n_6143)
);

AOI31xp33_ASAP7_75t_L g6144 ( 
.A1(n_6117),
.A2(n_1460),
.A3(n_1456),
.B(n_1459),
.Y(n_6144)
);

NOR2x1_ASAP7_75t_L g6145 ( 
.A(n_6115),
.B(n_6125),
.Y(n_6145)
);

OAI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_6110),
.A2(n_6126),
.B(n_6106),
.Y(n_6146)
);

NOR2x1_ASAP7_75t_L g6147 ( 
.A(n_6132),
.B(n_6120),
.Y(n_6147)
);

INVxp33_ASAP7_75t_L g6148 ( 
.A(n_6130),
.Y(n_6148)
);

NOR2x1_ASAP7_75t_L g6149 ( 
.A(n_6131),
.B(n_6122),
.Y(n_6149)
);

INVxp67_ASAP7_75t_L g6150 ( 
.A(n_6140),
.Y(n_6150)
);

AOI22xp5_ASAP7_75t_L g6151 ( 
.A1(n_6145),
.A2(n_6124),
.B1(n_6123),
.B2(n_6109),
.Y(n_6151)
);

NOR2x1_ASAP7_75t_L g6152 ( 
.A(n_6135),
.B(n_6119),
.Y(n_6152)
);

AO22x2_ASAP7_75t_L g6153 ( 
.A1(n_6133),
.A2(n_6121),
.B1(n_1464),
.B2(n_1462),
.Y(n_6153)
);

AND2x4_ASAP7_75t_L g6154 ( 
.A(n_6137),
.B(n_1463),
.Y(n_6154)
);

INVx1_ASAP7_75t_L g6155 ( 
.A(n_6127),
.Y(n_6155)
);

AOI22xp5_ASAP7_75t_L g6156 ( 
.A1(n_6136),
.A2(n_1468),
.B1(n_1466),
.B2(n_1467),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_6138),
.Y(n_6157)
);

AND3x1_ASAP7_75t_L g6158 ( 
.A(n_6149),
.B(n_6141),
.C(n_6143),
.Y(n_6158)
);

NOR2x1_ASAP7_75t_L g6159 ( 
.A(n_6154),
.B(n_6139),
.Y(n_6159)
);

AOI221xp5_ASAP7_75t_L g6160 ( 
.A1(n_6150),
.A2(n_6128),
.B1(n_6146),
.B2(n_6134),
.C(n_6144),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_6153),
.Y(n_6161)
);

AND2x2_ASAP7_75t_L g6162 ( 
.A(n_6155),
.B(n_6129),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_6147),
.Y(n_6163)
);

NAND2x1p5_ASAP7_75t_L g6164 ( 
.A(n_6152),
.B(n_6142),
.Y(n_6164)
);

OR2x2_ASAP7_75t_L g6165 ( 
.A(n_6148),
.B(n_6157),
.Y(n_6165)
);

OAI21xp33_ASAP7_75t_L g6166 ( 
.A1(n_6163),
.A2(n_6151),
.B(n_6156),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_6164),
.Y(n_6167)
);

AOI22xp5_ASAP7_75t_L g6168 ( 
.A1(n_6161),
.A2(n_6158),
.B1(n_6159),
.B2(n_6162),
.Y(n_6168)
);

AOI211xp5_ASAP7_75t_SL g6169 ( 
.A1(n_6165),
.A2(n_1474),
.B(n_1472),
.C(n_1473),
.Y(n_6169)
);

NAND5xp2_ASAP7_75t_L g6170 ( 
.A(n_6160),
.B(n_1475),
.C(n_1472),
.D(n_1474),
.E(n_1476),
.Y(n_6170)
);

BUFx2_ASAP7_75t_L g6171 ( 
.A(n_6167),
.Y(n_6171)
);

XOR2xp5_ASAP7_75t_L g6172 ( 
.A(n_6171),
.B(n_6168),
.Y(n_6172)
);

HB1xp67_ASAP7_75t_L g6173 ( 
.A(n_6172),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_6173),
.Y(n_6174)
);

INVx1_ASAP7_75t_SL g6175 ( 
.A(n_6174),
.Y(n_6175)
);

OAI21xp5_ASAP7_75t_SL g6176 ( 
.A1(n_6175),
.A2(n_6166),
.B(n_6169),
.Y(n_6176)
);

OAI31xp33_ASAP7_75t_L g6177 ( 
.A1(n_6176),
.A2(n_6170),
.A3(n_1482),
.B(n_1480),
.Y(n_6177)
);

AOI222xp33_ASAP7_75t_L g6178 ( 
.A1(n_6177),
.A2(n_1483),
.B1(n_1485),
.B2(n_1481),
.C1(n_1482),
.C2(n_1484),
.Y(n_6178)
);

AOI22xp5_ASAP7_75t_SL g6179 ( 
.A1(n_6178),
.A2(n_1487),
.B1(n_1485),
.B2(n_1486),
.Y(n_6179)
);

OR2x6_ASAP7_75t_L g6180 ( 
.A(n_6179),
.B(n_1486),
.Y(n_6180)
);

AOI21xp33_ASAP7_75t_SL g6181 ( 
.A1(n_6180),
.A2(n_1488),
.B(n_1489),
.Y(n_6181)
);

AOI211xp5_ASAP7_75t_L g6182 ( 
.A1(n_6181),
.A2(n_1700),
.B(n_1490),
.C(n_1489),
.Y(n_6182)
);


endmodule