module fake_netlist_6_650_n_106 (n_7, n_6, n_12, n_4, n_2, n_15, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_10, n_106);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_106;

wire n_52;
wire n_16;
wire n_91;
wire n_46;
wire n_21;
wire n_18;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_17;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_25;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVxp67_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OR2x6_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_27),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_26),
.B1(n_16),
.B2(n_28),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_35),
.B(n_41),
.C(n_34),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_36),
.B(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_30),
.B1(n_24),
.B2(n_18),
.Y(n_55)
);

CKINVDCx10_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_55),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_50),
.B(n_47),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_51),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_45),
.B(n_43),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_46),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_42),
.B(n_34),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_31),
.B(n_51),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_2),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_13),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_31),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NAND2x1_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_59),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_69),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_68),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_64),
.Y(n_83)
);

AOI211xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_65),
.B(n_64),
.C(n_62),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_75),
.B(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_65),
.B1(n_80),
.B2(n_66),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_65),
.B1(n_67),
.B2(n_66),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_66),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_84),
.B(n_87),
.Y(n_91)
);

AOI222xp33_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_87),
.B1(n_60),
.B2(n_66),
.C1(n_62),
.C2(n_7),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_88),
.B1(n_62),
.B2(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NOR4xp25_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_63),
.B(n_61),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_96),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_SL g103 ( 
.A(n_101),
.B(n_96),
.C(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_103),
.B1(n_67),
.B2(n_61),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_61),
.B(n_7),
.Y(n_106)
);


endmodule