module fake_jpeg_24336_n_230 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_33),
.B1(n_21),
.B2(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_26),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_17),
.B1(n_20),
.B2(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_13),
.B1(n_26),
.B2(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_60),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_36),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_36),
.B(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_62),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_71),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_87),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_57),
.B(n_58),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_83),
.B(n_85),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_89),
.B1(n_29),
.B2(n_60),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_65),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_18),
.B(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_14),
.B1(n_18),
.B2(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_39),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_19),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_70),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_102),
.B(n_82),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_39),
.B1(n_33),
.B2(n_31),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_90),
.B1(n_29),
.B2(n_84),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_31),
.B1(n_33),
.B2(n_45),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_106),
.B1(n_90),
.B2(n_62),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_52),
.C(n_48),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_112),
.C(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_35),
.C(n_44),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_129),
.C(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_120),
.B1(n_121),
.B2(n_130),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_82),
.B1(n_84),
.B2(n_78),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_102),
.B1(n_101),
.B2(n_104),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_75),
.B(n_78),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_80),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_87),
.C(n_88),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_91),
.B1(n_86),
.B2(n_19),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_71),
.B(n_69),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_22),
.B(n_15),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_95),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_107),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_152),
.B1(n_121),
.B2(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_98),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_91),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_99),
.B1(n_68),
.B2(n_22),
.Y(n_152)
);

INVxp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_129),
.C(n_131),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_147),
.C(n_135),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_114),
.B1(n_128),
.B2(n_116),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_142),
.B(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_168),
.B1(n_134),
.B2(n_148),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_133),
.B1(n_129),
.B2(n_114),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_172),
.C(n_179),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_181),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_180),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_128),
.B(n_152),
.C(n_116),
.D(n_35),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_177),
.B(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_44),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_15),
.C(n_23),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_16),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_24),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_153),
.B(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_159),
.B(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_153),
.B1(n_158),
.B2(n_165),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_193),
.B1(n_154),
.B2(n_35),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_0),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_154),
.B1(n_164),
.B2(n_55),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_184),
.B1(n_192),
.B2(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_24),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_200),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_8),
.B(n_1),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_204),
.B(n_2),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_24),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_24),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_204),
.C(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_8),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_7),
.B(n_2),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_23),
.C(n_14),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_193),
.B1(n_190),
.B2(n_183),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_195),
.C(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_9),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_9),
.B(n_3),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_3),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_4),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_5),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_222),
.C(n_5),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_226),
.B(n_10),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_10),
.C(n_11),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_11),
.C(n_12),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_0),
.B1(n_12),
.B2(n_216),
.Y(n_230)
);


endmodule