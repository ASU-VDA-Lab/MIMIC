module fake_ibex_1833_n_1420 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_105, n_187, n_1, n_154, n_182, n_196, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_57, n_301, n_296, n_120, n_168, n_155, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_55, n_291, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_119, n_72, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1420);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_55;
input n_291;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_119;
input n_72;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1420;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_891;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_1339;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_716;
wire n_923;
wire n_642;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_804;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1374;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1361;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_288),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_277),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_268),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_182),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_190),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_208),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_186),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_174),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_166),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_281),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_167),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_34),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_168),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_175),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_27),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_250),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_224),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_122),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_99),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_61),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_173),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_142),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_92),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_113),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_70),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_226),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_229),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_156),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_64),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_312),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_17),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_41),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_94),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_133),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_213),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_4),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_120),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_209),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_131),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_179),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_127),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_188),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_265),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_153),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_161),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_146),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_274),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_283),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_272),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_241),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_126),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_255),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_220),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_53),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_163),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_165),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_87),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_238),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_143),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_297),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_185),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_66),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_176),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_22),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_290),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_172),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_38),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_144),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_4),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_71),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_210),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_75),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_202),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_0),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_256),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_31),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_292),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_287),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_96),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_111),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_299),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_259),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_178),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_222),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_157),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_95),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_245),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_254),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_253),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_70),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_233),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_199),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_106),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_151),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_73),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_7),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_291),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_232),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_278),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_116),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_214),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_263),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_99),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_267),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_107),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_273),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_302),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_148),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_311),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_269),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_203),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_285),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_200),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_249),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_81),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_42),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_252),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_115),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_134),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_293),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_270),
.Y(n_441)
);

BUFx8_ASAP7_75t_SL g442 ( 
.A(n_279),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_239),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_170),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_294),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_114),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_204),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_271),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_158),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_298),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_128),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_261),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_196),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_56),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_78),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_93),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_286),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_66),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_205),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_88),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_240),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_284),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_149),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_29),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_125),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_81),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_295),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_280),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_212),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_309),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_211),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_155),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_307),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_39),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_52),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_47),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_110),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_25),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_71),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_51),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_46),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_236),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_223),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_169),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_83),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_160),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_304),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_121),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_86),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_109),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_177),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_192),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_104),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_219),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_9),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_38),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_296),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_289),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_306),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_234),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_201),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_129),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_92),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_42),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_246),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_187),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_251),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_218),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_300),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_154),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_96),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_257),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_310),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_266),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_282),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_262),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_164),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_207),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_46),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_206),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_356),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_520),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_352),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_0),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_329),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_442),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_352),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_478),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_442),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_370),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_317),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_394),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_333),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_313),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_482),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_313),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_410),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_337),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_1),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_337),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_498),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_318),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_334),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_328),
.B(n_1),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_320),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_330),
.B(n_2),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_424),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_318),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_424),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_425),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_425),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_426),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_426),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_339),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_325),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_440),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_503),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_421),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_345),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_374),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_321),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_421),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_382),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_343),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_455),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_346),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_384),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_349),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_455),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_387),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_389),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_390),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_377),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_392),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_396),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_406),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_399),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_415),
.Y(n_589)
);

INVxp33_ASAP7_75t_SL g590 ( 
.A(n_416),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_423),
.Y(n_591)
);

INVxp33_ASAP7_75t_SL g592 ( 
.A(n_435),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_586),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_586),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_586),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_544),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_591),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_567),
.B(n_571),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_534),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_551),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_570),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_540),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_522),
.B(n_515),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_565),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_548),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_542),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_545),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_553),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_554),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_523),
.B(n_454),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_575),
.B(n_321),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_582),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_561),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_587),
.B(n_368),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_562),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_524),
.A2(n_458),
.B1(n_466),
.B2(n_460),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_563),
.B(n_368),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_577),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_547),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_559),
.B(n_393),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_535),
.B(n_568),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_549),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_572),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_569),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_585),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_525),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_576),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_579),
.B(n_441),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_526),
.B(n_372),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_580),
.B(n_441),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_581),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_583),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_584),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_590),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_574),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_574),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_524),
.A2(n_474),
.B1(n_480),
.B2(n_475),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_578),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_550),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_552),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_589),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_556),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_589),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_557),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_558),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_560),
.B(n_372),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_564),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_531),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_537),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_543),
.B(n_484),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_536),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_536),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_538),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_538),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_555),
.B(n_496),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_528),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_529),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_541),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_586),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_504),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_586),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_541),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_541),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_541),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_586),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_541),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_541),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_541),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_541),
.Y(n_689)
);

BUFx8_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_548),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_541),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_532),
.B(n_484),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_532),
.B(n_508),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_586),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_541),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_541),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_586),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_541),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_586),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_586),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_541),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_586),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_532),
.B(n_519),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_591),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_541),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_586),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_592),
.B(n_314),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_541),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_586),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_541),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_541),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_586),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_591),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_521),
.B(n_315),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_521),
.B(n_316),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_586),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_548),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_541),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_681),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_631),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_707),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_634),
.B(n_633),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_635),
.B(n_320),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_603),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_681),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_681),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_633),
.A2(n_479),
.B1(n_485),
.B2(n_481),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_720),
.Y(n_731)
);

BUFx4f_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_690),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_634),
.B(n_319),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_607),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_720),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_634),
.B(n_365),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_630),
.B(n_323),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_626),
.B(n_430),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_720),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_675),
.B(n_324),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_716),
.A2(n_495),
.B1(n_489),
.B2(n_493),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_610),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_608),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_690),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_630),
.B(n_326),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_630),
.B(n_327),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_630),
.B(n_331),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_616),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_597),
.B(n_716),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_675),
.B(n_355),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_597),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_685),
.B(n_332),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_622),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_674),
.B(n_335),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_622),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_685),
.B(n_355),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_608),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_635),
.B(n_398),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_679),
.B(n_338),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_340),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_594),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_686),
.B(n_341),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_612),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_616),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_680),
.B(n_342),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_624),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_600),
.B(n_398),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_639),
.B(n_505),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_682),
.A2(n_336),
.B1(n_348),
.B2(n_347),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_611),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_615),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_624),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_700),
.B(n_344),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_632),
.B(n_505),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_624),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_627),
.B(n_453),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_620),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_632),
.B(n_468),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_683),
.B(n_358),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_598),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_708),
.B(n_359),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_611),
.Y(n_784)
);

CKINVDCx8_ASAP7_75t_R g785 ( 
.A(n_670),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_624),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_R g787 ( 
.A(n_652),
.B(n_364),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_629),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_596),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_628),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_601),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_639),
.B(n_350),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_596),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_602),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_668),
.B(n_3),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_606),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_721),
.B(n_367),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_687),
.B(n_371),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_603),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_688),
.B(n_351),
.Y(n_800)
);

AND2x2_ASAP7_75t_SL g801 ( 
.A(n_710),
.B(n_353),
.Y(n_801)
);

BUFx10_ASAP7_75t_L g802 ( 
.A(n_645),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_645),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_645),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_689),
.A2(n_354),
.B1(n_360),
.B2(n_357),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_605),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_605),
.Y(n_807)
);

BUFx8_ASAP7_75t_SL g808 ( 
.A(n_670),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_614),
.B(n_375),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_619),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_692),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_599),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_599),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_696),
.B(n_361),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_640),
.B(n_362),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_599),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_599),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_697),
.B(n_378),
.Y(n_818)
);

AO22x2_ASAP7_75t_L g819 ( 
.A1(n_664),
.A2(n_366),
.B1(n_369),
.B2(n_363),
.Y(n_819)
);

HAxp5_ASAP7_75t_SL g820 ( 
.A(n_673),
.B(n_373),
.CON(n_820),
.SN(n_820)
);

AO21x2_ASAP7_75t_L g821 ( 
.A1(n_618),
.A2(n_621),
.B(n_625),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_691),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_604),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_706),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_604),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_604),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_698),
.B(n_380),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_604),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_703),
.B(n_381),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_643),
.B(n_383),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_691),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_598),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_704),
.B(n_385),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_711),
.B(n_388),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_651),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_713),
.B(n_401),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_714),
.B(n_404),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_618),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_594),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_637),
.B(n_405),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_594),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_637),
.B(n_717),
.Y(n_842)
);

OR2x2_ASAP7_75t_SL g843 ( 
.A(n_670),
.B(n_376),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_594),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_641),
.B(n_379),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_718),
.B(n_407),
.Y(n_846)
);

AO22x2_ASAP7_75t_L g847 ( 
.A1(n_664),
.A2(n_395),
.B1(n_400),
.B2(n_386),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_609),
.A2(n_403),
.B1(n_409),
.B2(n_402),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_647),
.Y(n_849)
);

XOR2xp5_ASAP7_75t_L g850 ( 
.A(n_623),
.B(n_3),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_609),
.B(n_408),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_636),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_642),
.B(n_411),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_638),
.B(n_417),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_651),
.Y(n_855)
);

BUFx4f_ASAP7_75t_L g856 ( 
.A(n_655),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_651),
.Y(n_857)
);

CKINVDCx8_ASAP7_75t_R g858 ( 
.A(n_670),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_693),
.B(n_412),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_625),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_649),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_702),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_617),
.B(n_414),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_677),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_652),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_SL g866 ( 
.A1(n_654),
.A2(n_427),
.B1(n_429),
.B2(n_422),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_593),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_694),
.B(n_432),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_709),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_659),
.A2(n_420),
.B1(n_428),
.B2(n_419),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_659),
.B(n_431),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_593),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_709),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_595),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_709),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_661),
.B(n_434),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_669),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_595),
.Y(n_878)
);

INVx6_ASAP7_75t_L g879 ( 
.A(n_655),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_676),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_655),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_663),
.B(n_518),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_678),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_678),
.Y(n_884)
);

AND2x6_ASAP7_75t_L g885 ( 
.A(n_662),
.B(n_657),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_669),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_653),
.B(n_445),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_684),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_657),
.B(n_448),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_662),
.B(n_450),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_695),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_699),
.Y(n_892)
);

AND2x4_ASAP7_75t_SL g893 ( 
.A(n_653),
.B(n_646),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_701),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_654),
.B(n_5),
.Y(n_895)
);

AO22x2_ASAP7_75t_L g896 ( 
.A1(n_665),
.A2(n_438),
.B1(n_443),
.B2(n_437),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_658),
.B(n_451),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_701),
.Y(n_898)
);

AO22x2_ASAP7_75t_L g899 ( 
.A1(n_850),
.A2(n_752),
.B1(n_667),
.B2(n_666),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_725),
.Y(n_900)
);

AO22x2_ASAP7_75t_L g901 ( 
.A1(n_750),
.A2(n_672),
.B1(n_671),
.B2(n_656),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_723),
.B(n_648),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_733),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_811),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_735),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_743),
.Y(n_906)
);

OAI221xp5_ASAP7_75t_L g907 ( 
.A1(n_788),
.A2(n_644),
.B1(n_660),
.B2(n_650),
.C(n_447),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_855),
.B(n_644),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_807),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_722),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_810),
.Y(n_912)
);

INVx3_ASAP7_75t_R g913 ( 
.A(n_724),
.Y(n_913)
);

AO22x2_ASAP7_75t_L g914 ( 
.A1(n_745),
.A2(n_757),
.B1(n_751),
.B2(n_792),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_736),
.Y(n_915)
);

AO22x2_ASAP7_75t_L g916 ( 
.A1(n_751),
.A2(n_446),
.B1(n_449),
.B2(n_444),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_791),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_857),
.B(n_452),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_740),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_SL g920 ( 
.A(n_877),
.B(n_459),
.C(n_457),
.Y(n_920)
);

OAI221xp5_ASAP7_75t_L g921 ( 
.A1(n_842),
.A2(n_470),
.B1(n_472),
.B2(n_467),
.C(n_462),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_864),
.A2(n_491),
.B1(n_501),
.B2(n_490),
.C(n_488),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_794),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_849),
.B(n_502),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_796),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_849),
.B(n_461),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_744),
.Y(n_927)
);

AO22x2_ASAP7_75t_L g928 ( 
.A1(n_757),
.A2(n_516),
.B1(n_517),
.B2(n_514),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_783),
.B(n_463),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_758),
.Y(n_930)
);

OAI221xp5_ASAP7_75t_L g931 ( 
.A1(n_730),
.A2(n_418),
.B1(n_483),
.B2(n_477),
.C(n_391),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_L g932 ( 
.A(n_815),
.B(n_465),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_754),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_808),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_772),
.Y(n_935)
);

AO22x2_ASAP7_75t_L g936 ( 
.A1(n_895),
.A2(n_477),
.B1(n_483),
.B2(n_418),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_756),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_764),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_778),
.A2(n_507),
.B(n_712),
.C(n_705),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_790),
.B(n_852),
.Y(n_940)
);

OAI221xp5_ASAP7_75t_L g941 ( 
.A1(n_805),
.A2(n_473),
.B1(n_486),
.B2(n_471),
.C(n_469),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_800),
.B(n_814),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_784),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_865),
.B(n_5),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_876),
.B(n_487),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_780),
.B(n_6),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_770),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_845),
.A2(n_497),
.B1(n_500),
.B2(n_492),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_773),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_799),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_779),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_785),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_814),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_856),
.B(n_322),
.Y(n_954)
);

AO22x2_ASAP7_75t_L g955 ( 
.A1(n_820),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_819),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_845),
.A2(n_509),
.B1(n_510),
.B2(n_506),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_819),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_893),
.B(n_8),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_824),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_847),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_847),
.Y(n_962)
);

OAI221xp5_ASAP7_75t_L g963 ( 
.A1(n_848),
.A2(n_513),
.B1(n_512),
.B2(n_715),
.C(n_712),
.Y(n_963)
);

AO22x2_ASAP7_75t_L g964 ( 
.A1(n_871),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_768),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_871),
.A2(n_896),
.B1(n_843),
.B2(n_771),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_835),
.B(n_11),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_838),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_856),
.B(n_322),
.Y(n_969)
);

AO22x2_ASAP7_75t_L g970 ( 
.A1(n_896),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_860),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_787),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_776),
.B(n_14),
.Y(n_973)
);

AO22x2_ASAP7_75t_L g974 ( 
.A1(n_795),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_830),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_806),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_854),
.B(n_16),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_821),
.Y(n_978)
);

OAI221xp5_ASAP7_75t_L g979 ( 
.A1(n_870),
.A2(n_719),
.B1(n_715),
.B2(n_439),
.C(n_499),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_742),
.B(n_18),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_834),
.B(n_18),
.Y(n_981)
);

OR2x2_ASAP7_75t_SL g982 ( 
.A(n_861),
.B(n_322),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_859),
.B(n_19),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_867),
.Y(n_984)
);

AO22x2_ASAP7_75t_L g985 ( 
.A1(n_801),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_894),
.Y(n_986)
);

AO22x2_ASAP7_75t_L g987 ( 
.A1(n_782),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_987)
);

AO22x2_ASAP7_75t_L g988 ( 
.A1(n_832),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_765),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_737),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_854),
.B(n_322),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_732),
.B(n_433),
.Y(n_992)
);

AO22x2_ASAP7_75t_L g993 ( 
.A1(n_881),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_882),
.B(n_433),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_732),
.B(n_433),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_741),
.Y(n_996)
);

AO22x2_ASAP7_75t_L g997 ( 
.A1(n_887),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_753),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_734),
.B(n_30),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_815),
.B(n_30),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_761),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_763),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_775),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_798),
.A2(n_719),
.B1(n_439),
.B2(n_499),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_815),
.B(n_31),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_803),
.B(n_804),
.Y(n_1006)
);

AO22x2_ASAP7_75t_L g1007 ( 
.A1(n_858),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_739),
.B(n_868),
.Y(n_1008)
);

AO22x2_ASAP7_75t_L g1009 ( 
.A1(n_755),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_822),
.B(n_831),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_879),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_886),
.B(n_840),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_885),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_885),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_802),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_885),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_853),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_853),
.B(n_863),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_809),
.Y(n_1019)
);

AO22x2_ASAP7_75t_L g1020 ( 
.A1(n_760),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_802),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_872),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_766),
.B(n_40),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_851),
.B(n_43),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_781),
.B(n_439),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_874),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_797),
.B(n_499),
.Y(n_1027)
);

AO22x2_ASAP7_75t_L g1028 ( 
.A1(n_818),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_846),
.B(n_44),
.Y(n_1029)
);

AO22x2_ASAP7_75t_L g1030 ( 
.A1(n_827),
.A2(n_49),
.B1(n_45),
.B2(n_48),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_866),
.B(n_49),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_878),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_900),
.B(n_829),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_913),
.B(n_728),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1008),
.B(n_833),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_960),
.B(n_897),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_975),
.B(n_728),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_904),
.B(n_729),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_942),
.B(n_836),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_967),
.B(n_729),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_SL g1041 ( 
.A(n_967),
.B(n_731),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_905),
.B(n_837),
.Y(n_1042)
);

NAND2xp33_ASAP7_75t_SL g1043 ( 
.A(n_972),
.B(n_889),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_SL g1044 ( 
.A(n_956),
.B(n_738),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1015),
.B(n_892),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_924),
.B(n_892),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_996),
.B(n_890),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_958),
.B(n_746),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_961),
.B(n_747),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_977),
.B(n_762),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_SL g1051 ( 
.A(n_962),
.B(n_748),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_944),
.B(n_816),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_948),
.B(n_762),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_998),
.B(n_816),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_957),
.B(n_762),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_1010),
.B(n_888),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_990),
.B(n_888),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_902),
.B(n_898),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_1017),
.B(n_777),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_959),
.B(n_786),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1001),
.B(n_1002),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1003),
.B(n_786),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_940),
.B(n_823),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_1018),
.B(n_823),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_910),
.B(n_812),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_906),
.B(n_726),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_1019),
.B(n_844),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_912),
.B(n_726),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_929),
.B(n_965),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_999),
.B(n_869),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_953),
.B(n_883),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_999),
.B(n_869),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_946),
.B(n_873),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_914),
.B(n_884),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_983),
.B(n_1023),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_SL g1077 ( 
.A(n_903),
.B(n_749),
.Y(n_1077)
);

NAND2xp33_ASAP7_75t_SL g1078 ( 
.A(n_952),
.B(n_749),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_SL g1079 ( 
.A(n_1000),
.B(n_767),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_SL g1080 ( 
.A(n_1005),
.B(n_767),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_950),
.B(n_774),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_981),
.B(n_880),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_SL g1083 ( 
.A(n_945),
.B(n_891),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_917),
.B(n_759),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_973),
.B(n_813),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_914),
.B(n_759),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_923),
.B(n_841),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_925),
.B(n_841),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_SL g1089 ( 
.A(n_1024),
.B(n_934),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_984),
.B(n_986),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_976),
.B(n_817),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1006),
.B(n_825),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_938),
.B(n_825),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_1031),
.B(n_826),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_SL g1095 ( 
.A(n_980),
.B(n_828),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_947),
.B(n_789),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_966),
.B(n_769),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_933),
.B(n_769),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_949),
.B(n_793),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_SL g1100 ( 
.A(n_951),
.B(n_839),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1029),
.B(n_875),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_SL g1102 ( 
.A(n_1022),
.B(n_862),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_899),
.B(n_50),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_916),
.B(n_50),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1026),
.B(n_51),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1032),
.B(n_954),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_916),
.B(n_52),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_969),
.B(n_53),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_992),
.B(n_54),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_995),
.B(n_54),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_928),
.B(n_55),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_908),
.B(n_55),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_SL g1113 ( 
.A(n_926),
.B(n_57),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_927),
.B(n_57),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_930),
.B(n_58),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_935),
.B(n_943),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1013),
.B(n_59),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_899),
.B(n_59),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1014),
.B(n_60),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_SL g1120 ( 
.A(n_918),
.B(n_60),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1016),
.B(n_61),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_937),
.B(n_62),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_SL g1123 ( 
.A(n_932),
.B(n_62),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_928),
.B(n_63),
.Y(n_1124)
);

NAND2xp33_ASAP7_75t_SL g1125 ( 
.A(n_982),
.B(n_65),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1011),
.B(n_65),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_978),
.B(n_108),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1101),
.A2(n_939),
.B(n_989),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1090),
.Y(n_1129)
);

CKINVDCx14_ASAP7_75t_R g1130 ( 
.A(n_1089),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1039),
.B(n_901),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1035),
.B(n_901),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_L g1133 ( 
.A(n_1041),
.B(n_993),
.Y(n_1133)
);

CKINVDCx14_ASAP7_75t_R g1134 ( 
.A(n_1034),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_1127),
.A2(n_1004),
.B(n_931),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1125),
.B(n_921),
.C(n_922),
.Y(n_1136)
);

CKINVDCx11_ASAP7_75t_R g1137 ( 
.A(n_1122),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1097),
.A2(n_936),
.B(n_993),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1066),
.A2(n_915),
.B(n_911),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1062),
.B(n_936),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_1122),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1036),
.B(n_971),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1054),
.Y(n_1143)
);

NOR4xp25_ASAP7_75t_L g1144 ( 
.A(n_1104),
.B(n_907),
.C(n_970),
.D(n_997),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1047),
.B(n_968),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1052),
.Y(n_1146)
);

BUFx8_ASAP7_75t_L g1147 ( 
.A(n_1103),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1068),
.A2(n_919),
.B(n_909),
.Y(n_1148)
);

OA22x2_ASAP7_75t_L g1149 ( 
.A1(n_1118),
.A2(n_994),
.B1(n_1027),
.B2(n_1025),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1042),
.A2(n_991),
.B(n_963),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1063),
.A2(n_920),
.B(n_1009),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1054),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1084),
.Y(n_1153)
);

AOI221x1_ASAP7_75t_L g1154 ( 
.A1(n_1095),
.A2(n_970),
.B1(n_985),
.B2(n_988),
.C(n_987),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1047),
.B(n_974),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1100),
.A2(n_1027),
.B(n_1025),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1084),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1033),
.A2(n_979),
.B(n_941),
.Y(n_1158)
);

AO22x1_ASAP7_75t_L g1159 ( 
.A1(n_1107),
.A2(n_987),
.B1(n_988),
.B2(n_985),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1071),
.A2(n_1020),
.B(n_1009),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1076),
.B(n_974),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1111),
.A2(n_997),
.B(n_955),
.C(n_964),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1102),
.A2(n_1028),
.B(n_1020),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1106),
.A2(n_1030),
.B(n_1028),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1046),
.B(n_964),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1098),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1077),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1074),
.A2(n_1030),
.B(n_1007),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1070),
.B(n_955),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1086),
.Y(n_1170)
);

NAND3x1_ASAP7_75t_L g1171 ( 
.A(n_1124),
.B(n_1007),
.C(n_67),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1072),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1082),
.A2(n_117),
.B(n_112),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1056),
.B(n_67),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1067),
.A2(n_119),
.B(n_118),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1075),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1073),
.A2(n_72),
.B1(n_68),
.B2(n_69),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1069),
.A2(n_68),
.B(n_69),
.Y(n_1178)
);

AO21x1_ASAP7_75t_L g1179 ( 
.A1(n_1123),
.A2(n_72),
.B(n_73),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1098),
.B(n_74),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1057),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1085),
.A2(n_124),
.B(n_123),
.Y(n_1182)
);

NAND3x1_ASAP7_75t_L g1183 ( 
.A(n_1043),
.B(n_76),
.C(n_77),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1094),
.A2(n_77),
.B(n_79),
.C(n_80),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1065),
.A2(n_1099),
.B(n_1096),
.Y(n_1185)
);

NAND2x1p5_ASAP7_75t_L g1186 ( 
.A(n_1040),
.B(n_80),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1116),
.A2(n_132),
.B(n_130),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1050),
.B(n_82),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1061),
.B(n_84),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1059),
.B(n_85),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1091),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1112),
.A2(n_88),
.B(n_89),
.Y(n_1192)
);

AO32x2_ASAP7_75t_L g1193 ( 
.A1(n_1044),
.A2(n_89),
.A3(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1064),
.B(n_97),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1093),
.Y(n_1195)
);

OAI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1144),
.A2(n_1120),
.B1(n_1113),
.B2(n_1105),
.C(n_1049),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1175),
.A2(n_1092),
.B(n_1060),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1163),
.A2(n_1048),
.B(n_1051),
.C(n_1078),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1172),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1154),
.A2(n_1179),
.A3(n_1128),
.B(n_1184),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1129),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1133),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1157),
.B(n_1058),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1156),
.A2(n_1080),
.B(n_1079),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1142),
.B(n_1176),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1165),
.A2(n_1171),
.B1(n_1149),
.B2(n_1141),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1132),
.B(n_1053),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1137),
.B(n_97),
.Y(n_1208)
);

OR2x6_ASAP7_75t_L g1209 ( 
.A(n_1159),
.B(n_1146),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1162),
.A2(n_1126),
.B(n_1114),
.C(n_1115),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1143),
.B(n_1045),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1195),
.Y(n_1212)
);

AOI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1138),
.A2(n_1119),
.B(n_1117),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1189),
.Y(n_1214)
);

AND2x2_ASAP7_75t_SL g1215 ( 
.A(n_1180),
.B(n_1108),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1191),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1152),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1191),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1131),
.B(n_1055),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1147),
.A2(n_1121),
.B1(n_1110),
.B2(n_1109),
.Y(n_1220)
);

AND2x6_ASAP7_75t_L g1221 ( 
.A(n_1170),
.B(n_1083),
.Y(n_1221)
);

AOI222xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1160),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.C1(n_102),
.C2(n_103),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1147),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1145),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1130),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1168),
.B(n_1038),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1164),
.A2(n_1088),
.B(n_1087),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1169),
.B(n_1037),
.Y(n_1228)
);

INVx6_ASAP7_75t_L g1229 ( 
.A(n_1153),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1155),
.B(n_102),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1188),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1174),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1201),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1205),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1216),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1202),
.Y(n_1236)
);

AOI21xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1206),
.A2(n_1167),
.B(n_1161),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1218),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1212),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1207),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1207),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1224),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_1217),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_1229),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1199),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1204),
.A2(n_1148),
.B(n_1185),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1204),
.A2(n_1151),
.B(n_1178),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1219),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1202),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1227),
.Y(n_1250)
);

BUFx2_ASAP7_75t_SL g1251 ( 
.A(n_1221),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1214),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1219),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1231),
.B(n_1232),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1226),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1226),
.Y(n_1256)
);

INVx5_ASAP7_75t_SL g1257 ( 
.A(n_1209),
.Y(n_1257)
);

NAND2x1_ASAP7_75t_L g1258 ( 
.A(n_1209),
.B(n_1157),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1197),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1210),
.A2(n_1136),
.B(n_1183),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1227),
.Y(n_1261)
);

NAND2xp33_ASAP7_75t_R g1262 ( 
.A(n_1236),
.B(n_1225),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1245),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1234),
.B(n_1208),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1242),
.B(n_1230),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1252),
.B(n_1209),
.Y(n_1266)
);

XOR2xp5_ASAP7_75t_L g1267 ( 
.A(n_1254),
.B(n_1223),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1235),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1236),
.Y(n_1269)
);

INVx8_ASAP7_75t_L g1270 ( 
.A(n_1243),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1244),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_R g1272 ( 
.A(n_1249),
.B(n_1134),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1248),
.B(n_1206),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1249),
.B(n_1228),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1258),
.B(n_1203),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1235),
.Y(n_1276)
);

NOR2xp67_ASAP7_75t_L g1277 ( 
.A(n_1237),
.B(n_1196),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1248),
.B(n_1140),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1251),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1258),
.B(n_1203),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1253),
.B(n_1223),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1253),
.B(n_1200),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1244),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_R g1284 ( 
.A(n_1240),
.B(n_1215),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1239),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1240),
.B(n_1198),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1241),
.B(n_1200),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1241),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1267),
.A2(n_1260),
.B1(n_1196),
.B2(n_1251),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1268),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1275),
.B(n_1255),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1276),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1285),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1263),
.B(n_1288),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1282),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1266),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1283),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1274),
.B(n_1238),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1269),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1265),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1273),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1277),
.A2(n_1237),
.B1(n_1257),
.B2(n_1220),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1278),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1271),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1281),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1287),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1272),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1286),
.B(n_1255),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1286),
.Y(n_1309)
);

AOI211xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1302),
.A2(n_1264),
.B(n_1280),
.C(n_1275),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1289),
.A2(n_1279),
.B(n_1270),
.C(n_1280),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1298),
.B(n_1233),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1309),
.B(n_1250),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1294),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1309),
.B(n_1250),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1290),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1299),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1295),
.B(n_1250),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1301),
.B(n_1238),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1296),
.B(n_1300),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1289),
.A2(n_1257),
.B1(n_1270),
.B2(n_1284),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1303),
.B(n_1233),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1290),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1317),
.B(n_1307),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1312),
.B(n_1295),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1320),
.B(n_1314),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1319),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1322),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1318),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1316),
.B(n_1305),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1323),
.B(n_1304),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1313),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1313),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1315),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1315),
.B(n_1306),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1310),
.B(n_1292),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1321),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1311),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1338),
.A2(n_1304),
.B1(n_1262),
.B2(n_1293),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1337),
.B(n_1292),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1327),
.B(n_1308),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1336),
.B(n_1308),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1326),
.B(n_1291),
.Y(n_1343)
);

AO221x2_ASAP7_75t_L g1344 ( 
.A1(n_1336),
.A2(n_1311),
.B1(n_1293),
.B2(n_1257),
.C(n_1222),
.Y(n_1344)
);

AO221x2_ASAP7_75t_L g1345 ( 
.A1(n_1338),
.A2(n_1257),
.B1(n_1222),
.B2(n_1271),
.C(n_1192),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1331),
.A2(n_1297),
.B1(n_1291),
.B2(n_1283),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1340),
.B(n_1325),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1339),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1342),
.A2(n_1324),
.B1(n_1331),
.B2(n_1332),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1343),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1348),
.A2(n_1349),
.B1(n_1346),
.B2(n_1350),
.C(n_1344),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1347),
.A2(n_1345),
.B1(n_1341),
.B2(n_1328),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1347),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1353),
.A2(n_1291),
.B1(n_1330),
.B2(n_1283),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1351),
.B(n_1333),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1352),
.B(n_1334),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1353),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1357),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1355),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1356),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1354),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1354),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1358),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1362),
.B(n_1359),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1361),
.B(n_1335),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1360),
.B(n_1297),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1358),
.B(n_1329),
.Y(n_1367)
);

NOR3xp33_ASAP7_75t_SL g1368 ( 
.A(n_1358),
.B(n_1194),
.C(n_1190),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1363),
.A2(n_1177),
.B(n_1186),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1367),
.Y(n_1370)
);

NAND4xp25_ASAP7_75t_L g1371 ( 
.A(n_1365),
.B(n_1210),
.C(n_1150),
.D(n_1158),
.Y(n_1371)
);

OAI21xp33_ASAP7_75t_L g1372 ( 
.A1(n_1366),
.A2(n_1297),
.B(n_1256),
.Y(n_1372)
);

OAI211xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1368),
.A2(n_105),
.B(n_106),
.C(n_1166),
.Y(n_1373)
);

NAND4xp25_ASAP7_75t_L g1374 ( 
.A(n_1364),
.B(n_1187),
.C(n_1173),
.D(n_1182),
.Y(n_1374)
);

XNOR2x1_ASAP7_75t_L g1375 ( 
.A(n_1364),
.B(n_1211),
.Y(n_1375)
);

NOR2x1_ASAP7_75t_L g1376 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_L g1377 ( 
.A(n_1375),
.B(n_1081),
.Y(n_1377)
);

NOR2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1371),
.B(n_1153),
.Y(n_1378)
);

OAI211xp5_ASAP7_75t_L g1379 ( 
.A1(n_1369),
.A2(n_1193),
.B(n_1247),
.C(n_1135),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1372),
.B(n_135),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1374),
.Y(n_1381)
);

NOR2xp67_ASAP7_75t_L g1382 ( 
.A(n_1370),
.B(n_136),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1370),
.Y(n_1383)
);

XNOR2xp5_ASAP7_75t_L g1384 ( 
.A(n_1376),
.B(n_1213),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1381),
.B(n_1181),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_R g1386 ( 
.A(n_1378),
.B(n_137),
.Y(n_1386)
);

NAND2xp33_ASAP7_75t_R g1387 ( 
.A(n_1380),
.B(n_138),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1377),
.B(n_139),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1379),
.B(n_1259),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_R g1390 ( 
.A(n_1381),
.B(n_140),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_SL g1391 ( 
.A(n_1383),
.B(n_141),
.C(n_145),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1382),
.B(n_1261),
.Y(n_1392)
);

NOR2x1_ASAP7_75t_L g1393 ( 
.A(n_1391),
.B(n_147),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1386),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1390),
.B(n_1139),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1388),
.B(n_1246),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1384),
.B(n_150),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1392),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1385),
.B(n_152),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1399),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1394),
.A2(n_1387),
.B(n_1389),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1397),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_SL g1403 ( 
.A(n_1398),
.B(n_1393),
.Y(n_1403)
);

OAI22x1_ASAP7_75t_L g1404 ( 
.A1(n_1395),
.A2(n_159),
.B1(n_162),
.B2(n_171),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1396),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1405),
.A2(n_1400),
.B1(n_1402),
.B2(n_1401),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1404),
.Y(n_1407)
);

AOI221xp5_ASAP7_75t_L g1408 ( 
.A1(n_1403),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.C(n_184),
.Y(n_1408)
);

AOI31xp33_ASAP7_75t_L g1409 ( 
.A1(n_1407),
.A2(n_189),
.A3(n_191),
.B(n_193),
.Y(n_1409)
);

AOI31xp33_ASAP7_75t_L g1410 ( 
.A1(n_1406),
.A2(n_194),
.A3(n_197),
.B(n_198),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1408),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_1411)
);

OAI322xp33_ASAP7_75t_L g1412 ( 
.A1(n_1411),
.A2(n_221),
.A3(n_225),
.B1(n_227),
.B2(n_228),
.C1(n_230),
.C2(n_231),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1410),
.B(n_235),
.Y(n_1413)
);

XNOR2xp5_ASAP7_75t_L g1414 ( 
.A(n_1409),
.B(n_237),
.Y(n_1414)
);

INVxp67_ASAP7_75t_SL g1415 ( 
.A(n_1413),
.Y(n_1415)
);

AOI21xp33_ASAP7_75t_L g1416 ( 
.A1(n_1414),
.A2(n_242),
.B(n_243),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1415),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1416),
.Y(n_1418)
);

AOI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1417),
.A2(n_1412),
.B1(n_244),
.B2(n_247),
.C(n_248),
.Y(n_1419)
);

AOI211xp5_ASAP7_75t_L g1420 ( 
.A1(n_1419),
.A2(n_1418),
.B(n_258),
.C(n_264),
.Y(n_1420)
);


endmodule