module real_aes_6073_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_929, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_929;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_884;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_922;
wire n_633;
wire n_926;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_0), .A2(n_208), .B1(n_464), .B2(n_466), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_1), .A2(n_123), .B1(n_495), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_2), .A2(n_98), .B1(n_415), .B2(n_417), .Y(n_414) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_3), .Y(n_668) );
AND2x4_ASAP7_75t_L g678 ( .A(n_3), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g687 ( .A(n_3), .B(n_239), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_4), .A2(n_200), .B1(n_363), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_5), .A2(n_116), .B1(n_690), .B2(n_712), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_6), .A2(n_54), .B1(n_394), .B2(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g530 ( .A(n_7), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_8), .A2(n_246), .B1(n_326), .B2(n_344), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_9), .A2(n_218), .B1(n_385), .B2(n_387), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_10), .A2(n_53), .B1(n_376), .B2(n_377), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g890 ( .A1(n_11), .A2(n_498), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_12), .A2(n_169), .B1(n_487), .B2(n_488), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_13), .A2(n_109), .B1(n_412), .B2(n_413), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_14), .A2(n_17), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_15), .A2(n_149), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_16), .A2(n_244), .B1(n_478), .B2(n_479), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_18), .A2(n_50), .B1(n_363), .B2(n_364), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_19), .Y(n_688) );
XNOR2x1_ASAP7_75t_L g433 ( .A(n_20), .B(n_434), .Y(n_433) );
INVxp33_ASAP7_75t_SL g705 ( .A(n_20), .Y(n_705) );
AO22x2_ASAP7_75t_L g744 ( .A1(n_21), .A2(n_61), .B1(n_690), .B2(n_712), .Y(n_744) );
AO22x1_ASAP7_75t_L g745 ( .A1(n_22), .A2(n_248), .B1(n_717), .B2(n_723), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_23), .A2(n_190), .B1(n_366), .B2(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_24), .B(n_390), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_25), .A2(n_127), .B1(n_412), .B2(n_541), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_26), .A2(n_243), .B1(n_381), .B2(n_383), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_27), .A2(n_60), .B1(n_370), .B2(n_417), .Y(n_584) );
INVx1_ASAP7_75t_L g443 ( .A(n_28), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_29), .A2(n_214), .B1(n_478), .B2(n_479), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_30), .A2(n_47), .B1(n_260), .B2(n_420), .C(n_422), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_31), .A2(n_65), .B1(n_302), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_32), .A2(n_178), .B1(n_370), .B2(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g423 ( .A(n_33), .Y(n_423) );
INVx1_ASAP7_75t_L g570 ( .A(n_34), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_35), .A2(n_111), .B1(n_686), .B2(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g281 ( .A(n_36), .Y(n_281) );
INVxp67_ASAP7_75t_L g297 ( .A(n_36), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_36), .B(n_185), .Y(n_320) );
OA22x2_ASAP7_75t_L g474 ( .A1(n_37), .A2(n_475), .B1(n_500), .B2(n_501), .Y(n_474) );
INVx1_ASAP7_75t_L g501 ( .A(n_37), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_38), .A2(n_187), .B1(n_495), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_39), .A2(n_119), .B1(n_394), .B2(n_439), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_40), .A2(n_192), .B1(n_680), .B2(n_690), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_41), .A2(n_113), .B1(n_717), .B2(n_719), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_42), .A2(n_131), .B1(n_499), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_43), .A2(n_51), .B1(n_481), .B2(n_482), .Y(n_895) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_44), .B(n_265), .Y(n_277) );
INVx1_ASAP7_75t_L g451 ( .A(n_45), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_46), .A2(n_155), .B1(n_366), .B2(n_368), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_48), .A2(n_69), .B1(n_364), .B2(n_471), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_49), .A2(n_238), .B1(n_285), .B2(n_289), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_52), .A2(n_197), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_55), .A2(n_211), .B1(n_712), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_56), .A2(n_232), .B1(n_376), .B2(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g666 ( .A(n_57), .Y(n_666) );
INVxp33_ASAP7_75t_SL g691 ( .A(n_58), .Y(n_691) );
INVx1_ASAP7_75t_L g677 ( .A(n_59), .Y(n_677) );
AND2x4_ASAP7_75t_L g683 ( .A(n_59), .B(n_666), .Y(n_683) );
INVx1_ASAP7_75t_SL g718 ( .A(n_59), .Y(n_718) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_62), .A2(n_247), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_63), .A2(n_86), .B1(n_495), .B2(n_496), .Y(n_564) );
INVx1_ASAP7_75t_L g314 ( .A(n_64), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_66), .A2(n_223), .B1(n_353), .B2(n_417), .Y(n_554) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_67), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_68), .A2(n_73), .B1(n_363), .B2(n_412), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_70), .B(n_569), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_71), .A2(n_242), .B1(n_326), .B2(n_332), .Y(n_325) );
INVx1_ASAP7_75t_L g437 ( .A(n_72), .Y(n_437) );
AOI21x1_ASAP7_75t_SL g525 ( .A1(n_74), .A2(n_526), .B(n_529), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_75), .A2(n_153), .B1(n_387), .B2(n_427), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_76), .A2(n_213), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_77), .A2(n_108), .B1(n_431), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g269 ( .A(n_78), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_78), .B(n_184), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_79), .A2(n_104), .B1(n_484), .B2(n_487), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_80), .A2(n_130), .B1(n_394), .B2(n_396), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_81), .A2(n_160), .B1(n_370), .B2(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_82), .A2(n_180), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_83), .A2(n_145), .B1(n_549), .B2(n_550), .C(n_552), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_84), .B(n_260), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_85), .A2(n_138), .B1(n_491), .B2(n_499), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_87), .A2(n_139), .B1(n_690), .B2(n_712), .Y(n_720) );
AO221x2_ASAP7_75t_L g672 ( .A1(n_88), .A2(n_90), .B1(n_673), .B2(n_680), .C(n_684), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_89), .A2(n_240), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_91), .A2(n_122), .B1(n_300), .B2(n_302), .Y(n_299) );
AOI221xp5_ASAP7_75t_SL g489 ( .A1(n_92), .A2(n_221), .B1(n_490), .B2(n_491), .C(n_492), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_93), .A2(n_146), .B1(n_341), .B2(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_94), .B(n_311), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_95), .A2(n_245), .B1(n_675), .B2(n_712), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_96), .A2(n_210), .B1(n_410), .B2(n_469), .Y(n_583) );
INVx1_ASAP7_75t_L g923 ( .A(n_97), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g921 ( .A1(n_99), .A2(n_491), .B(n_922), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_100), .A2(n_236), .B1(n_484), .B2(n_485), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_101), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_102), .A2(n_165), .B1(n_495), .B2(n_496), .C(n_497), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_103), .A2(n_215), .B1(n_479), .B2(n_484), .Y(n_896) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_105), .A2(n_311), .B(n_313), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_106), .A2(n_212), .B1(n_366), .B2(n_368), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_107), .A2(n_162), .B1(n_609), .B2(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g619 ( .A(n_110), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_112), .B(n_490), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_114), .A2(n_166), .B1(n_391), .B2(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g915 ( .A1(n_115), .A2(n_174), .B1(n_487), .B2(n_488), .Y(n_915) );
INVx1_ASAP7_75t_L g578 ( .A(n_116), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_117), .A2(n_148), .B1(n_487), .B2(n_488), .Y(n_486) );
NAND2xp33_ASAP7_75t_L g638 ( .A(n_118), .B(n_326), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_120), .A2(n_140), .B1(n_481), .B2(n_482), .Y(n_913) );
INVx1_ASAP7_75t_L g892 ( .A(n_121), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_124), .A2(n_179), .B1(n_455), .B2(n_456), .Y(n_454) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_125), .A2(n_616), .B(n_618), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_126), .A2(n_176), .B1(n_429), .B2(n_431), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_128), .A2(n_189), .B1(n_717), .B2(n_719), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_129), .A2(n_161), .B1(n_336), .B2(n_341), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_132), .A2(n_230), .B1(n_478), .B2(n_491), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_133), .A2(n_216), .B1(n_364), .B2(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g533 ( .A(n_134), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_135), .A2(n_194), .B1(n_495), .B2(n_499), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_136), .A2(n_159), .B1(n_601), .B2(n_604), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_137), .A2(n_141), .B1(n_364), .B2(n_368), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_142), .A2(n_883), .B1(n_884), .B2(n_898), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_142), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_143), .A2(n_235), .B1(n_351), .B2(n_353), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_144), .A2(n_224), .B1(n_412), .B2(n_413), .Y(n_542) );
AO22x1_ASAP7_75t_L g497 ( .A1(n_147), .A2(n_206), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22x1_ASAP7_75t_L g596 ( .A1(n_150), .A2(n_597), .B1(n_598), .B2(n_631), .Y(n_596) );
INVx1_ASAP7_75t_L g631 ( .A(n_150), .Y(n_631) );
OAI22x1_ASAP7_75t_L g659 ( .A1(n_150), .A2(n_597), .B1(n_598), .B2(n_631), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_151), .A2(n_220), .B1(n_485), .B2(n_488), .Y(n_558) );
INVx1_ASAP7_75t_L g440 ( .A(n_152), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_154), .A2(n_237), .B1(n_344), .B2(n_348), .Y(n_343) );
XNOR2x1_ASAP7_75t_L g256 ( .A(n_156), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_157), .B(n_456), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_158), .A2(n_181), .B1(n_675), .B2(n_686), .Y(n_751) );
INVx1_ASAP7_75t_L g589 ( .A(n_163), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_164), .A2(n_196), .B1(n_485), .B2(n_496), .Y(n_887) );
OA22x2_ASAP7_75t_L g263 ( .A1(n_167), .A2(n_185), .B1(n_264), .B2(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g308 ( .A(n_167), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_168), .A2(n_182), .B1(n_351), .B2(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_170), .A2(n_201), .B1(n_445), .B2(n_587), .C(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g567 ( .A(n_171), .Y(n_567) );
XNOR2x1_ASAP7_75t_L g510 ( .A(n_172), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_173), .A2(n_225), .B1(n_368), .B2(n_410), .Y(n_409) );
AOI221x1_ASAP7_75t_L g639 ( .A1(n_175), .A2(n_222), .B1(n_344), .B2(n_353), .C(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g700 ( .A(n_177), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_183), .A2(n_191), .B1(n_675), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g283 ( .A(n_184), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_184), .B(n_306), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g309 ( .A1(n_185), .A2(n_198), .B(n_298), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_186), .A2(n_203), .B1(n_498), .B2(n_499), .Y(n_920) );
AND2x2_ASAP7_75t_L g640 ( .A(n_188), .B(n_342), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_189), .A2(n_904), .B1(n_907), .B2(n_924), .Y(n_903) );
XNOR2x2_ASAP7_75t_SL g909 ( .A(n_189), .B(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_193), .A2(n_207), .B1(n_387), .B2(n_532), .Y(n_593) );
INVx1_ASAP7_75t_SL g701 ( .A(n_195), .Y(n_701) );
INVx1_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_198), .B(n_233), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_199), .A2(n_229), .B1(n_481), .B2(n_482), .Y(n_561) );
INVx1_ASAP7_75t_L g553 ( .A(n_202), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_204), .B(n_645), .Y(n_644) );
XNOR2x1_ASAP7_75t_L g537 ( .A(n_205), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_209), .A2(n_219), .B1(n_623), .B2(n_625), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_217), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_226), .B(n_637), .C(n_641), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_226), .A2(n_641), .B1(n_647), .B2(n_929), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_226), .A2(n_637), .B(n_652), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_227), .A2(n_241), .B1(n_383), .B2(n_427), .Y(n_594) );
INVx1_ASAP7_75t_L g447 ( .A(n_228), .Y(n_447) );
INVx1_ASAP7_75t_L g358 ( .A(n_231), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_233), .B(n_276), .Y(n_275) );
AOI21xp33_ASAP7_75t_L g565 ( .A1(n_234), .A2(n_491), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g679 ( .A(n_239), .Y(n_679) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_239), .Y(n_926) );
XNOR2x1_ASAP7_75t_L g404 ( .A(n_245), .B(n_405), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_660), .B(n_669), .Y(n_249) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_503), .Y(n_250) );
XNOR2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_400), .Y(n_251) );
AOI22x1_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B1(n_355), .B2(n_398), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_258), .B(n_324), .Y(n_257) );
NAND4xp25_ASAP7_75t_L g258 ( .A(n_259), .B(n_284), .C(n_299), .D(n_310), .Y(n_258) );
BUFx8_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g382 ( .A(n_261), .Y(n_382) );
INVx2_ASAP7_75t_L g446 ( .A(n_261), .Y(n_446) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_261), .Y(n_490) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_261), .Y(n_624) );
BUFx3_ASAP7_75t_L g645 ( .A(n_261), .Y(n_645) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_272), .Y(n_261) );
AND2x4_ASAP7_75t_L g301 ( .A(n_262), .B(n_287), .Y(n_301) );
AND2x4_ASAP7_75t_L g491 ( .A(n_262), .B(n_287), .Y(n_491) );
AND2x2_ASAP7_75t_L g569 ( .A(n_262), .B(n_272), .Y(n_569) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
AND2x2_ASAP7_75t_L g288 ( .A(n_263), .B(n_267), .Y(n_288) );
AND2x2_ASAP7_75t_L g295 ( .A(n_263), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g347 ( .A(n_263), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_264), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp33_ASAP7_75t_L g268 ( .A(n_265), .B(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g276 ( .A(n_265), .Y(n_276) );
NAND2xp33_ASAP7_75t_L g282 ( .A(n_265), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
AND2x4_ASAP7_75t_L g346 ( .A(n_266), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_269), .B(n_308), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_271), .A2(n_297), .B(n_298), .Y(n_296) );
AND2x4_ASAP7_75t_L g303 ( .A(n_272), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g312 ( .A(n_272), .B(n_288), .Y(n_312) );
AND2x2_ASAP7_75t_L g352 ( .A(n_272), .B(n_346), .Y(n_352) );
AND2x4_ASAP7_75t_L g482 ( .A(n_272), .B(n_346), .Y(n_482) );
AND2x2_ASAP7_75t_L g498 ( .A(n_272), .B(n_288), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_272), .B(n_304), .Y(n_499) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g287 ( .A(n_274), .B(n_278), .Y(n_287) );
AND2x2_ASAP7_75t_L g291 ( .A(n_274), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g330 ( .A(n_274), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g339 ( .A(n_274), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_276), .B(n_281), .Y(n_280) );
INVxp67_ASAP7_75t_L g306 ( .A(n_276), .Y(n_306) );
NAND3xp33_ASAP7_75t_L g322 ( .A(n_277), .B(n_305), .C(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g388 ( .A(n_286), .Y(n_388) );
BUFx3_ASAP7_75t_L g630 ( .A(n_286), .Y(n_630) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x4_ASAP7_75t_L g354 ( .A(n_287), .B(n_346), .Y(n_354) );
AND2x4_ASAP7_75t_L g481 ( .A(n_287), .B(n_346), .Y(n_481) );
AND2x4_ASAP7_75t_L g495 ( .A(n_287), .B(n_288), .Y(n_495) );
AND2x4_ASAP7_75t_L g333 ( .A(n_288), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g342 ( .A(n_288), .B(n_339), .Y(n_342) );
AND2x2_ASAP7_75t_L g367 ( .A(n_288), .B(n_339), .Y(n_367) );
AND2x4_ASAP7_75t_L g478 ( .A(n_288), .B(n_339), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_288), .B(n_329), .Y(n_479) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx5_ASAP7_75t_L g395 ( .A(n_290), .Y(n_395) );
BUFx4f_ASAP7_75t_L g455 ( .A(n_290), .Y(n_455) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
AND2x2_ASAP7_75t_L g496 ( .A(n_291), .B(n_295), .Y(n_496) );
AND2x4_ASAP7_75t_L g918 ( .A(n_291), .B(n_295), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
BUFx2_ASAP7_75t_L g627 ( .A(n_300), .Y(n_627) );
BUFx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g386 ( .A(n_301), .Y(n_386) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_301), .Y(n_427) );
BUFx3_ASAP7_75t_L g439 ( .A(n_301), .Y(n_439) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_303), .Y(n_383) );
INVx3_ASAP7_75t_L g432 ( .A(n_303), .Y(n_432) );
AND2x4_ASAP7_75t_L g328 ( .A(n_304), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g338 ( .A(n_304), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g487 ( .A(n_304), .B(n_339), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_304), .B(n_329), .Y(n_488) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_309), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
BUFx3_ASAP7_75t_L g617 ( .A(n_311), .Y(n_617) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g392 ( .A(n_312), .Y(n_392) );
INVx3_ASAP7_75t_L g421 ( .A(n_312), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_315), .B(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g396 ( .A(n_316), .Y(n_396) );
INVx2_ASAP7_75t_L g425 ( .A(n_316), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_316), .B(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_316), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_316), .B(n_923), .Y(n_922) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx3_ASAP7_75t_L g458 ( .A(n_317), .Y(n_458) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B(n_322), .Y(n_317) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_319), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_325), .B(n_335), .C(n_343), .D(n_350), .Y(n_324) );
INVx5_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g408 ( .A(n_327), .Y(n_408) );
INVx6_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx12f_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
AND2x4_ASAP7_75t_L g345 ( .A(n_329), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g334 ( .A(n_330), .Y(n_334) );
INVx1_ASAP7_75t_L g340 ( .A(n_331), .Y(n_340) );
BUFx3_ASAP7_75t_L g607 ( .A(n_332), .Y(n_607) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_333), .Y(n_368) );
BUFx3_ASAP7_75t_L g462 ( .A(n_333), .Y(n_462) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_333), .Y(n_541) );
AND2x4_ASAP7_75t_L g485 ( .A(n_334), .B(n_346), .Y(n_485) );
BUFx2_ASAP7_75t_SL g613 ( .A(n_336), .Y(n_613) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx4_ASAP7_75t_L g377 ( .A(n_337), .Y(n_377) );
INVx2_ASAP7_75t_SL g413 ( .A(n_337), .Y(n_413) );
INVx4_ASAP7_75t_L g469 ( .A(n_337), .Y(n_469) );
INVx1_ASAP7_75t_L g515 ( .A(n_337), .Y(n_515) );
INVx4_ASAP7_75t_L g654 ( .A(n_337), .Y(n_654) );
INVx8_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g349 ( .A(n_339), .B(n_346), .Y(n_349) );
AND2x4_ASAP7_75t_L g484 ( .A(n_339), .B(n_346), .Y(n_484) );
BUFx4f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_342), .Y(n_606) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_345), .Y(n_363) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_345), .Y(n_471) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_345), .Y(n_603) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g374 ( .A(n_352), .Y(n_374) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
BUFx5_ASAP7_75t_L g520 ( .A(n_352), .Y(n_520) );
BUFx12f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_354), .Y(n_370) );
INVx3_ASAP7_75t_L g416 ( .A(n_354), .Y(n_416) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g399 ( .A(n_357), .Y(n_399) );
AO21x2_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B(n_397), .Y(n_357) );
NOR3xp33_ASAP7_75t_SL g397 ( .A(n_358), .B(n_361), .C(n_379), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_378), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND4xp25_ASAP7_75t_SL g361 ( .A(n_362), .B(n_365), .C(n_369), .D(n_375), .Y(n_361) );
BUFx3_ASAP7_75t_L g604 ( .A(n_364), .Y(n_604) );
BUFx8_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_373), .Y(n_466) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND4xp25_ASAP7_75t_L g379 ( .A(n_380), .B(n_384), .C(n_389), .D(n_393), .Y(n_379) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g549 ( .A(n_382), .Y(n_549) );
BUFx3_ASAP7_75t_L g625 ( .A(n_383), .Y(n_625) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g441 ( .A(n_387), .Y(n_441) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
INVx2_ASAP7_75t_L g643 ( .A(n_388), .Y(n_643) );
BUFx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_392), .Y(n_528) );
INVx4_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g532 ( .A(n_395), .Y(n_532) );
INVx2_ASAP7_75t_L g544 ( .A(n_395), .Y(n_544) );
INVx2_ASAP7_75t_SL g534 ( .A(n_396), .Y(n_534) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_472), .B2(n_502), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_433), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_418), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .C(n_411), .D(n_414), .Y(n_406) );
BUFx12f_ASAP7_75t_L g514 ( .A(n_412), .Y(n_514) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_412), .Y(n_612) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g465 ( .A(n_416), .Y(n_465) );
INVx1_ASAP7_75t_L g609 ( .A(n_416), .Y(n_609) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_417), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_426), .C(n_428), .Y(n_418) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g453 ( .A(n_421), .Y(n_453) );
INVx3_ASAP7_75t_SL g587 ( .A(n_421), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_459), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_442), .C(n_450), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g524 ( .A(n_446), .Y(n_524) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g620 ( .A(n_455), .Y(n_620) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_457), .B(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx4_ASAP7_75t_L g592 ( .A(n_458), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
BUFx4f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_SL g502 ( .A(n_472), .Y(n_502) );
BUFx4_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g500 ( .A(n_475), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_489), .C(n_494), .Y(n_475) );
AND4x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .C(n_483), .D(n_486), .Y(n_476) );
INVx2_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
XNOR2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_573), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI22xp33_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_507), .B1(n_535), .B2(n_536), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND4xp75_ASAP7_75t_SL g511 ( .A(n_512), .B(n_517), .C(n_521), .D(n_525), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_533), .B2(n_534), .Y(n_529) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OA22x2_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_555), .B1(n_571), .B2(n_572), .Y(n_536) );
INVx1_ASAP7_75t_L g571 ( .A(n_537), .Y(n_571) );
NOR2x1_ASAP7_75t_L g538 ( .A(n_539), .B(n_546), .Y(n_538) );
NAND4xp25_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .C(n_543), .D(n_545), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .C(n_554), .Y(n_546) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g572 ( .A(n_555), .Y(n_572) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_570), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .C(n_560), .D(n_561), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .C(n_565), .D(n_568), .Y(n_562) );
XOR2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_595), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
XNOR2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
NAND4xp25_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .C(n_583), .D(n_584), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_593), .C(n_594), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_592), .B(n_892), .Y(n_891) );
OA22x2_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_632), .B1(n_633), .B2(n_659), .Y(n_595) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_614), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g599 ( .A(n_600), .B(n_605), .C(n_608), .D(n_611), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_622), .C(n_626), .Y(n_614) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_621), .Y(n_618) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AO21x2_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_646), .B(n_656), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_642), .B(n_644), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_652), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2x1_ASAP7_75t_SL g652 ( .A(n_653), .B(n_655), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
BUFx10_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .C(n_668), .Y(n_663) );
AND2x2_ASAP7_75t_L g901 ( .A(n_664), .B(n_902), .Y(n_901) );
AND2x2_ASAP7_75t_L g905 ( .A(n_664), .B(n_906), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_664), .A2(n_668), .B(n_718), .Y(n_927) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AO21x1_ASAP7_75t_L g925 ( .A1(n_665), .A2(n_926), .B(n_927), .Y(n_925) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g676 ( .A(n_666), .B(n_677), .Y(n_676) );
AND3x4_ASAP7_75t_L g717 ( .A(n_666), .B(n_678), .C(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_667), .B(n_902), .Y(n_906) );
INVx1_ASAP7_75t_L g902 ( .A(n_668), .Y(n_902) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_880), .B1(n_882), .B2(n_899), .C(n_903), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_692), .B(n_799), .C(n_850), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_671), .A2(n_800), .B(n_832), .Y(n_799) );
INVx1_ASAP7_75t_L g868 ( .A(n_671), .Y(n_868) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI311xp33_ASAP7_75t_L g832 ( .A1(n_672), .A2(n_833), .A3(n_841), .B(n_843), .C(n_846), .Y(n_832) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_673), .Y(n_881) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_674), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
INVx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
AND2x4_ASAP7_75t_L g686 ( .A(n_676), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g719 ( .A(n_676), .B(n_687), .Y(n_719) );
AND2x2_ASAP7_75t_L g723 ( .A(n_676), .B(n_687), .Y(n_723) );
AND2x4_ASAP7_75t_L g682 ( .A(n_678), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_678), .B(n_683), .Y(n_704) );
AND2x4_ASAP7_75t_L g712 ( .A(n_678), .B(n_683), .Y(n_712) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g690 ( .A(n_683), .B(n_687), .Y(n_690) );
AND2x2_ASAP7_75t_L g710 ( .A(n_683), .B(n_687), .Y(n_710) );
AND2x2_ASAP7_75t_L g728 ( .A(n_683), .B(n_687), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_685), .A2(n_689), .B1(n_700), .B2(n_701), .Y(n_699) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND5xp2_ASAP7_75t_L g692 ( .A(n_693), .B(n_730), .C(n_739), .D(n_771), .E(n_792), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_725), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_706), .Y(n_696) );
AND2x2_ASAP7_75t_L g740 ( .A(n_697), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g758 ( .A(n_697), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_697), .B(n_708), .Y(n_775) );
AND2x2_ASAP7_75t_L g865 ( .A(n_697), .B(n_759), .Y(n_865) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_698), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g767 ( .A(n_698), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_698), .B(n_738), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_698), .B(n_726), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_698), .B(n_743), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_698), .B(n_770), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_698), .B(n_707), .Y(n_825) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_698), .Y(n_844) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g766 ( .A1(n_706), .A2(n_752), .B(n_767), .C(n_768), .Y(n_766) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_713), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_707), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_707), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g777 ( .A(n_707), .B(n_778), .Y(n_777) );
OR2x2_ASAP7_75t_L g788 ( .A(n_707), .B(n_735), .Y(n_788) );
OR2x2_ASAP7_75t_L g812 ( .A(n_707), .B(n_714), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_707), .B(n_721), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_707), .B(n_735), .Y(n_857) );
INVx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g764 ( .A(n_708), .B(n_721), .Y(n_764) );
INVx1_ASAP7_75t_L g782 ( .A(n_708), .Y(n_782) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_714), .B(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_721), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_715), .Y(n_735) );
AND2x2_ASAP7_75t_L g778 ( .A(n_715), .B(n_721), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_715), .A2(n_803), .B1(n_805), .B2(n_807), .Y(n_802) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_720), .Y(n_715) );
OR2x2_ASAP7_75t_L g734 ( .A(n_721), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g752 ( .A(n_721), .Y(n_752) );
AND2x2_ASAP7_75t_L g759 ( .A(n_721), .B(n_735), .Y(n_759) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_726), .Y(n_738) );
OR2x2_ASAP7_75t_L g742 ( .A(n_726), .B(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g762 ( .A(n_726), .Y(n_762) );
AND2x2_ASAP7_75t_L g770 ( .A(n_726), .B(n_743), .Y(n_770) );
AND2x4_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_736), .Y(n_731) );
INVx1_ASAP7_75t_L g876 ( .A(n_732), .Y(n_876) );
INVx1_ASAP7_75t_L g755 ( .A(n_734), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_734), .B(n_825), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_735), .B(n_781), .Y(n_780) );
OAI222xp33_ASAP7_75t_L g772 ( .A1(n_736), .A2(n_768), .B1(n_773), .B2(n_776), .C1(n_779), .C2(n_783), .Y(n_772) );
OAI211xp5_ASAP7_75t_L g833 ( .A1(n_736), .A2(n_834), .B(n_836), .C(n_839), .Y(n_833) );
AND2x2_ASAP7_75t_L g872 ( .A(n_736), .B(n_748), .Y(n_872) );
AND3x1_ASAP7_75t_L g877 ( .A(n_736), .B(n_781), .C(n_865), .Y(n_877) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g822 ( .A(n_737), .Y(n_822) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g791 ( .A(n_738), .B(n_743), .Y(n_791) );
AOI311xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_746), .A3(n_752), .B(n_753), .C(n_763), .Y(n_739) );
AOI222xp33_ASAP7_75t_L g792 ( .A1(n_741), .A2(n_743), .B1(n_759), .B2(n_793), .C1(n_795), .C2(n_796), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_741), .A2(n_814), .B1(n_817), .B2(n_818), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_741), .A2(n_863), .B1(n_866), .B2(n_869), .C(n_873), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_741), .B(n_823), .Y(n_874) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g765 ( .A(n_742), .B(n_749), .Y(n_765) );
INVx1_ASAP7_75t_L g786 ( .A(n_743), .Y(n_786) );
CKINVDCx6p67_ASAP7_75t_R g809 ( .A(n_743), .Y(n_809) );
OR2x2_ASAP7_75t_L g842 ( .A(n_743), .B(n_748), .Y(n_842) );
OR2x6_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_746), .B(n_791), .Y(n_811) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g771 ( .A1(n_747), .A2(n_772), .B1(n_781), .B2(n_784), .C1(n_787), .C2(n_789), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_747), .B(n_791), .Y(n_790) );
INVx5_ASAP7_75t_L g801 ( .A(n_747), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_747), .B(n_767), .Y(n_861) );
INVx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g761 ( .A(n_748), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g827 ( .A(n_748), .B(n_785), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_748), .B(n_809), .Y(n_849) );
INVx3_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g784 ( .A(n_749), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g845 ( .A(n_749), .B(n_769), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_752), .B(n_774), .Y(n_773) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B(n_760), .Y(n_753) );
INVx1_ASAP7_75t_L g854 ( .A(n_754), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_755), .B(n_774), .Y(n_815) );
O2A1O1Ixp33_ASAP7_75t_L g843 ( .A1(n_756), .A2(n_779), .B(n_844), .C(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g848 ( .A(n_757), .B(n_781), .Y(n_848) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_758), .B(n_787), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_758), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g817 ( .A(n_759), .B(n_781), .Y(n_817) );
AND2x2_ASAP7_75t_L g823 ( .A(n_759), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g858 ( .A(n_759), .Y(n_858) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g808 ( .A(n_762), .B(n_809), .Y(n_808) );
OAI21xp5_ASAP7_75t_SL g763 ( .A1(n_764), .A2(n_765), .B(n_766), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_SL g846 ( .A1(n_764), .A2(n_837), .B(n_847), .C(n_849), .Y(n_846) );
INVx1_ASAP7_75t_L g855 ( .A(n_765), .Y(n_855) );
AND2x2_ASAP7_75t_L g795 ( .A(n_767), .B(n_778), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g807 ( .A(n_767), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g837 ( .A(n_767), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_767), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_769), .B(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_777), .A2(n_818), .B(n_827), .Y(n_831) );
INVx1_ASAP7_75t_L g804 ( .A(n_778), .Y(n_804) );
AND2x2_ASAP7_75t_L g840 ( .A(n_778), .B(n_781), .Y(n_840) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_781), .B(n_865), .Y(n_864) );
INVx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_783), .A2(n_811), .B(n_812), .C(n_813), .Y(n_810) );
AOI211xp5_ASAP7_75t_L g851 ( .A1(n_784), .A2(n_793), .B(n_852), .C(n_856), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_785), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g878 ( .A1(n_788), .A2(n_790), .B(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_791), .A2(n_828), .B(n_840), .Y(n_879) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI211xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B(n_810), .C(n_820), .Y(n_800) );
O2A1O1Ixp33_ASAP7_75t_L g875 ( .A1(n_801), .A2(n_876), .B(n_877), .C(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g870 ( .A(n_808), .Y(n_870) );
INVx1_ASAP7_75t_L g838 ( .A(n_812), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND3xp33_ASAP7_75t_SL g820 ( .A(n_821), .B(n_826), .C(n_831), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g867 ( .A(n_837), .B(n_840), .C(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND3xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_862), .C(n_875), .Y(n_850) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
AOI21xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B(n_859), .Y(n_856) );
INVxp67_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NOR2x1_ASAP7_75t_L g885 ( .A(n_886), .B(n_893), .Y(n_885) );
NAND4xp25_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .C(n_889), .D(n_890), .Y(n_886) );
NAND4xp25_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .C(n_896), .D(n_897), .Y(n_893) );
INVx1_ASAP7_75t_SL g899 ( .A(n_900), .Y(n_899) );
BUFx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx3_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OR2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_916), .Y(n_910) );
NAND4xp25_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .C(n_914), .D(n_915), .Y(n_911) );
NAND4xp25_ASAP7_75t_L g916 ( .A(n_917), .B(n_919), .C(n_920), .D(n_921), .Y(n_916) );
BUFx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
endmodule