module fake_netlist_6_4015_n_1625 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1625);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1625;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_33),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_100),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_58),
.Y(n_150)
);

INVxp33_ASAP7_75t_R g151 ( 
.A(n_82),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_4),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_53),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_94),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_63),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_87),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_93),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_103),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_14),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_4),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_111),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

BUFx8_ASAP7_75t_SL g170 ( 
.A(n_76),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_57),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_112),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_32),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_18),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_32),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_27),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_84),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_67),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_25),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_40),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_116),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_85),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_51),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_109),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_31),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_96),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_80),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_2),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_3),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_51),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_31),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_72),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_77),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_70),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_25),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_88),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_124),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_26),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_46),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_22),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_108),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_46),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_2),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_75),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_60),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_101),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_41),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_52),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_55),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_35),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_98),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_126),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_132),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_65),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_14),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_3),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_92),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_102),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_39),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_29),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_97),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_68),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_66),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_86),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_37),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_45),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_107),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_83),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_71),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_11),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_11),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_136),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_50),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_22),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_44),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_143),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_105),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_79),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_27),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_10),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_47),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_117),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_28),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_0),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_174),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_170),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_174),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_148),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_268),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_174),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_237),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_149),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_199),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_174),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_155),
.B(n_1),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_195),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_216),
.B(n_1),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_152),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_216),
.B(n_6),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_160),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_169),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_171),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_262),
.B(n_7),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_172),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_9),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_147),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_147),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_183),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_178),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_178),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_184),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_150),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_186),
.B(n_10),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_186),
.B(n_12),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_190),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_205),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_276),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_191),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_205),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_196),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_221),
.Y(n_336)
);

BUFx2_ASAP7_75t_SL g337 ( 
.A(n_150),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_161),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_257),
.B(n_12),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_200),
.Y(n_340)
);

BUFx6f_ASAP7_75t_SL g341 ( 
.A(n_181),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_159),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_221),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_206),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_209),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_153),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_215),
.B(n_15),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_154),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_167),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_211),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_175),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_176),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_202),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_203),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_215),
.B(n_19),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_173),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_213),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_223),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_182),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_159),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_227),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_257),
.B(n_20),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_236),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_243),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_163),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_290),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_158),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_295),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_291),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_287),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_289),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_307),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_164),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_311),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_314),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_292),
.B(n_220),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_318),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_201),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_298),
.A2(n_286),
.B1(n_192),
.B2(n_166),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_293),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_293),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_289),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_301),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_322),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_261),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_297),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_303),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_305),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_305),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_306),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_310),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_330),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_310),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_312),
.B(n_220),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_312),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_335),
.B(n_235),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_319),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_327),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_340),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_315),
.B(n_185),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_345),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_168),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_321),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_346),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_300),
.B(n_193),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_271),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_212),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_294),
.B(n_163),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_321),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_R g428 ( 
.A(n_358),
.B(n_189),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_324),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_342),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_362),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_367),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_294),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_296),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_288),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_341),
.B(n_165),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_420),
.B(n_235),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_410),
.B(n_244),
.Y(n_440)
);

INVx4_ASAP7_75t_SL g441 ( 
.A(n_423),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_299),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_370),
.B(n_304),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_428),
.A2(n_274),
.B1(n_165),
.B2(n_259),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_377),
.B(n_370),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_392),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_385),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_313),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_369),
.B(n_244),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_259),
.B1(n_274),
.B2(n_208),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_371),
.B(n_255),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_385),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_388),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_384),
.B(n_329),
.C(n_328),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_337),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_341),
.Y(n_461)
);

BUFx4f_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_374),
.B(n_341),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_372),
.B(n_337),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_376),
.B(n_255),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_378),
.B(n_336),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_386),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_424),
.B(n_343),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_382),
.Y(n_474)
);

NOR2x1p5_ASAP7_75t_L g475 ( 
.A(n_379),
.B(n_343),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_381),
.B(n_344),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_193),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_408),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_390),
.A2(n_364),
.B1(n_339),
.B2(n_349),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_368),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_417),
.A2(n_258),
.B1(n_208),
.B2(n_357),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_401),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_408),
.B(n_193),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_405),
.B(n_193),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_411),
.B(n_258),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_384),
.B(n_344),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_347),
.Y(n_491)
);

CKINVDCx11_ASAP7_75t_R g492 ( 
.A(n_434),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_412),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_386),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_214),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_373),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_373),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g501 ( 
.A(n_438),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_413),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_423),
.B(n_375),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_387),
.B(n_224),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_432),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

INVx4_ASAP7_75t_SL g510 ( 
.A(n_386),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_419),
.B(n_347),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_422),
.B(n_348),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_430),
.B(n_366),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_429),
.B(n_193),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_429),
.B(n_198),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_386),
.Y(n_516)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_393),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_429),
.B(n_198),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_429),
.B(n_198),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_394),
.B(n_198),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_394),
.B(n_396),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

OR2x2_ASAP7_75t_SL g524 ( 
.A(n_437),
.B(n_151),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_397),
.B(n_350),
.Y(n_525)
);

BUFx8_ASAP7_75t_SL g526 ( 
.A(n_433),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_430),
.B(n_350),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g531 ( 
.A(n_430),
.B(n_281),
.C(n_280),
.Y(n_531)
);

BUFx4f_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_402),
.A2(n_284),
.B1(n_162),
.B2(n_157),
.Y(n_533)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_402),
.B(n_198),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_404),
.B(n_230),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_429),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_404),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_407),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_407),
.B(n_146),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_414),
.B(n_239),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_430),
.A2(n_366),
.B1(n_365),
.B2(n_363),
.Y(n_541)
);

AND3x2_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_156),
.C(n_177),
.Y(n_542)
);

BUFx8_ASAP7_75t_SL g543 ( 
.A(n_416),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_418),
.A2(n_233),
.B1(n_232),
.B2(n_234),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_386),
.B(n_218),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_398),
.B(n_353),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_421),
.A2(n_365),
.B1(n_363),
.B2(n_360),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_409),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_398),
.B(n_353),
.Y(n_551)
);

OAI22x1_ASAP7_75t_L g552 ( 
.A1(n_398),
.A2(n_250),
.B1(n_194),
.B2(n_204),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_427),
.B(n_240),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_427),
.B(n_241),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_427),
.A2(n_360),
.B1(n_359),
.B2(n_356),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_409),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_391),
.B(n_359),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_409),
.B(n_242),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_391),
.B(n_246),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_391),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_409),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_391),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_409),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_391),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_372),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_372),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_380),
.Y(n_567)
);

INVxp33_ASAP7_75t_SL g568 ( 
.A(n_438),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_420),
.B(n_218),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_385),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_443),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_512),
.B(n_181),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_478),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_442),
.B(n_252),
.Y(n_574)
);

BUFx4_ASAP7_75t_L g575 ( 
.A(n_526),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_442),
.B(n_181),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_481),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_481),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_447),
.B(n_179),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_448),
.B(n_254),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_458),
.A2(n_146),
.B1(n_166),
.B2(n_192),
.Y(n_582)
);

CKINVDCx8_ASAP7_75t_R g583 ( 
.A(n_486),
.Y(n_583)
);

AND2x4_ASAP7_75t_SL g584 ( 
.A(n_443),
.B(n_187),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_447),
.A2(n_264),
.B1(n_263),
.B2(n_265),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_459),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_462),
.B(n_218),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_444),
.B(n_229),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_468),
.B(n_283),
.C(n_267),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_450),
.B(n_188),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_467),
.B(n_197),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_491),
.B(n_207),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_449),
.B(n_210),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_439),
.A2(n_277),
.B1(n_247),
.B2(n_231),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_507),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_454),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_469),
.B(n_249),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_566),
.B(n_354),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_476),
.B(n_270),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_217),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_503),
.B(n_464),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_452),
.B(n_219),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_460),
.B(n_570),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_466),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_462),
.A2(n_218),
.B(n_278),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_460),
.B(n_278),
.Y(n_609)
);

AND2x6_ASAP7_75t_SL g610 ( 
.A(n_461),
.B(n_356),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_480),
.B(n_278),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_570),
.B(n_278),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_439),
.A2(n_228),
.B1(n_279),
.B2(n_238),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_452),
.B(n_222),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_567),
.A2(n_355),
.B(n_354),
.C(n_334),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_528),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_455),
.B(n_229),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_484),
.B(n_229),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_455),
.B(n_225),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_499),
.B(n_229),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_500),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_229),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_490),
.B(n_325),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_457),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_465),
.B(n_245),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_509),
.B(n_229),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_569),
.A2(n_228),
.B1(n_286),
.B2(n_238),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_473),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_548),
.A2(n_331),
.B(n_285),
.C(n_226),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_465),
.B(n_275),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_485),
.A2(n_279),
.B1(n_253),
.B2(n_272),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_488),
.B(n_273),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_457),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_488),
.B(n_251),
.Y(n_635)
);

AO221x1_ASAP7_75t_L g636 ( 
.A1(n_552),
.A2(n_533),
.B1(n_544),
.B2(n_530),
.C(n_529),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_538),
.B(n_266),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_456),
.B(n_505),
.Y(n_638)
);

NAND2x1_ASAP7_75t_L g639 ( 
.A(n_471),
.B(n_61),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_547),
.Y(n_640)
);

INVx8_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_440),
.B(n_62),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_440),
.B(n_187),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_475),
.B(n_272),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_557),
.B(n_59),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_479),
.Y(n_646)
);

AND2x6_ASAP7_75t_SL g647 ( 
.A(n_463),
.B(n_260),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_473),
.B(n_256),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_479),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_568),
.A2(n_260),
.B1(n_253),
.B2(n_256),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_483),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_506),
.B(n_187),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_463),
.B(n_539),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_513),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_565),
.B(n_20),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_446),
.B(n_21),
.Y(n_656)
);

AND2x4_ASAP7_75t_SL g657 ( 
.A(n_453),
.B(n_54),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_535),
.B(n_21),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_551),
.B(n_56),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_540),
.B(n_144),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_441),
.B(n_137),
.Y(n_661)
);

BUFx8_ASAP7_75t_L g662 ( 
.A(n_492),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_483),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_548),
.B(n_133),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_493),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_553),
.B(n_130),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_542),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_R g668 ( 
.A(n_474),
.B(n_95),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_501),
.B(n_23),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_501),
.B(n_24),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_554),
.B(n_129),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_496),
.B(n_24),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_521),
.B(n_122),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_527),
.B(n_26),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_508),
.B(n_28),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_556),
.B(n_89),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_495),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_558),
.B(n_81),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_527),
.B(n_74),
.Y(n_679)
);

AO22x1_ASAP7_75t_L g680 ( 
.A1(n_531),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_541),
.B(n_36),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_555),
.B(n_37),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_523),
.B(n_69),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_555),
.B(n_49),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_498),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_502),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_525),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_533),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_533),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_525),
.B(n_47),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_471),
.B(n_48),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_546),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_543),
.B(n_561),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_524),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_549),
.B(n_489),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_472),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_497),
.B(n_562),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_549),
.B(n_546),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_516),
.B(n_560),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_470),
.B(n_482),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_516),
.B(n_560),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_470),
.B(n_550),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_482),
.B(n_550),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_494),
.B(n_477),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_477),
.A2(n_487),
.B1(n_519),
.B2(n_518),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_514),
.B(n_519),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_494),
.B(n_477),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_472),
.B(n_564),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_708),
.A2(n_522),
.B(n_532),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_592),
.A2(n_514),
.B1(n_518),
.B2(n_515),
.Y(n_710)
);

OAI321xp33_ASAP7_75t_L g711 ( 
.A1(n_688),
.A2(n_515),
.A3(n_545),
.B1(n_472),
.B2(n_534),
.C(n_520),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_585),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_687),
.A2(n_545),
.B1(n_522),
.B2(n_532),
.Y(n_713)
);

OAI21xp33_ASAP7_75t_L g714 ( 
.A1(n_594),
.A2(n_559),
.B(n_472),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_576),
.B(n_441),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_687),
.B(n_594),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_700),
.A2(n_517),
.B(n_564),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_572),
.B(n_441),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_700),
.A2(n_517),
.B(n_563),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_625),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_702),
.A2(n_563),
.B(n_510),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_702),
.A2(n_563),
.B(n_510),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_563),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_585),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_652),
.B(n_629),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_703),
.A2(n_534),
.B(n_606),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_625),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_699),
.A2(n_701),
.B(n_697),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_645),
.A2(n_534),
.B(n_704),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_617),
.B(n_580),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_707),
.A2(n_659),
.B(n_696),
.Y(n_731)
);

BUFx12f_ASAP7_75t_L g732 ( 
.A(n_662),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_636),
.A2(n_589),
.B1(n_656),
.B2(n_689),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_652),
.B(n_633),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_605),
.A2(n_615),
.B(n_620),
.C(n_626),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_696),
.A2(n_588),
.B(n_678),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_698),
.A2(n_590),
.B1(n_607),
.B2(n_599),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_597),
.B(n_690),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_603),
.B(n_653),
.Y(n_739)
);

NOR2x1_ASAP7_75t_L g740 ( 
.A(n_604),
.B(n_694),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_682),
.A2(n_684),
.B(n_630),
.C(n_681),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_622),
.B(n_640),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_603),
.B(n_601),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_604),
.B(n_624),
.Y(n_744)
);

AOI21x1_ASAP7_75t_L g745 ( 
.A1(n_609),
.A2(n_613),
.B(n_664),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_573),
.B(n_577),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_574),
.B(n_658),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_696),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_666),
.A2(n_671),
.B(n_679),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_633),
.B(n_635),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_635),
.B(n_605),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_658),
.B(n_643),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_578),
.Y(n_753)
);

BUFx4f_ASAP7_75t_L g754 ( 
.A(n_641),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_683),
.A2(n_676),
.B(n_665),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_615),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_620),
.B(n_626),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_673),
.A2(n_660),
.B(n_642),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_661),
.A2(n_595),
.B(n_627),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_SL g760 ( 
.A(n_628),
.B(n_614),
.C(n_582),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_631),
.A2(n_591),
.B1(n_611),
.B2(n_638),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_614),
.B(n_628),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_604),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_631),
.B(n_579),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_624),
.B(n_584),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_SL g766 ( 
.A(n_583),
.B(n_641),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_L g767 ( 
.A1(n_618),
.A2(n_581),
.B(n_600),
.C(n_602),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_616),
.A2(n_674),
.B(n_669),
.C(n_661),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_619),
.A2(n_621),
.B(n_623),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_639),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_624),
.Y(n_771)
);

BUFx8_ASAP7_75t_L g772 ( 
.A(n_598),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_695),
.A2(n_670),
.B1(n_685),
.B2(n_674),
.Y(n_773)
);

BUFx12f_ASAP7_75t_L g774 ( 
.A(n_662),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_593),
.B(n_677),
.Y(n_775)
);

BUFx12f_ASAP7_75t_L g776 ( 
.A(n_667),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_591),
.B(n_657),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_646),
.B(n_649),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_691),
.Y(n_779)
);

AO32x1_ASAP7_75t_L g780 ( 
.A1(n_651),
.A2(n_663),
.A3(n_692),
.B1(n_686),
.B2(n_634),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_650),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_586),
.B(n_637),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_706),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_608),
.A2(n_648),
.B(n_705),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_638),
.B(n_596),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_688),
.A2(n_638),
.B1(n_655),
.B2(n_582),
.Y(n_786)
);

AO22x1_ASAP7_75t_L g787 ( 
.A1(n_693),
.A2(n_612),
.B1(n_680),
.B2(n_647),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_641),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_672),
.A2(n_675),
.B(n_644),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_668),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_610),
.B(n_644),
.Y(n_791)
);

BUFx8_ASAP7_75t_L g792 ( 
.A(n_575),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_641),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_572),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_687),
.B(n_442),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_687),
.B(n_442),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_687),
.B(n_442),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_687),
.B(n_442),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_571),
.B(n_443),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_629),
.B(n_622),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_687),
.B(n_442),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_687),
.B(n_442),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_588),
.A2(n_456),
.B(n_609),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_587),
.B(n_447),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_687),
.B(n_442),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_808)
);

BUFx8_ASAP7_75t_L g809 ( 
.A(n_571),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_587),
.B(n_447),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_612),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_590),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_583),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_687),
.B(n_442),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_687),
.B(n_442),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_592),
.A2(n_687),
.B1(n_654),
.B2(n_580),
.Y(n_816)
);

AO32x2_ASAP7_75t_L g817 ( 
.A1(n_689),
.A2(n_636),
.A3(n_480),
.B1(n_587),
.B2(n_257),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_585),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_687),
.B(n_442),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_696),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_612),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_636),
.A2(n_448),
.B1(n_442),
.B2(n_589),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_687),
.B(n_442),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_687),
.B(n_442),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_587),
.B(n_447),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_696),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_588),
.A2(n_456),
.B(n_609),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_SL g831 ( 
.A1(n_588),
.A2(n_664),
.B(n_642),
.C(n_659),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_590),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_696),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_687),
.B(n_442),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_571),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_L g836 ( 
.A(n_658),
.B(n_592),
.C(n_589),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_636),
.A2(n_448),
.B1(n_442),
.B2(n_589),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_571),
.B(n_443),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_687),
.B(n_442),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_585),
.Y(n_841)
);

AND2x6_ASAP7_75t_L g842 ( 
.A(n_681),
.B(n_705),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_696),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_L g845 ( 
.A(n_592),
.B(n_660),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_687),
.B(n_442),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_687),
.B(n_442),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_687),
.B(n_442),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_636),
.A2(n_448),
.B1(n_442),
.B2(n_589),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_687),
.B(n_442),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_687),
.B(n_442),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_585),
.B(n_629),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_687),
.B(n_442),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_708),
.A2(n_462),
.B(n_700),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_585),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_590),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_590),
.Y(n_860)
);

NAND2x1p5_ASAP7_75t_L g861 ( 
.A(n_585),
.B(n_629),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_687),
.B(n_442),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_687),
.B(n_442),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_696),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_585),
.B(n_629),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_748),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_812),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_845),
.A2(n_799),
.B(n_798),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_716),
.B(n_819),
.Y(n_869)
);

INVx5_ASAP7_75t_L g870 ( 
.A(n_748),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_862),
.B(n_795),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_801),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_808),
.A2(n_824),
.B(n_823),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_L g874 ( 
.A(n_735),
.B(n_756),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_736),
.A2(n_830),
.B(n_805),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_743),
.B(n_796),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_797),
.B(n_800),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_813),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_792),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_803),
.B(n_804),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_724),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_741),
.A2(n_757),
.B(n_752),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_807),
.B(n_814),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_811),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_739),
.A2(n_751),
.B(n_734),
.C(n_750),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_788),
.B(n_821),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_769),
.A2(n_729),
.B(n_745),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_815),
.B(n_826),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_825),
.A2(n_844),
.B(n_838),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_709),
.A2(n_759),
.B(n_847),
.Y(n_891)
);

OAI21x1_ASAP7_75t_L g892 ( 
.A1(n_851),
.A2(n_857),
.B(n_854),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_727),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_758),
.A2(n_749),
.B(n_714),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_714),
.A2(n_831),
.B(n_717),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_732),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_827),
.B(n_834),
.Y(n_898)
);

BUFx8_ASAP7_75t_L g899 ( 
.A(n_774),
.Y(n_899)
);

OAI21x1_ASAP7_75t_L g900 ( 
.A1(n_784),
.A2(n_719),
.B(n_726),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_832),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_L g902 ( 
.A1(n_762),
.A2(n_747),
.B(n_773),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_840),
.B(n_846),
.Y(n_903)
);

OAI22x1_ASAP7_75t_L g904 ( 
.A1(n_781),
.A2(n_786),
.B1(n_773),
.B2(n_791),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_721),
.A2(n_722),
.B(n_778),
.Y(n_905)
);

XNOR2xp5_ASAP7_75t_L g906 ( 
.A(n_760),
.B(n_740),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_835),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_848),
.B(n_849),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_724),
.B(n_858),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_852),
.B(n_853),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_786),
.A2(n_856),
.B1(n_863),
.B2(n_761),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_733),
.A2(n_837),
.B1(n_822),
.B2(n_850),
.Y(n_912)
);

OAI22x1_ASAP7_75t_L g913 ( 
.A1(n_777),
.A2(n_733),
.B1(n_822),
.B2(n_850),
.Y(n_913)
);

AO21x1_ASAP7_75t_L g914 ( 
.A1(n_768),
.A2(n_837),
.B(n_785),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_839),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_794),
.B(n_765),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_775),
.A2(n_782),
.B(n_764),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_713),
.A2(n_746),
.B(n_816),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_718),
.A2(n_738),
.B(n_836),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_790),
.B(n_730),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_802),
.B(n_763),
.Y(n_921)
);

OAI21x1_ASAP7_75t_L g922 ( 
.A1(n_767),
.A2(n_841),
.B(n_712),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_836),
.A2(n_711),
.B(n_742),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_SL g924 ( 
.A1(n_770),
.A2(n_833),
.B(n_864),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_842),
.B(n_737),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_842),
.B(n_783),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_L g927 ( 
.A(n_763),
.B(n_776),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_712),
.A2(n_818),
.B(n_841),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_859),
.A2(n_860),
.B(n_746),
.C(n_789),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_842),
.B(n_818),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_802),
.B(n_777),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_772),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_725),
.A2(n_828),
.B(n_810),
.C(n_806),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_820),
.B(n_864),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_772),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_771),
.B(n_744),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_779),
.A2(n_820),
.B(n_829),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_753),
.A2(n_723),
.B(n_779),
.C(n_770),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_809),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_855),
.B(n_865),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_861),
.A2(n_780),
.B(n_770),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_820),
.A2(n_864),
.B1(n_843),
.B2(n_833),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_817),
.A2(n_780),
.B(n_754),
.Y(n_943)
);

AO21x1_ASAP7_75t_L g944 ( 
.A1(n_817),
.A2(n_780),
.B(n_766),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_829),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_843),
.B(n_833),
.Y(n_946)
);

AO31x2_ASAP7_75t_L g947 ( 
.A1(n_817),
.A2(n_787),
.A3(n_829),
.B(n_843),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_809),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_766),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_788),
.Y(n_950)
);

BUFx2_ASAP7_75t_R g951 ( 
.A(n_792),
.Y(n_951)
);

NOR2x1_ASAP7_75t_L g952 ( 
.A(n_788),
.B(n_754),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_793),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_793),
.A2(n_728),
.B(n_755),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_720),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_801),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_735),
.A2(n_741),
.B(n_757),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_743),
.B(n_576),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_845),
.A2(n_462),
.B(n_798),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_748),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_798),
.A2(n_808),
.B(n_799),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_716),
.B(n_819),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_716),
.B(n_819),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_735),
.A2(n_710),
.A3(n_752),
.B(n_737),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_724),
.B(n_858),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_716),
.B(n_819),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_845),
.A2(n_462),
.B(n_798),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_748),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_716),
.B(n_819),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_716),
.B(n_819),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_819),
.B(n_862),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_716),
.B(n_819),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_735),
.A2(n_741),
.B(n_757),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_763),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_716),
.B(n_819),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_716),
.B(n_819),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_716),
.B(n_819),
.Y(n_978)
);

NAND2x1p5_ASAP7_75t_L g979 ( 
.A(n_724),
.B(n_858),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_798),
.A2(n_808),
.B(n_799),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_735),
.A2(n_756),
.B(n_757),
.C(n_739),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_813),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_735),
.A2(n_756),
.B1(n_762),
.B2(n_757),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_792),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_987)
);

AND2x6_ASAP7_75t_L g988 ( 
.A(n_715),
.B(n_718),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_743),
.B(n_576),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_798),
.A2(n_808),
.B(n_799),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_748),
.Y(n_991)
);

AND2x2_ASAP7_75t_SL g992 ( 
.A(n_762),
.B(n_446),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_993)
);

AO31x2_ASAP7_75t_L g994 ( 
.A1(n_735),
.A2(n_710),
.A3(n_752),
.B(n_737),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_845),
.A2(n_462),
.B(n_798),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_728),
.A2(n_755),
.B(n_731),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_716),
.B(n_819),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_845),
.A2(n_462),
.B(n_798),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_735),
.A2(n_741),
.B(n_757),
.Y(n_1000)
);

BUFx4_ASAP7_75t_SL g1001 ( 
.A(n_813),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_716),
.B(n_819),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_SL g1003 ( 
.A1(n_735),
.A2(n_757),
.B(n_756),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_835),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_931),
.B(n_921),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_1001),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_972),
.B(n_878),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_931),
.B(n_921),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_975),
.B(n_952),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_975),
.B(n_950),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_907),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_894),
.A2(n_1003),
.B(n_917),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_962),
.B(n_967),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_885),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_992),
.A2(n_989),
.B1(n_958),
.B2(n_877),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_904),
.B(n_881),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_899),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_874),
.A2(n_968),
.B(n_959),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_957),
.A2(n_1000),
.B(n_974),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_898),
.B(n_915),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_887),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_915),
.B(n_884),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_869),
.B(n_963),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_901),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_870),
.B(n_882),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_887),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_869),
.B(n_963),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_884),
.B(n_889),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_995),
.A2(n_999),
.B(n_868),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_970),
.B(n_1002),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_971),
.B(n_973),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_957),
.A2(n_974),
.B(n_1000),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_971),
.B(n_973),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_889),
.B(n_908),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_976),
.A2(n_977),
.B1(n_978),
.B2(n_998),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_899),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_976),
.B(n_977),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_978),
.B(n_998),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_982),
.A2(n_902),
.B(n_886),
.C(n_883),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_871),
.A2(n_908),
.B1(n_910),
.B2(n_985),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1004),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_887),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_883),
.A2(n_890),
.B(n_873),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_SL g1044 ( 
.A(n_870),
.B(n_942),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_879),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_983),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_895),
.A2(n_919),
.B(n_923),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_893),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_871),
.B(n_910),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_936),
.B(n_916),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_955),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_949),
.A2(n_906),
.B1(n_948),
.B2(n_880),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_903),
.B(n_902),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_922),
.A2(n_876),
.B(n_905),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_888),
.A2(n_924),
.B(n_997),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_872),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_911),
.B(n_912),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_911),
.B(n_912),
.Y(n_1058)
);

BUFx4f_ASAP7_75t_L g1059 ( 
.A(n_986),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_925),
.B(n_913),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_932),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_935),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_925),
.A2(n_933),
.B1(n_926),
.B2(n_938),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_956),
.B(n_949),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_920),
.B(n_929),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_926),
.B(n_930),
.Y(n_1066)
);

OAI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_940),
.A2(n_953),
.B(n_930),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_945),
.B(n_927),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_939),
.B(n_918),
.C(n_896),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_951),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_914),
.B(n_945),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_988),
.A2(n_942),
.B1(n_944),
.B2(n_937),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_870),
.B(n_991),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_946),
.B(n_969),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_875),
.A2(n_996),
.B(n_987),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_943),
.A2(n_909),
.B(n_979),
.C(n_965),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_870),
.B(n_991),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_994),
.B(n_964),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_965),
.A2(n_979),
.B1(n_934),
.B2(n_897),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_994),
.B(n_964),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_928),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_969),
.B(n_866),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_866),
.B(n_960),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_866),
.B(n_897),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_966),
.A2(n_980),
.B(n_993),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_964),
.B(n_994),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_960),
.B(n_934),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_947),
.A2(n_988),
.B(n_990),
.C(n_981),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_961),
.B(n_954),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_947),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_988),
.B(n_941),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_988),
.B(n_947),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_900),
.B(n_891),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_892),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_984),
.A2(n_972),
.B1(n_962),
.B2(n_970),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_866),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_894),
.A2(n_462),
.B(n_1003),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_877),
.B(n_958),
.Y(n_1098)
);

NAND2x1_ASAP7_75t_L g1099 ( 
.A(n_924),
.B(n_882),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_867),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_972),
.B(n_878),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_931),
.B(n_921),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_866),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_931),
.B(n_921),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_877),
.B(n_958),
.Y(n_1105)
);

AND2x6_ASAP7_75t_L g1106 ( 
.A(n_925),
.B(n_783),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_L g1107 ( 
.A1(n_985),
.A2(n_757),
.B(n_756),
.Y(n_1107)
);

CKINVDCx6p67_ASAP7_75t_R g1108 ( 
.A(n_880),
.Y(n_1108)
);

OAI21xp33_ASAP7_75t_L g1109 ( 
.A1(n_972),
.A2(n_446),
.B(n_442),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_887),
.B(n_641),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_972),
.A2(n_760),
.B1(n_757),
.B2(n_762),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_958),
.B(n_989),
.Y(n_1112)
);

BUFx2_ASAP7_75t_SL g1113 ( 
.A(n_927),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_877),
.B(n_958),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_867),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1001),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_972),
.B(n_878),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_972),
.B(n_762),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_957),
.A2(n_716),
.B(n_739),
.C(n_819),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_931),
.B(n_921),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_972),
.B(n_878),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_867),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_894),
.A2(n_462),
.B(n_1003),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_L g1124 ( 
.A(n_884),
.B(n_735),
.Y(n_1124)
);

BUFx8_ASAP7_75t_L g1125 ( 
.A(n_880),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_882),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_972),
.B(n_878),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_931),
.B(n_921),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_972),
.B(n_878),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_877),
.B(n_958),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_877),
.B(n_958),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_915),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_957),
.A2(n_735),
.B(n_1000),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_877),
.B(n_958),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_867),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_894),
.A2(n_462),
.B(n_1003),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_907),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_885),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_885),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1001),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_972),
.B(n_878),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_931),
.B(n_921),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_894),
.A2(n_462),
.B(n_1003),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1066),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_R g1145 ( 
.A(n_1006),
.B(n_1116),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1024),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_1140),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1135),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1111),
.B(n_1016),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1109),
.A2(n_1118),
.B1(n_1030),
.B2(n_1015),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1014),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1090),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1078),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1118),
.A2(n_1101),
.B1(n_1007),
.B2(n_1127),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1007),
.B(n_1117),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1055),
.A2(n_1054),
.B(n_1075),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1117),
.A2(n_1129),
.B1(n_1127),
.B2(n_1141),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1133),
.A2(n_1019),
.B1(n_1057),
.B2(n_1058),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1085),
.A2(n_1018),
.B(n_1029),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1133),
.A2(n_1019),
.B1(n_1058),
.B2(n_1057),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1106),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1106),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1060),
.B(n_1053),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_SL g1166 ( 
.A(n_1036),
.Y(n_1166)
);

BUFx8_ASAP7_75t_L g1167 ( 
.A(n_1139),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1106),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_1064),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1138),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1028),
.B(n_1034),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1009),
.B(n_1005),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_R g1173 ( 
.A(n_1070),
.B(n_1045),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1121),
.B(n_1129),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1080),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1097),
.A2(n_1143),
.B(n_1123),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1121),
.A2(n_1141),
.B1(n_1031),
.B2(n_1035),
.Y(n_1177)
);

INVx6_ASAP7_75t_L g1178 ( 
.A(n_1010),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1060),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1100),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1132),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1053),
.B(n_1022),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1013),
.B(n_1035),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1106),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1107),
.A2(n_1032),
.B(n_1039),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1132),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1098),
.B(n_1105),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1115),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1041),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1122),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1051),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1089),
.A2(n_1136),
.B(n_1047),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1033),
.A2(n_1038),
.B1(n_1037),
.B2(n_1023),
.Y(n_1193)
);

BUFx8_ASAP7_75t_SL g1194 ( 
.A(n_1017),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1124),
.A2(n_1114),
.B1(n_1134),
.B2(n_1131),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1096),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1073),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1012),
.A2(n_1043),
.B(n_1088),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1096),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1083),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1048),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1041),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1023),
.A2(n_1027),
.B1(n_1110),
.B2(n_1137),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1130),
.B(n_1086),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1107),
.A2(n_1112),
.B1(n_1067),
.B2(n_1069),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1065),
.A2(n_1092),
.B(n_1093),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1011),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1081),
.A2(n_1076),
.B(n_1063),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1056),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1092),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1063),
.A2(n_1050),
.B1(n_1071),
.B2(n_1020),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1083),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1087),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1126),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1027),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1025),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1119),
.B(n_1095),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1095),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1009),
.B(n_1005),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1072),
.A2(n_1079),
.B(n_1091),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1052),
.A2(n_1008),
.B1(n_1128),
.B2(n_1120),
.Y(n_1221)
);

CKINVDCx8_ASAP7_75t_R g1222 ( 
.A(n_1046),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1056),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1102),
.A2(n_1142),
.B1(n_1128),
.B2(n_1120),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1102),
.B(n_1104),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1094),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1104),
.B(n_1062),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1110),
.A2(n_1113),
.B1(n_1068),
.B2(n_1042),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1094),
.A2(n_1079),
.B(n_1074),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1077),
.A2(n_1021),
.B1(n_1026),
.B2(n_1044),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1094),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1082),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1083),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1084),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1077),
.A2(n_1103),
.B(n_1110),
.Y(n_1235)
);

BUFx2_ASAP7_75t_SL g1236 ( 
.A(n_1061),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1059),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1059),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1125),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1108),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1125),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1055),
.A2(n_1054),
.B(n_891),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1111),
.B(n_1016),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1024),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1109),
.A2(n_760),
.B1(n_762),
.B2(n_992),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1118),
.A2(n_762),
.B1(n_992),
.B2(n_316),
.Y(n_1246)
);

CKINVDCx6p67_ASAP7_75t_R g1247 ( 
.A(n_1036),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1065),
.B(n_1099),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1066),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1198),
.A2(n_1157),
.B(n_1176),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1217),
.A2(n_1218),
.A3(n_1153),
.B(n_1175),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1204),
.B(n_1182),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1176),
.B(n_1198),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1152),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1186),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1242),
.A2(n_1160),
.B(n_1192),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1200),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1241),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1185),
.A2(n_1208),
.B(n_1220),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1206),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1210),
.B(n_1156),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1156),
.B(n_1163),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1229),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1154),
.B(n_1174),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1179),
.B(n_1182),
.Y(n_1266)
);

AO21x1_ASAP7_75t_SL g1267 ( 
.A1(n_1205),
.A2(n_1183),
.B(n_1150),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1248),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1179),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1235),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1226),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1149),
.B(n_1243),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1159),
.A2(n_1161),
.B(n_1245),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1231),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1149),
.B(n_1243),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1231),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1203),
.A2(n_1165),
.B(n_1190),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1165),
.A2(n_1188),
.B(n_1180),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1162),
.A2(n_1164),
.B(n_1168),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1235),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1162),
.A2(n_1164),
.B(n_1184),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1194),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1229),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1168),
.B(n_1184),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1144),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1211),
.A2(n_1191),
.B(n_1215),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1171),
.B(n_1177),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1249),
.B(n_1171),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1187),
.B(n_1155),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1213),
.A2(n_1193),
.B(n_1146),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1189),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1202),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1223),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1148),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1244),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1201),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1187),
.B(n_1158),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1195),
.B(n_1214),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1194),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1181),
.B(n_1228),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1233),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1209),
.B(n_1170),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1246),
.B(n_1230),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1200),
.Y(n_1304)
);

INVxp33_ASAP7_75t_L g1305 ( 
.A(n_1227),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1207),
.B(n_1225),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1265),
.A2(n_1221),
.B1(n_1219),
.B2(n_1172),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1251),
.B(n_1236),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1267),
.A2(n_1273),
.B1(n_1303),
.B2(n_1297),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1293),
.Y(n_1310)
);

NOR2x1_ASAP7_75t_L g1311 ( 
.A(n_1290),
.B(n_1212),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1288),
.B(n_1169),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1251),
.B(n_1236),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1270),
.B(n_1268),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1251),
.B(n_1234),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1285),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1254),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1288),
.B(n_1169),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_SL g1319 ( 
.A(n_1303),
.B(n_1222),
.C(n_1238),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_R g1320 ( 
.A(n_1282),
.B(n_1299),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1262),
.B(n_1172),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1251),
.B(n_1151),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1285),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1255),
.B(n_1169),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1255),
.B(n_1151),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1266),
.B(n_1167),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1293),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1264),
.B(n_1216),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1251),
.B(n_1212),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1256),
.A2(n_1224),
.B(n_1232),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1253),
.A2(n_1212),
.B(n_1216),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1279),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1279),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1267),
.A2(n_1239),
.B1(n_1241),
.B2(n_1178),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1273),
.A2(n_1241),
.B1(n_1237),
.B2(n_1178),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1278),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1278),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1279),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1268),
.B(n_1197),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1291),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1300),
.A2(n_1178),
.B1(n_1240),
.B2(n_1237),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1261),
.B(n_1199),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1275),
.B(n_1199),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1275),
.B(n_1199),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1309),
.B(n_1287),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1342),
.B(n_1279),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1342),
.B(n_1279),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1328),
.B(n_1343),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1328),
.B(n_1281),
.Y(n_1349)
);

AOI211xp5_ASAP7_75t_L g1350 ( 
.A1(n_1319),
.A2(n_1300),
.B(n_1287),
.C(n_1305),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1317),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1343),
.B(n_1281),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_L g1353 ( 
.A(n_1334),
.B(n_1273),
.C(n_1306),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1327),
.B(n_1292),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1307),
.A2(n_1273),
.B1(n_1289),
.B2(n_1297),
.Y(n_1355)
);

NOR3xp33_ASAP7_75t_L g1356 ( 
.A(n_1341),
.B(n_1298),
.C(n_1292),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1317),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1324),
.B(n_1268),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1310),
.B(n_1266),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1344),
.B(n_1281),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1314),
.B(n_1281),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1314),
.B(n_1280),
.Y(n_1362)
);

AOI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1340),
.A2(n_1297),
.B1(n_1275),
.B2(n_1272),
.C(n_1298),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1314),
.B(n_1280),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1307),
.A2(n_1335),
.B1(n_1318),
.B2(n_1312),
.Y(n_1365)
);

AOI221xp5_ASAP7_75t_L g1366 ( 
.A1(n_1325),
.A2(n_1272),
.B1(n_1298),
.B2(n_1283),
.C(n_1263),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1316),
.B(n_1252),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1339),
.B(n_1268),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1323),
.B(n_1252),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1322),
.B(n_1273),
.C(n_1306),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1322),
.B(n_1313),
.C(n_1308),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1326),
.B(n_1302),
.Y(n_1372)
);

NAND3xp33_ASAP7_75t_L g1373 ( 
.A(n_1311),
.B(n_1313),
.C(n_1308),
.Y(n_1373)
);

NAND4xp25_ASAP7_75t_L g1374 ( 
.A(n_1315),
.B(n_1302),
.C(n_1294),
.D(n_1296),
.Y(n_1374)
);

NAND3xp33_ASAP7_75t_L g1375 ( 
.A(n_1311),
.B(n_1301),
.C(n_1294),
.Y(n_1375)
);

OAI221xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1329),
.A2(n_1263),
.B1(n_1283),
.B2(n_1247),
.C(n_1239),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1336),
.A2(n_1256),
.B(n_1250),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1323),
.B(n_1301),
.Y(n_1378)
);

NOR3xp33_ASAP7_75t_L g1379 ( 
.A(n_1331),
.B(n_1257),
.C(n_1304),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1339),
.A2(n_1268),
.B1(n_1284),
.B2(n_1277),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1332),
.A2(n_1269),
.B1(n_1296),
.B2(n_1271),
.C(n_1274),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1329),
.B(n_1286),
.C(n_1295),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1321),
.B(n_1222),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1332),
.A2(n_1269),
.B1(n_1276),
.B2(n_1274),
.C(n_1271),
.Y(n_1384)
);

NAND3xp33_ASAP7_75t_L g1385 ( 
.A(n_1315),
.B(n_1268),
.C(n_1286),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1361),
.B(n_1333),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1371),
.B(n_1382),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1361),
.B(n_1333),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1362),
.B(n_1364),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1351),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1362),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1349),
.B(n_1338),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1351),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1357),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1357),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1346),
.B(n_1330),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1377),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1375),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1346),
.B(n_1330),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1347),
.B(n_1330),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1371),
.B(n_1337),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1355),
.A2(n_1277),
.B1(n_1259),
.B2(n_1286),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1352),
.B(n_1277),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1347),
.B(n_1330),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1377),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1360),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1373),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1378),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1382),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1359),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1385),
.B(n_1260),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1393),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1387),
.A2(n_1350),
.B(n_1345),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1398),
.B(n_1366),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1398),
.B(n_1381),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1406),
.B(n_1348),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1390),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1387),
.B(n_1370),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1389),
.B(n_1379),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1387),
.B(n_1370),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1397),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1387),
.B(n_1354),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1397),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1409),
.B(n_1367),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1406),
.B(n_1380),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1393),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1393),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1395),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1397),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1395),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1408),
.Y(n_1431)
);

NOR3xp33_ASAP7_75t_L g1432 ( 
.A(n_1407),
.B(n_1350),
.C(n_1353),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1395),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1397),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1407),
.B(n_1409),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1390),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1407),
.B(n_1384),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1391),
.B(n_1356),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1409),
.B(n_1369),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1391),
.B(n_1372),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1389),
.B(n_1368),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1394),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1405),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1401),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1402),
.A2(n_1353),
.B(n_1375),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1405),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1440),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1415),
.B(n_1408),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1412),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1413),
.B(n_1376),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1417),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1412),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1426),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1426),
.Y(n_1454)
);

NAND2x1_ASAP7_75t_L g1455 ( 
.A(n_1419),
.B(n_1409),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1435),
.B(n_1403),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1441),
.B(n_1425),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1427),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1415),
.B(n_1414),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1414),
.B(n_1408),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1441),
.B(n_1386),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1435),
.B(n_1403),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1427),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1428),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1419),
.B(n_1386),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1428),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1431),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1430),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1430),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1425),
.B(n_1386),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1419),
.B(n_1438),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1419),
.B(n_1386),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_SL g1473 ( 
.A(n_1445),
.B(n_1241),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1417),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1433),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1432),
.B(n_1408),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1431),
.B(n_1388),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1432),
.B(n_1410),
.Y(n_1478)
);

AOI31xp33_ASAP7_75t_L g1479 ( 
.A1(n_1413),
.A2(n_1365),
.A3(n_1173),
.B(n_1383),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1433),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1431),
.B(n_1388),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1417),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1445),
.A2(n_1402),
.B(n_1358),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1437),
.B(n_1410),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1437),
.A2(n_1363),
.B(n_1411),
.C(n_1374),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1422),
.B(n_1401),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1438),
.B(n_1388),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1436),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1440),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1489),
.B(n_1471),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1468),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1468),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1247),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1489),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1455),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1447),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1471),
.B(n_1416),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1457),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1449),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1478),
.B(n_1422),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1442),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1476),
.A2(n_1420),
.B(n_1418),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1452),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1450),
.A2(n_1420),
.B1(n_1418),
.B2(n_1444),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1460),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1455),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1241),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1448),
.B(n_1424),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1453),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1483),
.A2(n_1424),
.B1(n_1439),
.B2(n_1411),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1477),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1454),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1485),
.B(n_1411),
.C(n_1401),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1477),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1477),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1481),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1484),
.B(n_1166),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1486),
.B(n_1439),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1457),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1465),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1481),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1485),
.B(n_1467),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1487),
.B(n_1416),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1481),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1498),
.B(n_1486),
.Y(n_1526)
);

AOI21xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1522),
.A2(n_1473),
.B(n_1462),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1496),
.B(n_1487),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1491),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1491),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1506),
.Y(n_1531)
);

AOI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1513),
.A2(n_1504),
.B1(n_1510),
.B2(n_1500),
.C(n_1505),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1492),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1490),
.B(n_1470),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1513),
.A2(n_1465),
.B1(n_1470),
.B2(n_1472),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1492),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_SL g1537 ( 
.A1(n_1506),
.A2(n_1482),
.B(n_1451),
.C(n_1474),
.Y(n_1537)
);

NOR4xp25_ASAP7_75t_SL g1538 ( 
.A(n_1499),
.B(n_1458),
.C(n_1480),
.D(n_1475),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1490),
.B(n_1472),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1493),
.B(n_1517),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1495),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1490),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1490),
.Y(n_1543)
);

AOI322xp5_ASAP7_75t_L g1544 ( 
.A1(n_1508),
.A2(n_1461),
.A3(n_1399),
.B1(n_1396),
.B2(n_1404),
.C1(n_1400),
.C2(n_1392),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1494),
.B(n_1461),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1525),
.A2(n_1411),
.B1(n_1456),
.B2(n_1462),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1521),
.Y(n_1547)
);

OAI21xp33_ASAP7_75t_L g1548 ( 
.A1(n_1519),
.A2(n_1456),
.B(n_1463),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1502),
.A2(n_1494),
.B1(n_1511),
.B2(n_1515),
.C(n_1516),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_SL g1550 ( 
.A(n_1524),
.B(n_1320),
.C(n_1451),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1521),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1529),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1530),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1540),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

CKINVDCx16_ASAP7_75t_R g1557 ( 
.A(n_1550),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1543),
.B(n_1497),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1536),
.Y(n_1559)
);

XNOR2xp5_ASAP7_75t_L g1560 ( 
.A(n_1532),
.B(n_1524),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1547),
.B(n_1523),
.Y(n_1561)
);

NOR2x1_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1502),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1551),
.B(n_1507),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1526),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1531),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1528),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1545),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1534),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1527),
.B(n_1495),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

AOI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1560),
.A2(n_1549),
.B1(n_1535),
.B2(n_1548),
.C(n_1537),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1565),
.Y(n_1573)
);

NAND3x1_ASAP7_75t_L g1574 ( 
.A(n_1562),
.B(n_1508),
.C(n_1520),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_SL g1575 ( 
.A(n_1555),
.B(n_1538),
.C(n_1541),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1570),
.B(n_1523),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1569),
.A2(n_1502),
.B(n_1546),
.C(n_1538),
.Y(n_1577)
);

OAI211xp5_ASAP7_75t_L g1578 ( 
.A1(n_1569),
.A2(n_1544),
.B(n_1514),
.C(n_1520),
.Y(n_1578)
);

NAND4xp25_ASAP7_75t_L g1579 ( 
.A(n_1563),
.B(n_1520),
.C(n_1518),
.D(n_1499),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1571),
.B(n_1514),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1564),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1566),
.B(n_1503),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1557),
.A2(n_1518),
.B1(n_1501),
.B2(n_1509),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_SL g1585 ( 
.A(n_1577),
.B(n_1555),
.C(n_1563),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1572),
.B(n_1561),
.C(n_1552),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_L g1587 ( 
.A(n_1575),
.B(n_1553),
.Y(n_1587)
);

NAND5xp2_ASAP7_75t_L g1588 ( 
.A(n_1578),
.B(n_1568),
.C(n_1567),
.D(n_1559),
.E(n_1556),
.Y(n_1588)
);

OA22x2_ASAP7_75t_L g1589 ( 
.A1(n_1584),
.A2(n_1554),
.B1(n_1501),
.B2(n_1509),
.Y(n_1589)
);

NOR2x1_ASAP7_75t_L g1590 ( 
.A(n_1573),
.B(n_1503),
.Y(n_1590)
);

NOR2xp67_ASAP7_75t_L g1591 ( 
.A(n_1579),
.B(n_1512),
.Y(n_1591)
);

AND3x4_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1501),
.C(n_1583),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1574),
.A2(n_1512),
.B1(n_1501),
.B2(n_1464),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1581),
.B(n_1237),
.Y(n_1594)
);

NOR3xp33_ASAP7_75t_L g1595 ( 
.A(n_1585),
.B(n_1580),
.C(n_1582),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1586),
.B(n_1147),
.Y(n_1596)
);

OAI211xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1587),
.A2(n_1469),
.B(n_1466),
.C(n_1488),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1588),
.A2(n_1482),
.B1(n_1474),
.B2(n_1446),
.C(n_1434),
.Y(n_1598)
);

NAND2x1_ASAP7_75t_L g1599 ( 
.A(n_1594),
.B(n_1442),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1597),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1599),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1595),
.Y(n_1602)
);

BUFx12f_ASAP7_75t_L g1603 ( 
.A(n_1596),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1598),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1597),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1601),
.B(n_1591),
.Y(n_1606)
);

NOR5xp2_ASAP7_75t_L g1607 ( 
.A(n_1602),
.B(n_1589),
.C(n_1592),
.D(n_1590),
.E(n_1593),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1600),
.Y(n_1608)
);

INVxp33_ASAP7_75t_L g1609 ( 
.A(n_1605),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1601),
.B(n_1237),
.Y(n_1610)
);

NAND3x2_ASAP7_75t_L g1611 ( 
.A(n_1606),
.B(n_1604),
.C(n_1603),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1608),
.A2(n_1603),
.B1(n_1147),
.B2(n_1258),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1610),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1613),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_1609),
.B(n_1612),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1615),
.Y(n_1616)
);

AOI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1615),
.A2(n_1611),
.B(n_1607),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1617),
.A2(n_1616),
.B(n_1240),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1616),
.B(n_1167),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1619),
.A2(n_1240),
.B1(n_1237),
.B2(n_1258),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1618),
.A2(n_1145),
.B(n_1240),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_L g1622 ( 
.A(n_1621),
.B(n_1240),
.C(n_1167),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1622),
.A2(n_1620),
.B1(n_1258),
.B2(n_1196),
.Y(n_1623)
);

OAI221xp5_ASAP7_75t_R g1624 ( 
.A1(n_1623),
.A2(n_1446),
.B1(n_1434),
.B2(n_1421),
.C(n_1443),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1421),
.B(n_1429),
.C(n_1423),
.Y(n_1625)
);


endmodule