module fake_jpeg_23044_n_207 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_207);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_13),
.B1(n_16),
.B2(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_13),
.B1(n_16),
.B2(n_24),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_34),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_23),
.B1(n_18),
.B2(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_50),
.B1(n_29),
.B2(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_41),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_48),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_58),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_26),
.A3(n_27),
.B1(n_17),
.B2(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_37),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_68),
.B1(n_46),
.B2(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_67),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_20),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_66),
.B(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_33),
.B1(n_46),
.B2(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_86),
.B1(n_38),
.B2(n_33),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_48),
.B(n_50),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_60),
.B(n_57),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_40),
.B(n_15),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_27),
.B(n_39),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_57),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_40),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_67),
.C(n_63),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_90),
.B(n_97),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_77),
.B1(n_70),
.B2(n_73),
.Y(n_112)
);

OA21x2_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_46),
.B(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_82),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_78),
.B(n_86),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_110),
.B(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_81),
.B(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_70),
.B1(n_80),
.B2(n_81),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_73),
.B1(n_56),
.B2(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_96),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_118),
.B1(n_116),
.B2(n_107),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_136),
.B1(n_139),
.B2(n_123),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_31),
.B1(n_19),
.B2(n_21),
.C(n_44),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_101),
.B1(n_95),
.B2(n_99),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_102),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_31),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_97),
.B1(n_104),
.B2(n_69),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_68),
.B1(n_55),
.B2(n_42),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_69),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_120),
.A3(n_105),
.B1(n_115),
.B2(n_119),
.C1(n_44),
.C2(n_56),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_144),
.B(n_153),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_105),
.B(n_120),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_92),
.C(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_149),
.C(n_140),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_92),
.C(n_122),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_36),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_55),
.B1(n_42),
.B2(n_44),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_44),
.B1(n_36),
.B2(n_51),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_136),
.A3(n_132),
.B1(n_126),
.B2(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_158),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_7),
.B(n_11),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_162),
.B(n_36),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_21),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_128),
.B(n_51),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_142),
.B1(n_144),
.B2(n_150),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_167),
.C(n_21),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_0),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_149),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_36),
.C(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_177),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_147),
.B1(n_1),
.B2(n_2),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_178),
.B1(n_12),
.B2(n_11),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_172),
.C(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_176),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_21),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_156),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_162),
.B(n_156),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_173),
.B1(n_8),
.B2(n_9),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_11),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_186),
.B(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_8),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_190),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_192),
.B(n_9),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_8),
.C(n_10),
.Y(n_193)
);

AOI21x1_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_180),
.B(n_10),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_181),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_179),
.C(n_10),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_191),
.B(n_12),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_202),
.C(n_197),
.Y(n_205)
);

AOI21x1_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_4),
.B(n_6),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_200),
.Y(n_207)
);


endmodule