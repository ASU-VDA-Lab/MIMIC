module fake_jpeg_1397_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_12),
.B1(n_13),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_16),
.C(n_11),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_22),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_19),
.B(n_2),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI321xp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_26),
.A3(n_1),
.B1(n_6),
.B2(n_8),
.C(n_5),
.Y(n_29)
);


endmodule