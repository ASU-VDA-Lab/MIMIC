module fake_jpeg_16576_n_349 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_21),
.A2(n_14),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_53),
.A2(n_57),
.B1(n_24),
.B2(n_29),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_73),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_19),
.B1(n_47),
.B2(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_27),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_78),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_19),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_105),
.B(n_58),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_19),
.A3(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_87),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_19),
.B1(n_39),
.B2(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_103),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_0),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_19),
.B1(n_49),
.B2(n_41),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_91),
.B1(n_102),
.B2(n_65),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_49),
.B1(n_24),
.B2(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_27),
.C(n_32),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_26),
.C(n_65),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_30),
.B1(n_24),
.B2(n_23),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_30),
.B1(n_24),
.B2(n_23),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_71),
.B1(n_66),
.B2(n_59),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_99),
.B1(n_101),
.B2(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_30),
.B1(n_26),
.B2(n_27),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

OR2x4_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_52),
.B(n_32),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_14),
.B1(n_29),
.B2(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_55),
.B1(n_54),
.B2(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_89),
.B1(n_105),
.B2(n_55),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_62),
.B1(n_59),
.B2(n_64),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_103),
.B1(n_78),
.B2(n_33),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_134),
.C(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_78),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_135),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_127),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_69),
.B(n_61),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_129),
.B1(n_97),
.B2(n_95),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_77),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_26),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_33),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_110),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_101),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_82),
.B1(n_81),
.B2(n_90),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_154),
.B1(n_130),
.B2(n_120),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_141),
.A2(n_144),
.B1(n_4),
.B2(n_5),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_82),
.B1(n_79),
.B2(n_81),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_92),
.B(n_98),
.C(n_85),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_157),
.C(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_89),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_100),
.B1(n_94),
.B2(n_96),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_33),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_7),
.C(n_9),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_106),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_119),
.B(n_111),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_0),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_147),
.B1(n_165),
.B2(n_146),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_156),
.B1(n_159),
.B2(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_13),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_103),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_119),
.B(n_2),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_171),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_194),
.B1(n_198),
.B2(n_202),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_111),
.A3(n_116),
.B1(n_135),
.B2(n_126),
.C1(n_123),
.C2(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_175),
.B(n_180),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_176),
.B(n_179),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_126),
.B1(n_116),
.B2(n_137),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_177),
.A2(n_181),
.B1(n_183),
.B2(n_193),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_126),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_131),
.B1(n_135),
.B2(n_109),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_187),
.B1(n_176),
.B2(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_109),
.B1(n_33),
.B2(n_4),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_2),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_185),
.B(n_206),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_2),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_3),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_191),
.B(n_166),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_3),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_203),
.B1(n_204),
.B2(n_163),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_145),
.B(n_6),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.C(n_205),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_9),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_139),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_10),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_207),
.B(n_208),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_151),
.B(n_140),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_154),
.B1(n_142),
.B2(n_140),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_221),
.B1(n_190),
.B2(n_196),
.Y(n_247)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_163),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_200),
.C(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_219),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_184),
.B(n_180),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_234),
.Y(n_242)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_151),
.B1(n_159),
.B2(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_143),
.B1(n_168),
.B2(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_178),
.B(n_143),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_183),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_204),
.Y(n_243)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_245),
.Y(n_280)
);

NAND4xp25_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_168),
.C(n_187),
.D(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_188),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_178),
.C(n_172),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_251),
.C(n_253),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_198),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_257),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_188),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_203),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_202),
.B1(n_193),
.B2(n_199),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_214),
.B1(n_222),
.B2(n_211),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_185),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_215),
.C(n_207),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_13),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_209),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_261),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_13),
.B1(n_214),
.B2(n_218),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_219),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_251),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_276),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_211),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_249),
.B(n_217),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_228),
.C(n_230),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_273),
.C(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_230),
.C(n_225),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_242),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_227),
.C(n_210),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_250),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_258),
.B1(n_238),
.B2(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_298),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_213),
.B(n_236),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_260),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_297),
.B1(n_236),
.B2(n_240),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_241),
.B1(n_244),
.B2(n_240),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_241),
.B1(n_244),
.B2(n_273),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_280),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_311),
.C(n_313),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_272),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_297),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_293),
.B1(n_287),
.B2(n_296),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_231),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_263),
.C(n_277),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_257),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_298),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_264),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_280),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_263),
.C(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_318),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_321),
.C(n_314),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_295),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_325),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_283),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_295),
.B1(n_268),
.B2(n_271),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_326),
.B1(n_311),
.B2(n_301),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_226),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_305),
.Y(n_327)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_333),
.C(n_319),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_334),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_303),
.C(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_307),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_309),
.B(n_255),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_320),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_332),
.A2(n_323),
.B(n_321),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_339),
.B(n_340),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_231),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_341),
.A2(n_333),
.B(n_330),
.C(n_329),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_341),
.C(n_337),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_344),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_336),
.B(n_342),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_347),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_256),
.Y(n_349)
);


endmodule