module fake_jpeg_18221_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_14),
.C(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_45),
.C(n_47),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_28),
.B1(n_18),
.B2(n_17),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_14),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_29),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_21),
.B1(n_26),
.B2(n_23),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_57),
.B1(n_15),
.B2(n_22),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_15),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_26),
.B1(n_23),
.B2(n_19),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_62),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_19),
.A3(n_28),
.B1(n_22),
.B2(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_76),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_34),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_41),
.C(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_33),
.B1(n_39),
.B2(n_27),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_72),
.B1(n_86),
.B2(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_30),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_33),
.B1(n_17),
.B2(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_79),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_13),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_1),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_96),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_80),
.B1(n_82),
.B2(n_63),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_65),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_59),
.B(n_9),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_11),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_83),
.Y(n_124)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_117),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_84),
.B(n_73),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_115),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_69),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_75),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_84),
.C(n_68),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_105),
.B1(n_106),
.B2(n_97),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_101),
.B1(n_95),
.B2(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_130),
.B1(n_137),
.B2(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_93),
.B1(n_92),
.B2(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_88),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_105),
.B1(n_97),
.B2(n_91),
.Y(n_137)
);

BUFx12f_ASAP7_75t_SL g138 ( 
.A(n_136),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_110),
.B(n_116),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_98),
.A3(n_112),
.B1(n_100),
.B2(n_121),
.C1(n_96),
.C2(n_117),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_133),
.C(n_126),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_137),
.C(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_129),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_123),
.B1(n_122),
.B2(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_147),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_124),
.C(n_120),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_135),
.C(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_153),
.C(n_145),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_160),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_143),
.B1(n_146),
.B2(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_90),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_157),
.A3(n_148),
.B1(n_158),
.B2(n_156),
.C1(n_139),
.C2(n_102),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_168),
.B(n_102),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_78),
.C(n_85),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_170),
.B(n_11),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_163),
.C(n_81),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_8),
.Y(n_172)
);


endmodule