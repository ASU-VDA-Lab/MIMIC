module real_jpeg_32773_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g296 ( 
.A(n_0),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.A3(n_30),
.B1(n_34),
.B2(n_42),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_43),
.B1(n_140),
.B2(n_144),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_1),
.B(n_148),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_1),
.A2(n_52),
.B1(n_290),
.B2(n_300),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_1),
.A2(n_331),
.B(n_335),
.C(n_337),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_1),
.B(n_336),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_44),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_84),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_2),
.A2(n_84),
.B1(n_275),
.B2(n_278),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_2),
.A2(n_84),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_3),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_3),
.Y(n_341)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_6),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_6),
.A2(n_155),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_6),
.A2(n_155),
.B1(n_276),
.B2(n_291),
.Y(n_290)
);

AO22x1_ASAP7_75t_L g320 ( 
.A1(n_6),
.A2(n_155),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_7),
.A2(n_183),
.B1(n_184),
.B2(n_188),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_7),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_7),
.A2(n_183),
.B1(n_217),
.B2(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_9),
.A2(n_384),
.B1(n_386),
.B2(n_387),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_9),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_10),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_11),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_199),
.B(n_202),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_11),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_11),
.A2(n_63),
.B1(n_416),
.B2(n_419),
.Y(n_415)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_12),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_13),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_13),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_14),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_14),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_15),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_15),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_15),
.A2(n_112),
.B1(n_223),
.B2(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_15),
.A2(n_112),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_16),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_16),
.A2(n_74),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_393),
.B1(n_394),
.B2(n_444),
.Y(n_18)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_19),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_207),
.B(n_311),
.C(n_391),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_156),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_21),
.B(n_156),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_122),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_22),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_50),
.B1(n_79),
.B2(n_80),
.Y(n_22)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_23),
.B(n_80),
.Y(n_194)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_29),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_29),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_29),
.Y(n_172)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

AO21x2_ASAP7_75t_L g124 ( 
.A1(n_34),
.A2(n_125),
.B(n_132),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_37),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_37),
.Y(n_418)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_39),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_SL g168 ( 
.A(n_43),
.B(n_169),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_43),
.A2(n_245),
.B(n_249),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_43),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_43),
.B(n_121),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_43),
.B(n_231),
.Y(n_303)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_49),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_49),
.Y(n_205)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_58),
.B1(n_68),
.B2(n_72),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_51),
.A2(n_72),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_51),
.A2(n_273),
.B1(n_282),
.B2(n_283),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_51),
.B(n_182),
.Y(n_389)
);

AO22x1_ASAP7_75t_L g426 ( 
.A1(n_51),
.A2(n_68),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_52),
.A2(n_222),
.B1(n_230),
.B2(n_234),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_52),
.A2(n_274),
.B1(n_290),
.B2(n_293),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_55),
.Y(n_233)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_55),
.Y(n_285)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_56),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_57),
.Y(n_187)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_57),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_58),
.Y(n_234)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_61),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_62),
.Y(n_385)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_65),
.Y(n_387)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_67),
.Y(n_277)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_68),
.Y(n_388)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_78),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_78),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_81),
.A2(n_122),
.B1(n_123),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_81),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_88),
.B1(n_111),
.B2(n_120),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_83),
.A2(n_89),
.B1(n_121),
.B2(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_88),
.A2(n_120),
.B1(n_213),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_89),
.A2(n_121),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_89),
.A2(n_121),
.B1(n_198),
.B2(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_89),
.Y(n_439)
);

AO21x2_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_97),
.B(n_102),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_96),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_97),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_118),
.Y(n_354)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

AO22x1_ASAP7_75t_SL g434 ( 
.A1(n_120),
.A2(n_435),
.B1(n_439),
.B2(n_440),
.Y(n_434)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_139),
.B1(n_147),
.B2(n_149),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_147),
.B1(n_149),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_124),
.A2(n_147),
.B1(n_159),
.B2(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_124),
.A2(n_147),
.B1(n_356),
.B2(n_415),
.Y(n_414)
);

NAND2xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_171),
.B1(n_173),
.B2(n_175),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_136),
.Y(n_351)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_146),
.Y(n_362)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_191),
.B1(n_192),
.B2(n_206),
.Y(n_156)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_158),
.B(n_168),
.C(n_177),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_161),
.Y(n_359)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_164),
.Y(n_375)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_165),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_177),
.B2(n_178),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g329 ( 
.A(n_169),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_170),
.B(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_173),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_174),
.Y(n_380)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_190),
.Y(n_430)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_193),
.B(n_196),
.C(n_206),
.Y(n_315)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_238),
.B(n_310),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_235),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_210),
.B(n_235),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.C(n_221),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_211),
.A2(n_219),
.B1(n_220),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_255),
.B1(n_265),
.B2(n_266),
.Y(n_254)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_270),
.B(n_309),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_267),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_241),
.B(n_267),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_253),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_242),
.A2(n_243),
.B1(n_253),
.B2(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_287),
.B(n_308),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_286),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_272),
.B(n_286),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx2_ASAP7_75t_SL g306 ( 
.A(n_277),
.Y(n_306)
);

BUFx2_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_298),
.B(n_307),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_297),
.Y(n_307)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_315),
.B(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_363),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_317),
.B(n_364),
.C(n_390),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_348),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_318),
.B(n_349),
.C(n_355),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_328),
.B(n_330),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22x1_ASAP7_75t_L g401 ( 
.A1(n_320),
.A2(n_329),
.B1(n_402),
.B2(n_413),
.Y(n_401)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_337),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_342),
.B1(n_345),
.B2(n_347),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_341),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_355),
.Y(n_348)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_390),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_382),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_382),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_370),
.B1(n_376),
.B2(n_381),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_388),
.B(n_389),
.Y(n_382)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_383),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_442),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_397),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_422),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_414),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_441),
.Y(n_422)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_434),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);


endmodule