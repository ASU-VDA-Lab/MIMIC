module fake_jpeg_10408_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_25),
.Y(n_32)
);

CKINVDCx9p33_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_38),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_11),
.B1(n_20),
.B2(n_19),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_18),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_20),
.B1(n_11),
.B2(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_16),
.B1(n_14),
.B2(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_28),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_45),
.B1(n_49),
.B2(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_14),
.B1(n_16),
.B2(n_10),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_31),
.C(n_26),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_43),
.B1(n_60),
.B2(n_12),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_31),
.C(n_22),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_29),
.B(n_23),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_53),
.B(n_58),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_37),
.Y(n_56)
);

OAI322xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_21),
.A3(n_27),
.B1(n_17),
.B2(n_15),
.C1(n_24),
.C2(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_21),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_42),
.B1(n_41),
.B2(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_56),
.B1(n_54),
.B2(n_50),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_68),
.Y(n_74)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_17),
.CI(n_15),
.CON(n_77),
.SN(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_76),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_27),
.C(n_24),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_74),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_82),
.B(n_78),
.C(n_2),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_73),
.B(n_77),
.C(n_72),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_84),
.B(n_3),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_SL g84 ( 
.A(n_82),
.B(n_2),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_6),
.B(n_8),
.Y(n_86)
);

OAI33xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_60),
.B3(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_9),
.Y(n_88)
);


endmodule