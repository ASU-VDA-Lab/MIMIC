module fake_jpeg_11777_n_65 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_65);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_14),
.Y(n_30)
);

OR2x2_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_21),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_17),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_24),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.C(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_30),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_19),
.B(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

XOR2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_18),
.B1(n_38),
.B2(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_39),
.C(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_30),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_47),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_55),
.B1(n_49),
.B2(n_7),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_48),
.C(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_53),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_49),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_1),
.B(n_2),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_1),
.B(n_2),
.C(n_3),
.D(n_62),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_3),
.B(n_30),
.Y(n_65)
);


endmodule