module fake_jpeg_436_n_505 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_505);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_505;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_11),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_5),
.B(n_1),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_51),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_49),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_73),
.Y(n_131)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_34),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_76),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_38),
.A2(n_48),
.B(n_45),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_45),
.C(n_47),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_38),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_37),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_28),
.B(n_0),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g192 ( 
.A(n_101),
.B(n_37),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_23),
.B1(n_29),
.B2(n_25),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_110),
.A2(n_126),
.B1(n_144),
.B2(n_145),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_138),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_29),
.B1(n_25),
.B2(n_47),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_125),
.A2(n_133),
.B1(n_26),
.B2(n_19),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_59),
.A2(n_47),
.B1(n_29),
.B2(n_25),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_51),
.B(n_43),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_60),
.A2(n_29),
.B1(n_25),
.B2(n_47),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_46),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_49),
.B(n_43),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_139),
.B(n_84),
.Y(n_199)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_46),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_44),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_81),
.A2(n_42),
.B1(n_40),
.B2(n_22),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_53),
.B(n_24),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_26),
.Y(n_206)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_54),
.B(n_31),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_33),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_157),
.Y(n_249)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_158),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_160),
.A2(n_168),
.B1(n_129),
.B2(n_149),
.Y(n_240)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_90),
.B1(n_85),
.B2(n_61),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_170),
.B(n_180),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_131),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_174),
.B(n_176),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_96),
.B(n_33),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_58),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_179),
.B(n_185),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_58),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_187),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_32),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_115),
.A2(n_93),
.B1(n_19),
.B2(n_31),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_189),
.A2(n_198),
.B1(n_209),
.B2(n_16),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_32),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_191),
.B(n_196),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_192),
.B(n_194),
.C(n_203),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

OR2x2_ASAP7_75t_SL g194 ( 
.A(n_106),
.B(n_24),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_130),
.A2(n_24),
.B(n_26),
.C(n_37),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_111),
.B(n_103),
.C(n_112),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_30),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_75),
.B1(n_79),
.B2(n_76),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_199),
.A2(n_207),
.B1(n_173),
.B2(n_203),
.Y(n_229)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_143),
.B(n_30),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_139),
.B(n_75),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_6),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_107),
.B(n_0),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_107),
.B(n_1),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_1),
.Y(n_227)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_99),
.Y(n_212)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_127),
.B(n_149),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_214),
.A2(n_252),
.B(n_171),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_220),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_210),
.A2(n_153),
.B1(n_108),
.B2(n_146),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_223),
.A2(n_237),
.B1(n_239),
.B2(n_243),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_227),
.B(n_9),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_229),
.A2(n_244),
.B1(n_254),
.B2(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_121),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_242),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_135),
.B(n_127),
.C(n_123),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_233),
.A2(n_242),
.B(n_220),
.C(n_261),
.D(n_252),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_168),
.B1(n_164),
.B2(n_162),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_161),
.A2(n_146),
.B1(n_108),
.B2(n_135),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_240),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_199),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_160),
.A2(n_129),
.B1(n_19),
.B2(n_7),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_166),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_189),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_195),
.A2(n_6),
.B(n_7),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_175),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_165),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_262),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_255),
.C(n_248),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_273),
.C(n_308),
.Y(n_330)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_167),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_274),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_159),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_234),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_256),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_277),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_183),
.C(n_163),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_266),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_200),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_285),
.Y(n_337)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_198),
.B1(n_205),
.B2(n_213),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_294),
.B1(n_240),
.B2(n_245),
.Y(n_315)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_284),
.B(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_197),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_157),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_290),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_180),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_292),
.B(n_299),
.Y(n_327)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_233),
.A2(n_190),
.B1(n_184),
.B2(n_180),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_295),
.B(n_297),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_262),
.A2(n_212),
.B1(n_188),
.B2(n_158),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_310),
.B1(n_243),
.B2(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_298),
.B(n_300),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_247),
.B(n_9),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_219),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_304),
.Y(n_344)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_306),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_247),
.B(n_219),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_216),
.B(n_221),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_241),
.B(n_188),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_261),
.B(n_11),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_241),
.A2(n_193),
.B1(n_172),
.B2(n_14),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_214),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_311),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_220),
.B(n_263),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_313),
.A2(n_296),
.B(n_283),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_314),
.B(n_324),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_315),
.A2(n_325),
.B1(n_326),
.B2(n_297),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_239),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_338),
.C(n_341),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_263),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_270),
.A2(n_257),
.B1(n_254),
.B2(n_244),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_285),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_339),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_275),
.A2(n_222),
.B(n_217),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_331),
.B(n_310),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_270),
.A2(n_251),
.B1(n_226),
.B2(n_238),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_351),
.B1(n_275),
.B2(n_280),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_333),
.A2(n_294),
.B(n_272),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_267),
.B(n_222),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_274),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_279),
.C(n_303),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_250),
.C(n_221),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_348),
.C(n_295),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_217),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_349),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_265),
.B(n_216),
.C(n_249),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_276),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_291),
.A2(n_251),
.B1(n_238),
.B2(n_226),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_344),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_356),
.B1(n_363),
.B2(n_364),
.Y(n_387)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_359),
.A2(n_360),
.B(n_348),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_281),
.B1(n_271),
.B2(n_269),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_382),
.B1(n_336),
.B2(n_320),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_324),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_332),
.A2(n_316),
.B1(n_331),
.B2(n_333),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_350),
.B(n_284),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_304),
.C(n_300),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_372),
.C(n_376),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_352),
.Y(n_368)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_344),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_371),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_312),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_268),
.C(n_282),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_316),
.A2(n_322),
.B1(n_323),
.B2(n_337),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_373),
.A2(n_379),
.B1(n_343),
.B2(n_342),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_313),
.A2(n_293),
.B(n_290),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_12),
.B(n_13),
.Y(n_413)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_268),
.C(n_288),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_286),
.C(n_249),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_381),
.C(n_386),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_305),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_378),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_218),
.C(n_232),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_321),
.A2(n_302),
.B1(n_246),
.B2(n_228),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_346),
.B(n_218),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_321),
.B(n_246),
.Y(n_384)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_337),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_193),
.C(n_172),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_370),
.A2(n_385),
.B1(n_364),
.B2(n_360),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_388),
.A2(n_394),
.B1(n_411),
.B2(n_374),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_389),
.A2(n_397),
.B(n_405),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_365),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_401),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_356),
.A2(n_325),
.B1(n_342),
.B2(n_331),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_367),
.C(n_372),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_368),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_345),
.B1(n_319),
.B2(n_340),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_402),
.A2(n_375),
.B1(n_386),
.B2(n_359),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_369),
.A2(n_351),
.B1(n_319),
.B2(n_336),
.Y(n_405)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_355),
.B(n_320),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_409),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_355),
.B(n_335),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_373),
.A2(n_352),
.B1(n_335),
.B2(n_334),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_334),
.B1(n_228),
.B2(n_14),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_412),
.A2(n_358),
.B1(n_380),
.B2(n_357),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_12),
.B(n_13),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_383),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_418),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_375),
.B1(n_362),
.B2(n_382),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_419),
.A2(n_414),
.B1(n_412),
.B2(n_398),
.Y(n_445)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_391),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_391),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_366),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_423),
.B(n_428),
.Y(n_446)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_392),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_426),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_430),
.Y(n_453)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_393),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_377),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_397),
.A2(n_395),
.B(n_388),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_429),
.A2(n_395),
.B(n_405),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_376),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_431),
.A2(n_410),
.B1(n_400),
.B2(n_406),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_436),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_354),
.C(n_381),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_433),
.B(n_434),
.C(n_435),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_403),
.B(n_354),
.C(n_14),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_12),
.C(n_15),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_413),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_441),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_422),
.C(n_424),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_436),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_438),
.B(n_410),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_451),
.Y(n_459)
);

AO221x1_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_411),
.B1(n_394),
.B2(n_392),
.C(n_396),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_448),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_396),
.B1(n_393),
.B2(n_16),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_420),
.A2(n_419),
.B1(n_429),
.B2(n_423),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_456),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_437),
.C(n_433),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_15),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_416),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_15),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_432),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_449),
.B(n_434),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_460),
.B(n_464),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_430),
.C(n_428),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_462),
.C(n_456),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_427),
.C(n_435),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_472),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_418),
.B(n_415),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_468),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_421),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_470),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_454),
.B(n_426),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_443),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g472 ( 
.A1(n_439),
.A2(n_16),
.A3(n_440),
.B1(n_446),
.B2(n_450),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_473),
.Y(n_474)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_474),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_441),
.B(n_446),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_481),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_465),
.A2(n_450),
.B1(n_440),
.B2(n_439),
.Y(n_476)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_483),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_473),
.A2(n_448),
.B1(n_455),
.B2(n_445),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_466),
.A2(n_451),
.B(n_452),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_484),
.A2(n_457),
.B(n_16),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_480),
.A2(n_459),
.B1(n_462),
.B2(n_461),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_484),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_471),
.C(n_452),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_482),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_489),
.B(n_478),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_492),
.B(n_495),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_494),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_477),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_490),
.Y(n_496)
);

AOI21xp33_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_475),
.B(n_480),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_493),
.B(n_488),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_500),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g501 ( 
.A1(n_499),
.A2(n_491),
.B(n_481),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_498),
.B1(n_501),
.B2(n_488),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_485),
.C(n_474),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_476),
.Y(n_505)
);


endmodule