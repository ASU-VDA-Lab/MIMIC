module fake_jpeg_14145_n_236 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_0),
.B(n_1),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_17),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_60),
.B(n_30),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_63),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

OR2x4_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_24),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_55),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_27),
.B(n_21),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_36),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_37),
.B1(n_44),
.B2(n_40),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_95),
.B1(n_75),
.B2(n_72),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_98),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_73),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_37),
.B1(n_45),
.B2(n_41),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_48),
.B(n_36),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_33),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_25),
.B1(n_30),
.B2(n_17),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_45),
.B1(n_41),
.B2(n_33),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_106),
.B1(n_109),
.B2(n_112),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_29),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_103),
.Y(n_136)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_114),
.Y(n_117)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_71),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_88),
.B(n_86),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_100),
.C(n_105),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_126),
.B(n_135),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_89),
.B(n_85),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_127),
.B1(n_139),
.B2(n_121),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_71),
.B1(n_78),
.B2(n_75),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_110),
.B1(n_115),
.B2(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_86),
.B(n_80),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_95),
.A2(n_94),
.B1(n_96),
.B2(n_100),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_108),
.B1(n_87),
.B2(n_111),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_98),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_150),
.C(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_148),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_130),
.B1(n_138),
.B2(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_156),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_99),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_106),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_157),
.C(n_3),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_117),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_100),
.C(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_136),
.C(n_117),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_120),
.B(n_138),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_170),
.B(n_174),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_131),
.B(n_119),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_146),
.B1(n_150),
.B2(n_145),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_132),
.B1(n_124),
.B2(n_122),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_171),
.B1(n_172),
.B2(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_126),
.B1(n_130),
.B2(n_78),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_107),
.B(n_2),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_1),
.B(n_2),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_11),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_181),
.B(n_11),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_151),
.B1(n_160),
.B2(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_183),
.A2(n_187),
.B1(n_189),
.B2(n_191),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_171),
.B2(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_145),
.C(n_12),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_177),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_165),
.B(n_170),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_204),
.B(n_207),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_166),
.C(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_180),
.B(n_176),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_210),
.C(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_188),
.C(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_196),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_185),
.C(n_195),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_216),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_195),
.B1(n_192),
.B2(n_189),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_198),
.B(n_191),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_194),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_205),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_219),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_209),
.B(n_210),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_208),
.B(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_200),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_227),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_225),
.B1(n_173),
.B2(n_5),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_222),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_193),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_198),
.B(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_3),
.B(n_4),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_4),
.Y(n_232)
);

AOI321xp33_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_228),
.A3(n_230),
.B1(n_7),
.B2(n_5),
.C(n_6),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_233),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_7),
.Y(n_236)
);


endmodule