module real_jpeg_10106_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_308, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_308;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx24_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_1),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_58),
.B1(n_65),
.B2(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_40),
.B1(n_50),
.B2(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_2),
.A2(n_58),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_58),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_2),
.A2(n_27),
.B1(n_33),
.B2(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_2),
.B(n_52),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_2),
.A2(n_42),
.B(n_46),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_2),
.A2(n_40),
.B1(n_50),
.B2(n_163),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_7),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_40),
.B1(n_50),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_54),
.B1(n_58),
.B2(n_65),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_10),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_58),
.B1(n_65),
.B2(n_145),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_145),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_10),
.A2(n_40),
.B1(n_50),
.B2(n_145),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_58),
.B1(n_65),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_11),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_154),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_154),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_11),
.A2(n_40),
.B1(n_50),
.B2(n_154),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_12),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_66),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_40),
.B1(n_50),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_13),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_103),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_13),
.A2(n_58),
.B1(n_65),
.B2(n_103),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_103),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_15),
.A2(n_36),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_15),
.A2(n_36),
.B1(n_58),
.B2(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_15),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_20),
.B(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_91),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_21),
.A2(n_22),
.B1(n_71),
.B2(n_72),
.Y(n_299)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_55),
.B2(n_70),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_25),
.A2(n_38),
.B(n_70),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_25),
.A2(n_26),
.B1(n_56),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_27),
.A2(n_33),
.B1(n_144),
.B2(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_27),
.A2(n_97),
.B(n_147),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_27),
.A2(n_34),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_27),
.A2(n_33),
.B1(n_210),
.B2(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_27),
.A2(n_196),
.B(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_28),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_28),
.A2(n_32),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_29),
.A2(n_30),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_29),
.B(n_63),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_29),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_30),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_155)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_32),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_32),
.B(n_96),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_33),
.B(n_163),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_33),
.A2(n_95),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_48),
.B(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_39),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_39),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_39),
.A2(n_44),
.B1(n_246),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_39),
.A2(n_44),
.B1(n_102),
.B2(n_255),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_40),
.A2(n_41),
.B(n_163),
.C(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_44),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_78),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g188 ( 
.A(n_46),
.B(n_163),
.CON(n_188),
.SN(n_188)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_49),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_52),
.A2(n_119),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_53),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_56),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_64),
.B(n_67),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_62),
.B1(n_64),
.B2(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_57),
.A2(n_62),
.B(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_62),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_57),
.A2(n_62),
.B1(n_153),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_57),
.A2(n_62),
.B1(n_178),
.B2(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_57),
.A2(n_84),
.B(n_186),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_60),
.Y(n_61)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_65),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_58),
.B(n_78),
.Y(n_194)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_62),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_62),
.A2(n_87),
.B(n_99),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_65),
.A2(n_80),
.B1(n_188),
.B2(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_68),
.A2(n_86),
.B(n_89),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_83),
.B(n_90),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_77),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_77),
.A2(n_81),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_77),
.A2(n_126),
.B(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_81),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_113),
.B1(n_114),
.B2(n_131),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_91),
.A2(n_92),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.C(n_105),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_93),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_94),
.B(n_98),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_107),
.A2(n_123),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_107),
.A2(n_123),
.B1(n_206),
.B2(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_132),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_123),
.A2(n_242),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_283),
.A3(n_295),
.B1(n_300),
.B2(n_306),
.C(n_308),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_248),
.C(n_279),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_222),
.B(n_247),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_199),
.B(n_221),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_181),
.B(n_198),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_172),
.B(n_180),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_160),
.B(n_171),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_148),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_159),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_166),
.B(n_170),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_162),
.B(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_182),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.CI(n_179),
.CON(n_175),
.SN(n_175)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_192),
.B2(n_197),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_191),
.C(n_197),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_215),
.B2(n_216),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_218),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_214),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.C(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_217),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_224),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_236),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_226),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_235),
.C(n_236),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_231),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_233),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_240),
.C(n_243),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_266),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_266),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.C(n_264),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_253),
.C(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_259),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_256),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_275),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_275),
.C(n_276),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_271),
.C(n_274),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_301),
.B(n_305),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_286),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_292),
.C(n_294),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_301)
);


endmodule