module real_jpeg_4267_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_46),
.B1(n_71),
.B2(n_76),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_46),
.B1(n_125),
.B2(n_129),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_2),
.A2(n_46),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_3),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_30),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_30),
.B1(n_68),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_3),
.B(n_96),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_3),
.A2(n_252),
.B(n_254),
.C(n_260),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_3),
.B(n_40),
.C(n_85),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_3),
.B(n_131),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_3),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_3),
.B(n_51),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_4),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_4),
.A2(n_109),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_4),
.A2(n_109),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_4),
.A2(n_109),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_6),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_10),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_10),
.A2(n_40),
.B1(n_64),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_10),
.A2(n_64),
.B1(n_98),
.B2(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_357),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_219),
.B(n_355),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_189),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_15),
.B(n_189),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_15),
.B(n_359),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_15),
.B(n_359),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_154),
.CI(n_162),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_87),
.B2(n_88),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_17),
.B(n_89),
.C(n_122),
.Y(n_381)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_19),
.B(n_49),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_20),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_21),
.Y(n_156)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_25),
.A2(n_37),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_25),
.B(n_37),
.Y(n_230)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_30),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_30),
.B(n_94),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_30),
.A2(n_255),
.B(n_257),
.Y(n_254)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_31),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_35),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_36),
.A2(n_165),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_37),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_37),
.B(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_42),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_48),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_58),
.B(n_69),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_50),
.A2(n_159),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_50),
.B(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_51),
.B(n_70),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_51),
.B(n_267),
.Y(n_283)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_54),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_63),
.Y(n_259)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_69),
.B(n_283),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_69),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_79),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_73),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_75),
.Y(n_271)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_79),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_79),
.B(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_83),
.Y(n_268)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_122),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_106),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_91),
.B(n_111),
.Y(n_235)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_91),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_94),
.Y(n_110)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_96),
.B(n_107),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_96),
.B(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_96),
.Y(n_370)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_97),
.B(n_148),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_106),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_111),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_120),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_140),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_123),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_130),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_141),
.B(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_131),
.B(n_215),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_131),
.A2(n_239),
.B(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_135),
.Y(n_256)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_140),
.B(n_241),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_141),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_142),
.B(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_145),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_148),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_149),
.Y(n_213)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_155),
.A2(n_161),
.B1(n_251),
.B2(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_155),
.B(n_158),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_155),
.A2(n_161),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_160),
.B(n_266),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_179),
.C(n_181),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_172),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_164),
.B(n_172),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B(n_168),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_168),
.B(n_287),
.Y(n_317)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_173),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_188),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_218),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_190),
.B(n_218),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_193),
.B(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.C(n_210),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_194),
.B(n_210),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_196),
.B(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_200),
.Y(n_232)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_204),
.A3(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_339),
.B(n_352),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_272),
.B(n_338),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_246),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_222),
.B(n_246),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_231),
.B2(n_232),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_225),
.B(n_231),
.C(n_233),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.C(n_229),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_230),
.B(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_234),
.B(n_237),
.C(n_243),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_262),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_247),
.B(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_250),
.A2(n_262),
.B1(n_263),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_251),
.Y(n_330)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_265),
.B(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_332),
.B(n_337),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_322),
.B(n_331),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_298),
.B(n_321),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_284),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_278),
.B1(n_282),
.B2(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_305),
.Y(n_304)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_296),
.C(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_307),
.B(n_320),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_302),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_316),
.B(n_319),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_315),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_325),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_336),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_345),
.C(n_346),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_353),
.B(n_354),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_351),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_382),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_381),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_372),
.B2(n_373),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B(n_371),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_378),
.B(n_380),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_374),
.B(n_378),
.Y(n_380)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);


endmodule