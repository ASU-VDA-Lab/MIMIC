module fake_aes_5693_n_533 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_533);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_533;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g77 ( .A(n_16), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_50), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_56), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_20), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_57), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_55), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_42), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_31), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_15), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_23), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_3), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_17), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_14), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
BUFx2_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_9), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_38), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_24), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_19), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_25), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_49), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_14), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_26), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_53), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_43), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_35), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_59), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_13), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_99), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_99), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_84), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
AND2x6_ASAP7_75t_L g118 ( .A(n_78), .B(n_36), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_96), .B(n_0), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_84), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_96), .Y(n_125) );
BUFx2_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_100), .B(n_1), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
AND2x4_ASAP7_75t_SL g130 ( .A(n_104), .B(n_39), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_89), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_90), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_131), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
OAI22xp33_ASAP7_75t_L g138 ( .A1(n_125), .A2(n_91), .B1(n_97), .B2(n_111), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_125), .B(n_98), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_114), .B(n_89), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_126), .B(n_81), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_114), .B(n_109), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_126), .B(n_109), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_113), .B(n_83), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_127), .B(n_103), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_131), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
INVx1_ASAP7_75t_SL g153 ( .A(n_128), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_134), .B(n_83), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_127), .B(n_79), .Y(n_156) );
BUFx4f_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_115), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_135), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_148), .B(n_128), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_152), .B(n_120), .Y(n_164) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_157), .B(n_130), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_153), .B(n_130), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_136), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_136), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_148), .B(n_130), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_157), .A2(n_123), .B(n_122), .C(n_91), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_152), .B(n_92), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_156), .B(n_122), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_143), .B(n_118), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_141), .B(n_118), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_157), .A2(n_123), .B(n_92), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_138), .B(n_112), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_144), .Y(n_188) );
AND2x6_ASAP7_75t_SL g189 ( .A(n_149), .B(n_97), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_152), .B(n_77), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
AOI222xp33_ASAP7_75t_L g193 ( .A1(n_163), .A2(n_154), .B1(n_86), .B2(n_88), .C1(n_157), .C2(n_118), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_192), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_161), .Y(n_195) );
BUFx2_ASAP7_75t_SL g196 ( .A(n_173), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_183), .B(n_152), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_177), .B(n_85), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_165), .A2(n_163), .B1(n_173), .B2(n_184), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_182), .B(n_118), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_165), .A2(n_80), .B1(n_108), .B2(n_94), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_185), .A2(n_159), .B(n_158), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_174), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_163), .A2(n_108), .B1(n_94), .B2(n_95), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_174), .Y(n_206) );
INVx8_ASAP7_75t_L g207 ( .A(n_190), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_187), .A2(n_95), .B(n_101), .C(n_106), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_173), .B(n_101), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_160), .B(n_93), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_162), .B(n_102), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_168), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_166), .A2(n_106), .B1(n_107), .B2(n_155), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_169), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g218 ( .A1(n_189), .A2(n_190), .B1(n_167), .B2(n_181), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
BUFx12f_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_175), .A2(n_107), .B(n_158), .C(n_155), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_190), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_206), .Y(n_225) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_223), .A2(n_186), .B(n_164), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_204), .B(n_178), .Y(n_227) );
CKINVDCx11_ASAP7_75t_R g228 ( .A(n_222), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_206), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_203), .A2(n_164), .B(n_176), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_217), .Y(n_231) );
CKINVDCx6p67_ASAP7_75t_R g232 ( .A(n_222), .Y(n_232) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_204), .A2(n_176), .B(n_191), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_204), .A2(n_181), .B(n_121), .Y(n_235) );
NOR2x1_ASAP7_75t_SL g236 ( .A(n_196), .B(n_194), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_217), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_208), .A2(n_175), .B(n_115), .C(n_119), .Y(n_238) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_195), .A2(n_121), .B(n_124), .Y(n_239) );
INVx6_ASAP7_75t_L g240 ( .A(n_207), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_194), .B(n_172), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_198), .A2(n_121), .B(n_124), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_214), .A2(n_172), .B1(n_170), .B2(n_178), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_216), .B(n_170), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_200), .B(n_178), .Y(n_245) );
CKINVDCx11_ASAP7_75t_R g246 ( .A(n_207), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_198), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_219), .A2(n_124), .B(n_147), .Y(n_249) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_219), .A2(n_147), .B(n_145), .Y(n_250) );
OAI211xp5_ASAP7_75t_L g251 ( .A1(n_246), .A2(n_218), .B(n_205), .C(n_193), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_245), .A2(n_214), .B1(n_196), .B2(n_202), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_231), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_234), .Y(n_254) );
AOI222xp33_ASAP7_75t_L g255 ( .A1(n_231), .A2(n_210), .B1(n_209), .B2(n_207), .C1(n_199), .C2(n_212), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_240), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_247), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_237), .B(n_209), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_238), .A2(n_200), .B(n_197), .C(n_225), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_238), .A2(n_229), .B(n_225), .C(n_244), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_211), .B(n_201), .C(n_224), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_229), .B(n_205), .Y(n_262) );
OAI221xp5_ASAP7_75t_SL g263 ( .A1(n_232), .A2(n_215), .B1(n_221), .B2(n_220), .C(n_119), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_245), .A2(n_207), .B1(n_220), .B2(n_221), .Y(n_264) );
OAI221xp5_ASAP7_75t_L g265 ( .A1(n_244), .A2(n_119), .B1(n_105), .B2(n_110), .C(n_132), .Y(n_265) );
HB1xp67_ASAP7_75t_SL g266 ( .A(n_247), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_247), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_248), .A2(n_213), .B1(n_119), .B2(n_132), .Y(n_268) );
AOI22xp33_ASAP7_75t_SL g269 ( .A1(n_236), .A2(n_213), .B1(n_133), .B2(n_132), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_248), .B(n_213), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g271 ( .A1(n_230), .A2(n_159), .B1(n_132), .B2(n_133), .C(n_213), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_253), .B(n_234), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_253), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_254), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_257), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_267), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_270), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_267), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_270), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_262), .B(n_234), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_262), .B(n_245), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_258), .B(n_259), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_258), .B(n_245), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
INVx4_ASAP7_75t_R g290 ( .A(n_266), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_264), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_256), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_275), .B(n_235), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_275), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_286), .B(n_235), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_291), .A2(n_255), .B1(n_252), .B2(n_240), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_273), .B(n_255), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_291), .A2(n_240), .B1(n_256), .B2(n_241), .Y(n_303) );
AOI222xp33_ASAP7_75t_L g304 ( .A1(n_287), .A2(n_251), .B1(n_236), .B2(n_228), .C1(n_265), .C2(n_240), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_286), .B(n_226), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_286), .B(n_226), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_285), .B(n_261), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_276), .B(n_250), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_280), .B(n_263), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_285), .B(n_230), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_232), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_285), .B(n_2), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_272), .Y(n_313) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_293), .A2(n_268), .B(n_265), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_282), .B(n_3), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_274), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_274), .Y(n_319) );
AOI21xp5_ASAP7_75t_SL g320 ( .A1(n_277), .A2(n_241), .B(n_271), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_272), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_287), .B(n_240), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_282), .B(n_269), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_311), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_313), .B(n_282), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_312), .B(n_277), .Y(n_328) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_304), .B(n_284), .C(n_288), .D(n_277), .Y(n_329) );
AND4x1_ASAP7_75t_L g330 ( .A(n_304), .B(n_290), .C(n_5), .D(n_6), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_296), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_302), .B(n_282), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_302), .B(n_288), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_313), .B(n_278), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_312), .B(n_278), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_317), .B(n_284), .Y(n_336) );
NAND2xp33_ASAP7_75t_SL g337 ( .A(n_299), .B(n_290), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_317), .B(n_274), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_296), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_321), .B(n_274), .Y(n_341) );
OAI33xp33_ASAP7_75t_L g342 ( .A1(n_311), .A2(n_289), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_301), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g344 ( .A(n_299), .B(n_283), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_321), .B(n_283), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_299), .B(n_279), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_295), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_297), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_309), .B(n_292), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_316), .B(n_292), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_301), .B(n_289), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_279), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g353 ( .A(n_300), .B(n_289), .C(n_7), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_305), .B(n_279), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_301), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_307), .B(n_289), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
AOI21xp33_ASAP7_75t_L g359 ( .A1(n_322), .A2(n_292), .B(n_281), .Y(n_359) );
NOR2xp67_ASAP7_75t_L g360 ( .A(n_315), .B(n_281), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_315), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_307), .B(n_279), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_308), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_309), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_305), .B(n_292), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_306), .B(n_292), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_364), .B(n_310), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_357), .B(n_306), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_367), .B(n_298), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_357), .B(n_298), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_361), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_358), .B(n_363), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_324), .B(n_298), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_330), .B(n_4), .Y(n_378) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_325), .B(n_318), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_332), .B(n_294), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_354), .B(n_318), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_325), .B(n_294), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_366), .B(n_294), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_325), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_356), .B(n_319), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_351), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_337), .B(n_281), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_361), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_365), .B(n_319), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_338), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_328), .B(n_319), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_335), .B(n_323), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_325), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_341), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_344), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_360), .B(n_323), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_327), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_346), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_333), .B(n_303), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_349), .B(n_4), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_347), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_345), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_346), .B(n_281), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_337), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_352), .B(n_314), .Y(n_409) );
NOR2x1p5_ASAP7_75t_L g410 ( .A(n_353), .B(n_281), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_348), .B(n_314), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_349), .B(n_314), .Y(n_412) );
NOR2x1_ASAP7_75t_R g413 ( .A(n_326), .B(n_241), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_340), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_326), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_362), .B(n_293), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_348), .B(n_314), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_340), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_397), .A2(n_320), .B1(n_350), .B2(n_359), .Y(n_420) );
OA22x2_ASAP7_75t_L g421 ( .A1(n_408), .A2(n_397), .B1(n_415), .B2(n_400), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_415), .B(n_293), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_378), .A2(n_329), .B1(n_320), .B2(n_132), .C(n_133), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_404), .B(n_342), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_402), .A2(n_342), .B(n_241), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_413), .A2(n_8), .B(n_9), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_404), .A2(n_133), .B1(n_117), .B2(n_129), .C(n_147), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_376), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_250), .B1(n_133), .B2(n_117), .Y(n_431) );
AOI31xp33_ASAP7_75t_SL g432 ( .A1(n_370), .A2(n_10), .A3(n_11), .B(n_12), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_410), .A2(n_243), .B1(n_227), .B2(n_250), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_394), .A2(n_250), .B1(n_117), .B2(n_129), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_400), .A2(n_129), .B1(n_117), .B2(n_227), .Y(n_435) );
NAND3x1_ASAP7_75t_L g436 ( .A(n_385), .B(n_10), .C(n_11), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_376), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_368), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_368), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_369), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_375), .A2(n_242), .B(n_239), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_379), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_382), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_369), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_394), .B(n_12), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_SL g446 ( .A1(n_389), .A2(n_15), .B(n_16), .C(n_17), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_416), .A2(n_227), .B1(n_129), .B2(n_117), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_388), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_129), .B1(n_233), .B2(n_242), .C1(n_239), .C2(n_249), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_407), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_383), .A2(n_213), .B1(n_145), .B2(n_142), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_396), .B(n_233), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_379), .Y(n_455) );
AOI322xp5_ASAP7_75t_L g456 ( .A1(n_384), .A2(n_145), .A3(n_142), .B1(n_140), .B2(n_137), .C1(n_29), .C2(n_30), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_399), .B(n_21), .Y(n_458) );
XNOR2x1_ASAP7_75t_L g459 ( .A(n_370), .B(n_22), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_405), .A2(n_142), .B1(n_140), .B2(n_137), .C(n_34), .Y(n_460) );
OAI21xp5_ASAP7_75t_SL g461 ( .A1(n_398), .A2(n_27), .B(n_28), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_398), .A2(n_140), .B(n_137), .C(n_249), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_390), .A2(n_32), .B(n_37), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_442), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_425), .B(n_419), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_452), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_461), .A2(n_406), .B(n_385), .C(n_383), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_457), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_421), .B(n_385), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_438), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_447), .B(n_419), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_439), .Y(n_473) );
XOR2x2_ASAP7_75t_L g474 ( .A(n_459), .B(n_377), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_423), .A2(n_398), .B1(n_409), .B2(n_373), .Y(n_475) );
AOI321xp33_ASAP7_75t_L g476 ( .A1(n_420), .A2(n_409), .A3(n_411), .B1(n_418), .B2(n_417), .C(n_405), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_445), .A2(n_399), .B1(n_396), .B2(n_387), .C(n_403), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_449), .A2(n_387), .B1(n_381), .B2(n_411), .C(n_418), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_426), .B(n_443), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_442), .B(n_395), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_430), .B(n_372), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_451), .A2(n_381), .B1(n_384), .B2(n_380), .C(n_391), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
AOI322xp5_ASAP7_75t_L g484 ( .A1(n_437), .A2(n_374), .A3(n_372), .B1(n_392), .B2(n_391), .C1(n_393), .C2(n_417), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_444), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_454), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_422), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_434), .B(n_392), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_428), .A2(n_417), .B1(n_383), .B2(n_406), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_455), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_427), .A2(n_393), .B1(n_374), .B2(n_406), .Y(n_491) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_434), .A2(n_386), .B(n_395), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_464), .B(n_490), .Y(n_493) );
AOI322xp5_ASAP7_75t_L g494 ( .A1(n_491), .A2(n_458), .A3(n_455), .B1(n_371), .B2(n_432), .C1(n_431), .C2(n_460), .Y(n_494) );
OAI21xp33_ASAP7_75t_SL g495 ( .A1(n_469), .A2(n_433), .B(n_463), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_483), .Y(n_496) );
OAI221xp5_ASAP7_75t_SL g497 ( .A1(n_476), .A2(n_456), .B1(n_462), .B2(n_386), .C(n_431), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_467), .A2(n_436), .B1(n_435), .B2(n_371), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_465), .B(n_441), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_469), .A2(n_448), .B1(n_453), .B2(n_446), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_489), .A2(n_429), .B1(n_450), .B2(n_140), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_485), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_485), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_480), .Y(n_504) );
NAND4xp25_ASAP7_75t_SL g505 ( .A(n_467), .B(n_40), .C(n_44), .D(n_46), .Y(n_505) );
OAI321xp33_ASAP7_75t_L g506 ( .A1(n_489), .A2(n_140), .A3(n_137), .B1(n_52), .B2(n_54), .C(n_60), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_474), .A2(n_140), .B1(n_137), .B2(n_61), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_488), .A2(n_137), .B1(n_51), .B2(n_62), .Y(n_508) );
AOI211xp5_ASAP7_75t_L g509 ( .A1(n_480), .A2(n_48), .B(n_63), .C(n_64), .Y(n_509) );
AOI311xp33_ASAP7_75t_L g510 ( .A1(n_498), .A2(n_477), .A3(n_478), .B(n_482), .C(n_487), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_495), .A2(n_484), .B(n_475), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_493), .B(n_481), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_500), .B(n_492), .C(n_486), .Y(n_513) );
OAI211xp5_ASAP7_75t_SL g514 ( .A1(n_494), .A2(n_472), .B(n_471), .C(n_468), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_504), .A2(n_466), .B1(n_473), .B2(n_470), .C(n_479), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_509), .B(n_503), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_502), .B(n_65), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_497), .A2(n_66), .B1(n_68), .B2(n_69), .C(n_70), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_516), .A2(n_505), .B(n_509), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_514), .B(n_499), .Y(n_520) );
XNOR2x1_ASAP7_75t_L g521 ( .A(n_510), .B(n_507), .Y(n_521) );
AND4x2_ASAP7_75t_L g522 ( .A(n_518), .B(n_506), .C(n_501), .D(n_508), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_512), .Y(n_523) );
OR4x2_ASAP7_75t_L g524 ( .A(n_521), .B(n_511), .C(n_513), .D(n_515), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_523), .B(n_496), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_519), .A2(n_517), .B1(n_72), .B2(n_73), .C(n_75), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_525), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_524), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_527), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g530 ( .A1(n_529), .A2(n_528), .B1(n_527), .B2(n_520), .Y(n_530) );
INVx4_ASAP7_75t_L g531 ( .A(n_530), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_531), .A2(n_528), .B1(n_526), .B2(n_522), .Y(n_532) );
AOI222xp33_ASAP7_75t_SL g533 ( .A1(n_532), .A2(n_71), .B1(n_76), .B2(n_528), .C1(n_530), .C2(n_529), .Y(n_533) );
endmodule