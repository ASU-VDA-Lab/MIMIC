module fake_aes_980_n_54 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_54);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_54;
wire n_53;
wire n_45;
wire n_38;
wire n_20;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_48;
wire n_30;
wire n_26;
wire n_33;
wire n_25;
wire n_50;
wire n_52;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_51;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_4), .B(n_15), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_7), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_9), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_4), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_0), .Y(n_22) );
AOI22x1_ASAP7_75t_SL g23 ( .A1(n_11), .A2(n_13), .B1(n_6), .B2(n_1), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_16), .Y(n_24) );
OA21x2_ASAP7_75t_L g25 ( .A1(n_12), .A2(n_8), .B(n_1), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_19), .B(n_0), .Y(n_27) );
BUFx8_ASAP7_75t_L g28 ( .A(n_21), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_22), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
OAI21x1_ASAP7_75t_L g31 ( .A1(n_27), .A2(n_24), .B(n_17), .Y(n_31) );
AND2x4_ASAP7_75t_L g32 ( .A(n_29), .B(n_22), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_32), .B(n_27), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_33), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
OAI21xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_31), .B(n_34), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_36), .B(n_33), .Y(n_39) );
OAI221xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_30), .B1(n_19), .B2(n_18), .C(n_24), .Y(n_40) );
OAI22xp33_ASAP7_75t_L g41 ( .A1(n_37), .A2(n_23), .B1(n_30), .B2(n_25), .Y(n_41) );
AOI22xp5_ASAP7_75t_L g42 ( .A1(n_37), .A2(n_28), .B1(n_23), .B2(n_32), .Y(n_42) );
AOI22xp5_ASAP7_75t_L g43 ( .A1(n_38), .A2(n_28), .B1(n_32), .B2(n_31), .Y(n_43) );
AND2x2_ASAP7_75t_L g44 ( .A(n_42), .B(n_32), .Y(n_44) );
NAND3xp33_ASAP7_75t_L g45 ( .A(n_41), .B(n_32), .C(n_25), .Y(n_45) );
AOI221xp5_ASAP7_75t_L g46 ( .A1(n_40), .A2(n_32), .B1(n_17), .B2(n_20), .C(n_31), .Y(n_46) );
O2A1O1Ixp33_ASAP7_75t_L g47 ( .A1(n_43), .A2(n_32), .B(n_20), .C(n_25), .Y(n_47) );
NOR2x1p5_ASAP7_75t_L g48 ( .A(n_45), .B(n_2), .Y(n_48) );
NAND3xp33_ASAP7_75t_L g49 ( .A(n_44), .B(n_31), .C(n_3), .Y(n_49) );
AND2x4_ASAP7_75t_L g50 ( .A(n_46), .B(n_2), .Y(n_50) );
OAI22xp5_ASAP7_75t_L g51 ( .A1(n_48), .A2(n_47), .B1(n_5), .B2(n_6), .Y(n_51) );
INVx1_ASAP7_75t_L g52 ( .A(n_50), .Y(n_52) );
OAI22xp5_ASAP7_75t_L g53 ( .A1(n_52), .A2(n_49), .B1(n_5), .B2(n_3), .Y(n_53) );
OAI21xp33_ASAP7_75t_L g54 ( .A1(n_53), .A2(n_51), .B(n_14), .Y(n_54) );
endmodule