module real_aes_7795_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g433 ( .A(n_0), .Y(n_433) );
INVx1_ASAP7_75t_L g534 ( .A(n_1), .Y(n_534) );
INVx1_ASAP7_75t_L g140 ( .A(n_2), .Y(n_140) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_3), .A2(n_447), .B1(n_732), .B2(n_733), .C1(n_742), .C2(n_744), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_4), .A2(n_39), .B1(n_165), .B2(n_480), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g172 ( .A1(n_5), .A2(n_156), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_6), .B(n_154), .Y(n_546) );
AND2x6_ASAP7_75t_L g133 ( .A(n_7), .B(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_8), .A2(n_243), .B(n_244), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_9), .B(n_40), .Y(n_434) );
INVx1_ASAP7_75t_L g178 ( .A(n_10), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_11), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g125 ( .A(n_12), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_13), .B(n_146), .Y(n_489) );
INVx1_ASAP7_75t_L g249 ( .A(n_14), .Y(n_249) );
INVx1_ASAP7_75t_L g528 ( .A(n_15), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_16), .B(n_121), .Y(n_517) );
AO32x2_ASAP7_75t_L g501 ( .A1(n_17), .A2(n_120), .A3(n_154), .B1(n_482), .B2(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_18), .B(n_165), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_19), .B(n_161), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_20), .B(n_121), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_21), .A2(n_50), .B1(n_165), .B2(n_480), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_22), .B(n_156), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_23), .A2(n_99), .B1(n_739), .B2(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_23), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_24), .A2(n_76), .B1(n_146), .B2(n_165), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_25), .B(n_165), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_26), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_27), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_28), .B(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_29), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_30), .B(n_151), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_31), .B(n_144), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g110 ( .A1(n_32), .A2(n_89), .B1(n_111), .B2(n_112), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_32), .Y(n_111) );
INVx1_ASAP7_75t_L g193 ( .A(n_33), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_34), .B(n_151), .Y(n_473) );
INVx2_ASAP7_75t_L g131 ( .A(n_35), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_36), .B(n_165), .Y(n_550) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_37), .A2(n_104), .B1(n_438), .B2(n_445), .C1(n_747), .C2(n_750), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_37), .A2(n_69), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_37), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_37), .B(n_151), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_38), .A2(n_133), .B(n_136), .C(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g191 ( .A(n_41), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_42), .B(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_43), .B(n_165), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_44), .A2(n_87), .B1(n_213), .B2(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_45), .B(n_165), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_46), .B(n_165), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_47), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_48), .B(n_533), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_49), .B(n_156), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_51), .A2(n_61), .B1(n_146), .B2(n_165), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_52), .A2(n_737), .B1(n_738), .B2(n_741), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_52), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_53), .A2(n_136), .B1(n_146), .B2(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_54), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_55), .B(n_165), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_56), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_57), .B(n_165), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_58), .A2(n_164), .B(n_176), .C(n_177), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_59), .Y(n_226) );
INVx1_ASAP7_75t_L g174 ( .A(n_60), .Y(n_174) );
INVx1_ASAP7_75t_L g134 ( .A(n_62), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_63), .B(n_165), .Y(n_535) );
INVx1_ASAP7_75t_L g124 ( .A(n_64), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_65), .Y(n_441) );
AO32x2_ASAP7_75t_L g477 ( .A1(n_66), .A2(n_154), .A3(n_229), .B1(n_478), .B2(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g553 ( .A(n_67), .Y(n_553) );
INVx1_ASAP7_75t_L g468 ( .A(n_68), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_69), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_SL g160 ( .A1(n_70), .A2(n_161), .B(n_162), .C(n_164), .Y(n_160) );
INVxp67_ASAP7_75t_L g163 ( .A(n_71), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_72), .B(n_146), .Y(n_469) );
INVx1_ASAP7_75t_L g444 ( .A(n_73), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_74), .Y(n_196) );
INVx1_ASAP7_75t_L g219 ( .A(n_75), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_77), .A2(n_133), .B(n_136), .C(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_78), .B(n_480), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_79), .B(n_146), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_80), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_80), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_81), .B(n_141), .Y(n_209) );
INVx2_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_83), .B(n_161), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_84), .B(n_146), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_85), .A2(n_133), .B(n_136), .C(n_139), .Y(n_135) );
OR2x2_ASAP7_75t_L g430 ( .A(n_86), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g450 ( .A(n_86), .B(n_432), .Y(n_450) );
INVx2_ASAP7_75t_L g455 ( .A(n_86), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_88), .A2(n_102), .B1(n_146), .B2(n_147), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_89), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_90), .B(n_151), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_91), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_92), .A2(n_133), .B(n_136), .C(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_93), .Y(n_239) );
INVx1_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_95), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_96), .B(n_141), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_97), .B(n_146), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_98), .B(n_154), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_99), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_100), .A2(n_156), .B(n_157), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_101), .B(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_427), .B(n_435), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B1(n_425), .B2(n_426), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_106), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_109), .Y(n_426) );
XNOR2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .Y(n_109) );
INVx1_ASAP7_75t_L g451 ( .A(n_113), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_113), .A2(n_452), .B1(n_457), .B2(n_743), .Y(n_742) );
NAND2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_341), .Y(n_113) );
NOR5xp2_ASAP7_75t_L g114 ( .A(n_115), .B(n_264), .C(n_296), .D(n_311), .E(n_328), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_180), .B(n_201), .C(n_252), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_152), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_117), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_117), .B(n_316), .Y(n_379) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_118), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_118), .B(n_198), .Y(n_265) );
AND2x2_ASAP7_75t_L g306 ( .A(n_118), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_118), .B(n_275), .Y(n_310) );
OR2x2_ASAP7_75t_L g347 ( .A(n_118), .B(n_186), .Y(n_347) );
INVx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g185 ( .A(n_119), .B(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g255 ( .A(n_119), .Y(n_255) );
OR2x2_ASAP7_75t_L g418 ( .A(n_119), .B(n_258), .Y(n_418) );
AO21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_126), .B(n_148), .Y(n_119) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_120), .A2(n_187), .B(n_195), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_120), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g214 ( .A(n_120), .Y(n_214) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_122), .B(n_123), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_135), .Y(n_126) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_128), .A2(n_166), .B1(n_188), .B2(n_194), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_128), .A2(n_219), .B(n_220), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
AND2x4_ASAP7_75t_L g156 ( .A(n_129), .B(n_133), .Y(n_156) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g533 ( .A(n_130), .Y(n_533) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx1_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
INVx3_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
INVx1_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_132), .Y(n_190) );
INVx4_ASAP7_75t_SL g166 ( .A(n_133), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_133), .A2(n_467), .B(n_470), .Y(n_466) );
BUFx3_ASAP7_75t_L g482 ( .A(n_133), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_133), .A2(n_487), .B(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_133), .A2(n_527), .B(n_531), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_133), .A2(n_540), .B(n_543), .Y(n_539) );
INVx5_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
BUFx3_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
INVx1_ASAP7_75t_L g480 ( .A(n_137), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_143), .C(n_145), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_SL g467 ( .A1(n_141), .A2(n_164), .B(n_468), .C(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g504 ( .A(n_141), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_141), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_141), .A2(n_550), .B(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_142), .B(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_142), .B(n_178), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g478 ( .A1(n_142), .A2(n_144), .B1(n_479), .B2(n_481), .Y(n_478) );
INVx2_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx4_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_144), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_144), .A2(n_504), .B1(n_520), .B2(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_145), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_150), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_150), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_151), .A2(n_242), .B(n_251), .Y(n_241) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_151), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_151), .A2(n_486), .B(n_494), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_152), .A2(n_321), .B1(n_322), .B2(n_325), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_152), .B(n_255), .Y(n_404) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_170), .Y(n_152) );
AND2x2_ASAP7_75t_L g200 ( .A(n_153), .B(n_186), .Y(n_200) );
AND2x2_ASAP7_75t_L g257 ( .A(n_153), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g262 ( .A(n_153), .Y(n_262) );
INVx3_ASAP7_75t_L g275 ( .A(n_153), .Y(n_275) );
OR2x2_ASAP7_75t_L g295 ( .A(n_153), .B(n_258), .Y(n_295) );
AND2x2_ASAP7_75t_L g314 ( .A(n_153), .B(n_171), .Y(n_314) );
BUFx2_ASAP7_75t_L g346 ( .A(n_153), .Y(n_346) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_167), .Y(n_153) );
INVx4_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_154), .A2(n_539), .B(n_546), .Y(n_538) );
BUFx2_ASAP7_75t_L g243 ( .A(n_156), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_160), .C(n_166), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_158), .A2(n_166), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_158), .A2(n_166), .B(n_245), .C(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g490 ( .A(n_161), .Y(n_490) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_165), .Y(n_236) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_168), .A2(n_172), .B(n_179), .Y(n_171) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_169), .B(n_216), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_169), .B(n_482), .C(n_519), .Y(n_518) );
AO21x1_ASAP7_75t_L g608 ( .A1(n_169), .A2(n_519), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g261 ( .A(n_170), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
BUFx2_ASAP7_75t_L g184 ( .A(n_171), .Y(n_184) );
INVx2_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
OR2x2_ASAP7_75t_L g277 ( .A(n_171), .B(n_258), .Y(n_277) );
AND2x2_ASAP7_75t_L g307 ( .A(n_171), .B(n_186), .Y(n_307) );
AND2x2_ASAP7_75t_L g324 ( .A(n_171), .B(n_255), .Y(n_324) );
AND2x2_ASAP7_75t_L g364 ( .A(n_171), .B(n_275), .Y(n_364) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_171), .B(n_200), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_176), .A2(n_492), .B(n_493), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g552 ( .A1(n_176), .A2(n_532), .B(n_553), .C(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp33_ASAP7_75t_SL g181 ( .A(n_182), .B(n_197), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_185), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_183), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OAI21xp33_ASAP7_75t_L g338 ( .A1(n_184), .A2(n_200), .B(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_184), .B(n_186), .Y(n_394) );
AND2x2_ASAP7_75t_L g330 ( .A(n_185), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_186), .Y(n_356) );
OAI22xp5_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_189) );
INVx2_ASAP7_75t_L g192 ( .A(n_190), .Y(n_192) );
INVx4_ASAP7_75t_L g247 ( .A(n_190), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_197), .B(n_255), .Y(n_423) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_198), .A2(n_366), .B1(n_367), .B2(n_372), .Y(n_365) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AND2x2_ASAP7_75t_L g256 ( .A(n_199), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g294 ( .A(n_199), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g331 ( .A(n_199), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_200), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g385 ( .A(n_200), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_227), .Y(n_202) );
INVx4_ASAP7_75t_L g271 ( .A(n_203), .Y(n_271) );
AND2x2_ASAP7_75t_L g349 ( .A(n_203), .B(n_316), .Y(n_349) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_217), .Y(n_203) );
INVx3_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_204), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
INVx2_ASAP7_75t_L g300 ( .A(n_204), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_204), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g357 ( .A(n_204), .B(n_352), .Y(n_357) );
AND2x2_ASAP7_75t_L g422 ( .A(n_204), .B(n_392), .Y(n_422) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
AOI21xp5_ASAP7_75t_SL g205 ( .A1(n_206), .A2(n_207), .B(n_214), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
INVx1_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_214), .A2(n_526), .B(n_536), .Y(n_525) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_214), .A2(n_548), .B(n_555), .Y(n_547) );
AND2x2_ASAP7_75t_L g263 ( .A(n_217), .B(n_241), .Y(n_263) );
INVx2_ASAP7_75t_L g283 ( .A(n_217), .Y(n_283) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
INVx1_ASAP7_75t_L g288 ( .A(n_227), .Y(n_288) );
AND2x2_ASAP7_75t_L g334 ( .A(n_227), .B(n_282), .Y(n_334) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_240), .Y(n_227) );
INVx2_ASAP7_75t_L g273 ( .A(n_228), .Y(n_273) );
INVx1_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
AND2x2_ASAP7_75t_L g299 ( .A(n_228), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_228), .B(n_283), .Y(n_337) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_236), .Y(n_232) );
AND2x2_ASAP7_75t_L g316 ( .A(n_240), .B(n_273), .Y(n_316) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
AND2x2_ASAP7_75t_L g352 ( .A(n_241), .B(n_283), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_247), .B(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_247), .A2(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g530 ( .A(n_247), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_259), .B(n_263), .Y(n_252) );
INVx1_ASAP7_75t_SL g297 ( .A(n_253), .Y(n_297) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_254), .B(n_261), .Y(n_354) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g303 ( .A(n_255), .B(n_258), .Y(n_303) );
AND2x2_ASAP7_75t_L g332 ( .A(n_255), .B(n_276), .Y(n_332) );
OR2x2_ASAP7_75t_L g335 ( .A(n_255), .B(n_295), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_256), .A2(n_348), .B1(n_400), .B2(n_401), .C1(n_403), .C2(n_405), .Y(n_399) );
BUFx2_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g302 ( .A(n_261), .B(n_303), .Y(n_302) );
INVx3_ASAP7_75t_SL g319 ( .A(n_261), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_261), .B(n_313), .Y(n_373) );
AND2x2_ASAP7_75t_L g308 ( .A(n_263), .B(n_268), .Y(n_308) );
INVx1_ASAP7_75t_L g327 ( .A(n_263), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g264 ( .A1(n_265), .A2(n_266), .B1(n_270), .B2(n_274), .C(n_278), .Y(n_264) );
OR2x2_ASAP7_75t_L g336 ( .A(n_266), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_291), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_268), .B(n_281), .Y(n_361) );
AND2x2_ASAP7_75t_L g366 ( .A(n_268), .B(n_316), .Y(n_366) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_268), .Y(n_376) );
NAND2x1_ASAP7_75t_SL g387 ( .A(n_268), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g272 ( .A(n_269), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_269), .B(n_287), .Y(n_318) );
INVx1_ASAP7_75t_L g384 ( .A(n_269), .Y(n_384) );
INVx1_ASAP7_75t_L g359 ( .A(n_270), .Y(n_359) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g371 ( .A(n_271), .Y(n_371) );
NOR2xp67_ASAP7_75t_L g383 ( .A(n_271), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g388 ( .A(n_272), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_272), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g291 ( .A(n_273), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_273), .B(n_283), .Y(n_304) );
INVx1_ASAP7_75t_L g370 ( .A(n_273), .Y(n_370) );
INVx1_ASAP7_75t_L g391 ( .A(n_274), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_284), .B(n_293), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
AND2x2_ASAP7_75t_L g424 ( .A(n_280), .B(n_357), .Y(n_424) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g392 ( .A(n_281), .B(n_352), .Y(n_392) );
AOI32xp33_ASAP7_75t_L g305 ( .A1(n_282), .A2(n_288), .A3(n_306), .B1(n_308), .B2(n_309), .Y(n_305) );
AOI322xp5_ASAP7_75t_L g407 ( .A1(n_282), .A2(n_314), .A3(n_397), .B1(n_408), .B2(n_409), .C1(n_410), .C2(n_412), .Y(n_407) );
INVx2_ASAP7_75t_L g287 ( .A(n_283), .Y(n_287) );
INVx1_ASAP7_75t_L g397 ( .A(n_283), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B1(n_289), .B2(n_290), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_285), .B(n_291), .Y(n_340) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_286), .B(n_352), .Y(n_402) );
INVx1_ASAP7_75t_L g289 ( .A(n_287), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_287), .B(n_316), .Y(n_406) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_295), .B(n_390), .Y(n_389) );
OAI221xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_298), .B1(n_301), .B2(n_304), .C(n_305), .Y(n_296) );
OR2x2_ASAP7_75t_L g317 ( .A(n_298), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g351 ( .A(n_299), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g355 ( .A(n_309), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_317), .B2(n_319), .C(n_320), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_313), .A2(n_344), .B1(n_348), .B2(n_349), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_314), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_314), .Y(n_419) );
INVx1_ASAP7_75t_L g413 ( .A(n_316), .Y(n_413) );
INVx1_ASAP7_75t_SL g348 ( .A(n_317), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_319), .B(n_347), .Y(n_409) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_324), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g390 ( .A(n_324), .Y(n_390) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
OAI221xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_333), .B1(n_335), .B2(n_336), .C(n_338), .Y(n_328) );
NOR2xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_330), .A2(n_348), .B1(n_394), .B2(n_395), .Y(n_393) );
CKINVDCx14_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_335), .A2(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR3xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_374), .C(n_398), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_350), .C(n_358), .D(n_365), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g421 ( .A(n_346), .Y(n_421) );
INVx3_ASAP7_75t_SL g415 ( .A(n_347), .Y(n_415) );
OR2x2_ASAP7_75t_L g420 ( .A(n_347), .B(n_421), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B1(n_355), .B2(n_357), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_352), .B(n_370), .Y(n_411) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI21xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_360), .B(n_362), .Y(n_358) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_377), .B(n_380), .C(n_393), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B1(n_386), .B2(n_389), .C1(n_391), .C2(n_392), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND4xp25_ASAP7_75t_SL g417 ( .A(n_390), .B(n_418), .C(n_419), .D(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND3xp33_ASAP7_75t_SL g398 ( .A(n_399), .B(n_407), .C(n_416), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_416) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp33_ASAP7_75t_L g748 ( .A(n_428), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_431), .B(n_455), .Y(n_746) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g454 ( .A(n_432), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_437), .A2(n_441), .B(n_442), .Y(n_751) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g749 ( .A(n_441), .B(n_443), .Y(n_749) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B1(n_452), .B2(n_456), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g743 ( .A(n_449), .Y(n_743) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_653), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_602), .C(n_644), .Y(n_458) );
AOI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_511), .B(n_556), .C(n_578), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_474), .B(n_495), .C(n_506), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_462), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g665 ( .A(n_462), .B(n_582), .Y(n_665) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g567 ( .A(n_463), .B(n_498), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_463), .B(n_485), .Y(n_684) );
INVx1_ASAP7_75t_L g702 ( .A(n_463), .Y(n_702) );
AND2x2_ASAP7_75t_L g711 ( .A(n_463), .B(n_599), .Y(n_711) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g594 ( .A(n_464), .B(n_485), .Y(n_594) );
AND2x2_ASAP7_75t_L g652 ( .A(n_464), .B(n_599), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_464), .Y(n_696) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g573 ( .A(n_465), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g581 ( .A(n_465), .Y(n_581) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_465), .Y(n_621) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
AND2x2_ASAP7_75t_L g560 ( .A(n_476), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g593 ( .A(n_476), .Y(n_593) );
OR2x2_ASAP7_75t_L g719 ( .A(n_476), .B(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_476), .B(n_485), .Y(n_723) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx1_ASAP7_75t_L g509 ( .A(n_477), .Y(n_509) );
AND2x2_ASAP7_75t_L g582 ( .A(n_477), .B(n_500), .Y(n_582) );
AND2x2_ASAP7_75t_L g622 ( .A(n_477), .B(n_501), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_482), .A2(n_549), .B(n_552), .Y(n_548) );
INVxp67_ASAP7_75t_L g664 ( .A(n_483), .Y(n_664) );
AND2x4_ASAP7_75t_L g689 ( .A(n_483), .B(n_582), .Y(n_689) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_484), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g499 ( .A(n_485), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g568 ( .A(n_485), .B(n_501), .Y(n_568) );
INVx1_ASAP7_75t_L g574 ( .A(n_485), .Y(n_574) );
INVx2_ASAP7_75t_L g600 ( .A(n_485), .Y(n_600) );
AND2x2_ASAP7_75t_L g616 ( .A(n_485), .B(n_617), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_496), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
AND2x2_ASAP7_75t_L g679 ( .A(n_498), .B(n_500), .Y(n_679) );
AND2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_581), .Y(n_596) );
AND2x2_ASAP7_75t_L g695 ( .A(n_499), .B(n_696), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_500), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g720 ( .A(n_500), .B(n_581), .Y(n_720) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g510 ( .A(n_501), .Y(n_510) );
AND2x2_ASAP7_75t_L g599 ( .A(n_501), .B(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_504), .A2(n_532), .B(n_534), .C(n_535), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_504), .A2(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AND2x2_ASAP7_75t_L g645 ( .A(n_508), .B(n_580), .Y(n_645) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_509), .B(n_581), .Y(n_630) );
INVx2_ASAP7_75t_L g629 ( .A(n_510), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_510), .A2(n_573), .B1(n_634), .B2(n_636), .C1(n_637), .C2(n_640), .Y(n_633) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g558 ( .A(n_515), .Y(n_558) );
OR2x2_ASAP7_75t_L g669 ( .A(n_515), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_516), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g648 ( .A(n_516), .B(n_562), .Y(n_648) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_522), .A2(n_612), .B1(n_651), .B2(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_537), .Y(n_522) );
INVx3_ASAP7_75t_L g584 ( .A(n_523), .Y(n_584) );
OR2x2_ASAP7_75t_L g717 ( .A(n_523), .B(n_593), .Y(n_717) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g590 ( .A(n_524), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g606 ( .A(n_524), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g614 ( .A(n_524), .B(n_562), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_524), .B(n_538), .Y(n_670) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g561 ( .A(n_525), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g565 ( .A(n_525), .B(n_538), .Y(n_565) );
AND2x2_ASAP7_75t_L g641 ( .A(n_525), .B(n_588), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_525), .B(n_547), .Y(n_681) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_537), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_558), .Y(n_597) );
AND2x2_ASAP7_75t_L g601 ( .A(n_537), .B(n_591), .Y(n_601) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
INVx3_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
AND2x2_ASAP7_75t_L g587 ( .A(n_538), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g722 ( .A(n_538), .B(n_705), .Y(n_722) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_547), .Y(n_576) );
INVx2_ASAP7_75t_L g588 ( .A(n_547), .Y(n_588) );
AND2x2_ASAP7_75t_L g632 ( .A(n_547), .B(n_608), .Y(n_632) );
INVx1_ASAP7_75t_L g675 ( .A(n_547), .Y(n_675) );
OR2x2_ASAP7_75t_L g706 ( .A(n_547), .B(n_608), .Y(n_706) );
AND2x2_ASAP7_75t_L g726 ( .A(n_547), .B(n_562), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g564 ( .A(n_558), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_558), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g683 ( .A(n_560), .Y(n_683) );
INVx2_ASAP7_75t_SL g577 ( .A(n_561), .Y(n_577) );
AND2x2_ASAP7_75t_L g697 ( .A(n_561), .B(n_591), .Y(n_697) );
INVx2_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_562), .B(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_569), .B2(n_575), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_565), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g731 ( .A(n_565), .Y(n_731) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g656 ( .A(n_567), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_567), .B(n_599), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_568), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_568), .B(n_621), .Y(n_672) );
INVx2_ASAP7_75t_L g728 ( .A(n_568), .Y(n_728) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_571), .B(n_616), .Y(n_649) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_573), .B(n_593), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g710 ( .A(n_576), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_577), .A2(n_661), .B(n_663), .C(n_666), .Y(n_660) );
OR2x2_ASAP7_75t_L g687 ( .A(n_577), .B(n_591), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_583), .B1(n_585), .B2(n_592), .C(n_595), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_580), .B(n_629), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_580), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g714 ( .A(n_580), .Y(n_714) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_581), .Y(n_605) );
INVx1_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_584), .B(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g692 ( .A(n_584), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_584), .B(n_632), .Y(n_708) );
INVx2_ASAP7_75t_L g694 ( .A(n_585), .Y(n_694) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g635 ( .A(n_587), .B(n_606), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_587), .A2(n_603), .B(n_645), .C(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g613 ( .A(n_588), .B(n_608), .Y(n_613) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_592), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g661 ( .A(n_593), .B(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_598), .B2(n_601), .Y(n_595) );
INVx1_ASAP7_75t_L g715 ( .A(n_597), .Y(n_715) );
INVx1_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
AOI211xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_606), .B(n_610), .C(n_633), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g625 ( .A(n_605), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g676 ( .A(n_606), .Y(n_676) );
AND2x2_ASAP7_75t_L g725 ( .A(n_606), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_615), .B(n_623), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx2_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_613), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g631 ( .A(n_614), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g707 ( .A(n_614), .Y(n_707) );
OAI32xp33_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_666), .A3(n_673), .B1(n_714), .B2(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_SL g686 ( .A(n_616), .Y(n_686) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g626 ( .A(n_622), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_631), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_625), .A2(n_673), .B1(n_699), .B2(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_629), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g666 ( .A(n_632), .Y(n_666) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_652), .A2(n_694), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g653 ( .A(n_654), .B(n_677), .C(n_693), .D(n_703), .E(n_721), .Y(n_653) );
AOI211xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_667), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g724 ( .A(n_661), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_SL g700 ( .A(n_670), .Y(n_700) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_673), .A2(n_683), .A3(n_684), .B1(n_685), .B2(n_686), .C1(n_687), .C2(n_688), .Y(n_682) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g685 ( .A(n_675), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_675), .B(n_700), .Y(n_699) );
AOI211xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_680), .B(n_682), .C(n_690), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_686), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g729 ( .A(n_696), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_711), .B1(n_712), .B2(n_716), .C(n_718), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_708), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g730 ( .A(n_706), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .C(n_727), .Y(n_721) );
AOI21xp33_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_729), .B(n_730), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
endmodule